
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_jnc, ABINPUT, ABINPUT000, ABINPUT000000);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  input [8:0] ABINPUT;
  input [16:0] ABINPUT000;
  input [16:0] ABINPUT000000;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire cy_reg;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [16:0] \oc8051_top_1.ABINPUT000 ;
  wire [16:0] \oc8051_top_1.ABINPUT000000 ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire \oc8051_top_1.decoder_new_valid_pc ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT000 ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire \oc8051_top_1.oc8051_alu1.divOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.mulOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire \oc8051_top_1.oc8051_decoder1.new_valid_pc ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire \oc8051_top_1.pc_log_change ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  wire pc_log_change;
  wire pc_log_change_r;
  output property_invalid_jnc;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not _13450_ (_05110_, rst);
  not _13451_ (_05111_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not _13452_ (_05112_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  not _13453_ (_05113_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _13454_ (_05114_, _05113_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand _13455_ (_05115_, _05114_, _05112_);
  or _13456_ (_05116_, _05115_, _05111_);
  not _13457_ (_05117_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not _13458_ (_05118_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _13459_ (_05119_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], _05113_);
  nand _13460_ (_05120_, _05119_, _05118_);
  or _13461_ (_05121_, _05120_, _05117_);
  and _13462_ (_05122_, _05121_, _05116_);
  not _13463_ (_05123_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _13464_ (_05124_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _13465_ (_05125_, _05124_, _05113_);
  nor _13466_ (_05126_, _05125_, _05123_);
  and _13467_ (_05127_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand _13468_ (_05128_, _05127_, _05112_);
  not _13469_ (_05129_, _05128_);
  and _13470_ (_05130_, _05129_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _13471_ (_05131_, _05130_, _05126_);
  and _13472_ (_05132_, _05131_, _05122_);
  nor _13473_ (_05133_, _05124_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not _13474_ (_05134_, _05133_);
  not _13475_ (_05135_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _13476_ (_05136_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _05135_);
  or _13477_ (_05137_, _05136_, ABINPUT[5]);
  nand _13478_ (_05138_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _05135_);
  or _13479_ (_05139_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _13480_ (_05140_, _05139_, _05137_);
  or _13481_ (_05141_, _05140_, _05134_);
  not _13482_ (_05142_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _13483_ (_05143_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand _13484_ (_05144_, _05143_, _05113_);
  nor _13485_ (_05145_, _05144_, _05142_);
  and _13486_ (_05146_, _05127_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _13487_ (_05147_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor _13488_ (_05148_, _05147_, _05145_);
  and _13489_ (_05149_, _05148_, _05141_);
  and _13490_ (_05150_, _05149_, _05132_);
  not _13491_ (_05151_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _13492_ (_05152_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _05151_);
  and _13493_ (_05153_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _05151_);
  nor _13494_ (_05154_, _05153_, _05152_);
  and _13495_ (_05155_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _05151_);
  and _13496_ (_05156_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _05151_);
  nor _13497_ (_05157_, _05156_, _05155_);
  and _13498_ (_05158_, _05157_, _05154_);
  not _13499_ (_05159_, _05158_);
  not _13500_ (_05160_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  not _13501_ (_05162_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _13502_ (_05163_, _05152_, _05162_);
  nand _13503_ (_05164_, _05163_, _05160_);
  nand _13504_ (_05165_, _05154_, _05156_);
  and _13505_ (_05166_, _05165_, _05164_);
  and _13506_ (_05167_, _05166_, _05159_);
  and _13507_ (_05168_, _05153_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  nand _13508_ (_05169_, _05168_, _05160_);
  not _13509_ (_05170_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _13510_ (_05171_, _05153_, _05170_);
  and _13511_ (_05172_, _05171_, _05155_);
  not _13512_ (_05174_, _05172_);
  and _13513_ (_05175_, _05174_, _05169_);
  and _13514_ (_05176_, _05175_, _05167_);
  nor _13515_ (_05177_, _05176_, _05150_);
  not _13516_ (_05178_, _05177_);
  and _13517_ (_05180_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _13518_ (_05181_, _05180_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _13519_ (_05182_, _05181_);
  or _13520_ (_05183_, _05136_, ABINPUT[0]);
  or _13521_ (_05184_, _05138_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and _13522_ (_05185_, _05184_, _05183_);
  or _13523_ (_05186_, _05185_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and _13524_ (_05187_, _05186_, _05182_);
  not _13525_ (_05188_, _05187_);
  not _13526_ (_05189_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or _13527_ (_05190_, _05115_, _05189_);
  not _13528_ (_05191_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or _13529_ (_05192_, _05120_, _05191_);
  and _13530_ (_05193_, _05192_, _05190_);
  nand _13531_ (_05194_, _05129_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _13532_ (_05195_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _13533_ (_05196_, _05125_, _05195_);
  and _13534_ (_05197_, _05196_, _05194_);
  and _13535_ (_05198_, _05197_, _05193_);
  or _13536_ (_05199_, _05136_, ABINPUT[4]);
  or _13537_ (_05200_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _13538_ (_05201_, _05200_, _05199_);
  or _13539_ (_05202_, _05201_, _05134_);
  nand _13540_ (_05203_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  not _13541_ (_05204_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _13542_ (_05206_, _05144_, _05204_);
  and _13543_ (_05207_, _05206_, _05203_);
  and _13544_ (_05209_, _05207_, _05202_);
  and _13545_ (_05210_, _05209_, _05198_);
  not _13546_ (_05211_, _05210_);
  not _13547_ (_05212_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or _13548_ (_05213_, _05115_, _05212_);
  not _13549_ (_05214_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  or _13550_ (_05215_, _05120_, _05214_);
  and _13551_ (_05217_, _05215_, _05213_);
  not _13552_ (_05218_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _13553_ (_05219_, _05125_, _05218_);
  not _13554_ (_05220_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _13555_ (_05221_, _05128_, _05220_);
  and _13556_ (_05222_, _05221_, _05219_);
  and _13557_ (_05223_, _05222_, _05217_);
  or _13558_ (_05224_, _05136_, ABINPUT[3]);
  or _13559_ (_05225_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _13560_ (_05226_, _05225_, _05224_);
  or _13561_ (_05227_, _05226_, _05134_);
  not _13562_ (_05228_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _13563_ (_05229_, _05144_, _05228_);
  nand _13564_ (_05230_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  and _13565_ (_05231_, _05230_, _05229_);
  and _13566_ (_05232_, _05231_, _05227_);
  and _13567_ (_05233_, _05232_, _05223_);
  not _13568_ (_05234_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  or _13569_ (_05235_, _05115_, _05234_);
  not _13570_ (_05236_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  or _13571_ (_05237_, _05120_, _05236_);
  and _13572_ (_05238_, _05237_, _05235_);
  nand _13573_ (_05239_, _05129_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _13574_ (_05240_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _13575_ (_05241_, _05125_, _05240_);
  and _13576_ (_05242_, _05241_, _05239_);
  and _13577_ (_05243_, _05242_, _05238_);
  or _13578_ (_05244_, _05136_, ABINPUT[1]);
  or _13579_ (_05245_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand _13580_ (_05246_, _05245_, _05244_);
  or _13581_ (_05247_, _05246_, _05134_);
  nand _13582_ (_05248_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  not _13583_ (_05249_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _13584_ (_05250_, _05144_, _05249_);
  and _13585_ (_05251_, _05250_, _05248_);
  and _13586_ (_05252_, _05251_, _05247_);
  and _13587_ (_05253_, _05252_, _05243_);
  or _13588_ (_05254_, _05136_, ABINPUT[2]);
  or _13589_ (_05255_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _13590_ (_05256_, _05255_, _05254_);
  or _13591_ (_05257_, _05256_, _05134_);
  not _13592_ (_05258_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or _13593_ (_05259_, _05115_, _05258_);
  not _13594_ (_05260_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  or _13595_ (_05261_, _05120_, _05260_);
  and _13596_ (_05262_, _05261_, _05259_);
  and _13597_ (_05263_, _05262_, _05257_);
  not _13598_ (_05264_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _13599_ (_05265_, _05125_, _05264_);
  not _13600_ (_05266_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _13601_ (_05267_, _05128_, _05266_);
  and _13602_ (_05268_, _05267_, _05265_);
  not _13603_ (_05269_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _13604_ (_05270_, _05144_, _05269_);
  nand _13605_ (_05271_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _13606_ (_05272_, _05271_, _05270_);
  and _13607_ (_05273_, _05272_, _05268_);
  and _13608_ (_05274_, _05273_, _05263_);
  and _13609_ (_05275_, _05274_, _05253_);
  nand _13610_ (_05276_, _05275_, _05233_);
  or _13611_ (_05277_, _05276_, _05211_);
  or _13612_ (_05278_, _05277_, _05188_);
  not _13613_ (_05279_, _05233_);
  nand _13614_ (_05280_, _05252_, _05243_);
  nand _13615_ (_05281_, _05273_, _05263_);
  and _13616_ (_05282_, _05281_, _05280_);
  nand _13617_ (_05283_, _05282_, _05279_);
  or _13618_ (_05284_, _05283_, _05210_);
  or _13619_ (_05285_, _05284_, _05187_);
  and _13620_ (_05286_, _05285_, _05278_);
  or _13621_ (_05287_, _05286_, _05150_);
  not _13622_ (_05288_, _05155_);
  nor _13623_ (_05290_, _05288_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _13624_ (_05291_, _05168_, _05290_);
  nand _13625_ (_05292_, _05286_, _05150_);
  and _13626_ (_05293_, _05292_, _05291_);
  nand _13627_ (_05294_, _05293_, _05287_);
  and _13628_ (_05295_, _05171_, _05157_);
  nor _13629_ (_05296_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not _13630_ (_05297_, _05296_);
  nor _13631_ (_05298_, _05297_, _05140_);
  not _13632_ (_05299_, _05298_);
  and _13633_ (_05300_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _13634_ (_05301_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  not _13635_ (_05302_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _13636_ (_05303_, _05302_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _13637_ (_05304_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _13638_ (_05305_, _05304_, _05301_);
  and _13639_ (_05306_, _05305_, _05299_);
  nor _13640_ (_05307_, _05306_, _05150_);
  and _13641_ (_05308_, _05306_, _05150_);
  nor _13642_ (_05309_, _05308_, _05307_);
  nand _13643_ (_05310_, _05309_, _05295_);
  and _13644_ (_05311_, _05155_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _13645_ (_05312_, _05311_, _05163_);
  and _13646_ (_05313_, _05312_, _05307_);
  and _13647_ (_05314_, _05290_, _05163_);
  and _13648_ (_05316_, _05314_, _05150_);
  nor _13649_ (_05317_, _05316_, _05313_);
  and _13650_ (_05318_, _05188_, _05150_);
  not _13651_ (_05319_, _05318_);
  and _13652_ (_05320_, _05168_, _05311_);
  not _13653_ (_05321_, _05320_);
  and _13654_ (_05322_, _05306_, _05187_);
  nor _13655_ (_05323_, _05322_, _05321_);
  and _13656_ (_05324_, _05323_, _05319_);
  and _13657_ (_05325_, _05156_, _05160_);
  and _13658_ (_05326_, _05171_, _05325_);
  not _13659_ (_05327_, _05326_);
  nor _13660_ (_05328_, _05327_, _05308_);
  nor _13661_ (_05329_, _05328_, _05324_);
  and _13662_ (_05330_, _05329_, _05317_);
  and _13663_ (_05332_, _05330_, _05310_);
  and _13664_ (_05333_, _05332_, _05294_);
  and _13665_ (_05334_, _05333_, _05178_);
  not _13666_ (_05335_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _13667_ (_05336_, \oc8051_top_1.oc8051_decoder1.wr , _05151_);
  and _13668_ (_05337_, _05336_, _05335_);
  not _13669_ (_05338_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _13670_ (_05339_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _05151_);
  and _13671_ (_05340_, _05339_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _13672_ (_05341_, _05340_, _05338_);
  and _13673_ (_05343_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _13674_ (_05344_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _13675_ (_05345_, _05344_, _05343_);
  and _13676_ (_05346_, _05345_, _05341_);
  and _13677_ (_05347_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _05151_);
  nor _13678_ (_05348_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _13679_ (_05349_, _05348_, _05347_);
  and _13680_ (_05350_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor _13681_ (_05351_, _05350_, _05346_);
  not _13682_ (_05352_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _13683_ (_05353_, _05339_, _05352_);
  nand _13684_ (_05354_, _05353_, _05338_);
  or _13685_ (_05355_, _05354_, _05258_);
  and _13686_ (_05356_, _05353_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nand _13687_ (_05357_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nor _13688_ (_05358_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nor _13689_ (_05359_, _05358_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _13690_ (_05361_, _05359_, _05339_);
  nand _13691_ (_05362_, _05361_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and _13692_ (_05363_, _05362_, _05357_);
  and _13693_ (_05364_, _05363_, _05355_);
  and _13694_ (_05365_, _05364_, _05351_);
  and _13695_ (_05366_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _13696_ (_05367_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _13697_ (_05368_, _05367_, _05366_);
  not _13698_ (_05369_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _13699_ (_05370_, _05341_, _05369_);
  or _13700_ (_05371_, _05354_, _05234_);
  nand _13701_ (_05372_, _05361_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nand _13702_ (_05373_, _05372_, _05371_);
  nor _13703_ (_05374_, _05373_, _05370_);
  and _13704_ (_05375_, _05374_, _05368_);
  and _13705_ (_05376_, _05375_, _05365_);
  nand _13706_ (_05377_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or _13707_ (_05378_, _05354_, _05189_);
  and _13708_ (_05379_, _05378_, _05377_);
  and _13709_ (_05380_, _05343_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nand _13710_ (_05381_, _05380_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  or _13711_ (_05382_, _05380_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _13712_ (_05383_, _05382_, _05381_);
  nand _13713_ (_05384_, _05383_, _05341_);
  nand _13714_ (_05385_, _05361_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nand _13715_ (_05386_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  and _13716_ (_05387_, _05386_, _05385_);
  and _13717_ (_05388_, _05387_, _05384_);
  and _13718_ (_05389_, _05388_, _05379_);
  not _13719_ (_05390_, _05389_);
  nor _13720_ (_05391_, _05343_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _13721_ (_05392_, _05391_, _05380_);
  and _13722_ (_05393_, _05392_, _05341_);
  and _13723_ (_05394_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _13724_ (_05395_, _05394_, _05393_);
  or _13725_ (_05396_, _05354_, _05212_);
  nand _13726_ (_05397_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  nand _13727_ (_05398_, _05361_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  and _13728_ (_05399_, _05398_, _05397_);
  and _13729_ (_05400_, _05399_, _05396_);
  and _13730_ (_05401_, _05400_, _05395_);
  and _13731_ (_05402_, _05401_, _05390_);
  and _13732_ (_05403_, _05402_, _05376_);
  and _13733_ (_05404_, _05380_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _13734_ (_05405_, _05404_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or _13735_ (_05406_, _05404_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nand _13736_ (_05407_, _05406_, _05341_);
  or _13737_ (_05408_, _05407_, _05405_);
  nand _13738_ (_05409_, _05356_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nand _13739_ (_05410_, _05340_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nand _13740_ (_05411_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  and _13741_ (_05412_, _05411_, _05410_);
  and _13742_ (_05413_, _05412_, _05409_);
  or _13743_ (_05414_, _05354_, _05111_);
  nand _13744_ (_05415_, _05361_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and _13745_ (_05416_, _05415_, _05414_);
  and _13746_ (_05417_, _05416_, _05413_);
  and _13747_ (_05418_, _05417_, _05408_);
  not _13748_ (_05419_, _05418_);
  nand _13749_ (_05420_, _05405_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  or _13750_ (_05421_, _05405_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _13751_ (_05422_, _05421_, _05341_);
  nand _13752_ (_05423_, _05422_, _05420_);
  nand _13753_ (_05424_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  not _13754_ (_05425_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or _13755_ (_05426_, _05354_, _05425_);
  nand _13756_ (_05427_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _13757_ (_05429_, _05427_, _05410_);
  and _13758_ (_05431_, _05429_, _05426_);
  and _13759_ (_05432_, _05431_, _05424_);
  and _13760_ (_05433_, _05432_, _05423_);
  and _13761_ (_05434_, _05433_, _05419_);
  and _13762_ (_05435_, _05405_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nand _13763_ (_05436_, _05435_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  or _13764_ (_05437_, _05435_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and _13765_ (_05438_, _05437_, _05341_);
  nand _13766_ (_05439_, _05438_, _05436_);
  nand _13767_ (_05440_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not _13768_ (_05441_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  or _13769_ (_05442_, _05354_, _05441_);
  nand _13770_ (_05443_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _13771_ (_05444_, _05443_, _05410_);
  and _13772_ (_05445_, _05444_, _05442_);
  and _13773_ (_05446_, _05445_, _05440_);
  and _13774_ (_05447_, _05446_, _05439_);
  not _13775_ (_05448_, _05447_);
  nand _13776_ (_05449_, _05436_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  or _13777_ (_05450_, _05436_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand _13778_ (_05451_, _05450_, _05449_);
  nand _13779_ (_05452_, _05451_, _05341_);
  nand _13780_ (_05453_, _05356_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  not _13781_ (_05454_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  or _13782_ (_05455_, _05354_, _05454_);
  nand _13783_ (_05456_, _05349_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and _13784_ (_05457_, _05456_, _05410_);
  and _13785_ (_05458_, _05457_, _05455_);
  and _13786_ (_05459_, _05458_, _05453_);
  nand _13787_ (_05460_, _05459_, _05452_);
  nor _13788_ (_05461_, _05460_, _05448_);
  and _13789_ (_05462_, _05461_, _05434_);
  and _13790_ (_05463_, _05462_, _05403_);
  and _13791_ (_05464_, _05463_, _05337_);
  not _13792_ (_05465_, _05464_);
  nor _13793_ (_05466_, _05465_, _05334_);
  not _13794_ (_05467_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor _13795_ (_05468_, _05464_, _05467_);
  or _13796_ (_05469_, _05468_, _05466_);
  and _13797_ (_05161_, _05469_, _05110_);
  not _13798_ (_05470_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  nor _13799_ (_05471_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _13800_ (_05472_, _05471_, _05470_);
  nor _13801_ (_05473_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  and _13802_ (_05474_, _05473_, _05151_);
  and _13803_ (_05475_, _05474_, _05472_);
  and _13804_ (pc_log_change, _05475_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or _13805_ (_05476_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  not _13806_ (_05478_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _13807_ (_05479_, pc_log_change, _05478_);
  and _13808_ (_05480_, _05479_, _05110_);
  and _13809_ (_06782_, _05480_, _05476_);
  and _13810_ (_05481_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _13811_ (_05482_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _13812_ (_05483_, pc_log_change, _05482_);
  or _13813_ (_05484_, _05483_, _05481_);
  and _13814_ (_06919_, _05484_, _05110_);
  not _13815_ (_05485_, _05401_);
  not _13816_ (_05486_, _05365_);
  and _13817_ (_05487_, _05375_, _05486_);
  and _13818_ (_05488_, _05487_, _05485_);
  and _13819_ (_05489_, _05325_, _05154_);
  not _13820_ (_05490_, _05489_);
  nor _13821_ (_05491_, _05115_, _05454_);
  not _13822_ (_05492_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor _13823_ (_05493_, _05120_, _05492_);
  nor _13824_ (_05494_, _05493_, _05491_);
  and _13825_ (_05495_, _05129_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not _13826_ (_05496_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _13827_ (_05497_, _05125_, _05496_);
  nor _13828_ (_05498_, _05497_, _05495_);
  and _13829_ (_05499_, _05498_, _05494_);
  nor _13830_ (_05500_, _05136_, ABINPUT[8]);
  nor _13831_ (_05501_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nor _13832_ (_05502_, _05501_, _05500_);
  and _13833_ (_05503_, _05502_, _05133_);
  not _13834_ (_05504_, _05503_);
  and _13835_ (_05505_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  not _13836_ (_05506_, _05144_);
  and _13837_ (_05507_, _05506_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _13838_ (_05508_, _05507_, _05505_);
  and _13839_ (_05509_, _05508_, _05504_);
  and _13840_ (_05510_, _05509_, _05499_);
  and _13841_ (_05511_, _05502_, _05296_);
  not _13842_ (_05512_, _05511_);
  and _13843_ (_05514_, _05300_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and _13844_ (_05515_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _13845_ (_05516_, _05515_, _05514_);
  and _13846_ (_05517_, _05516_, _05512_);
  nor _13847_ (_05518_, _05517_, _05510_);
  not _13848_ (_05519_, _05518_);
  and _13849_ (_05520_, _05517_, _05510_);
  or _13850_ (_05521_, _05297_, _05201_);
  and _13851_ (_05522_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _13852_ (_05523_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _13853_ (_05524_, _05523_, _05522_);
  and _13854_ (_05526_, _05524_, _05521_);
  nor _13855_ (_05527_, _05526_, _05210_);
  and _13856_ (_05528_, _05526_, _05210_);
  nor _13857_ (_05529_, _05528_, _05527_);
  or _13858_ (_05530_, _05297_, _05226_);
  and _13859_ (_05531_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and _13860_ (_05532_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _13861_ (_05533_, _05532_, _05531_);
  and _13862_ (_05534_, _05533_, _05530_);
  nor _13863_ (_05535_, _05534_, _05233_);
  not _13864_ (_05536_, _05535_);
  and _13865_ (_05537_, _05534_, _05233_);
  nor _13866_ (_05538_, _05537_, _05535_);
  or _13867_ (_05539_, _05297_, _05256_);
  nand _13868_ (_05540_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand _13869_ (_05541_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _13870_ (_05542_, _05541_, _05540_);
  nand _13871_ (_05543_, _05542_, _05539_);
  and _13872_ (_05544_, _05543_, _05281_);
  or _13873_ (_05545_, _05297_, _05246_);
  nand _13874_ (_05546_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nand _13875_ (_05547_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _13876_ (_05548_, _05547_, _05546_);
  and _13877_ (_05549_, _05548_, _05545_);
  not _13878_ (_05550_, _05549_);
  and _13879_ (_05551_, _05550_, _05280_);
  and _13880_ (_05552_, _05542_, _05539_);
  and _13881_ (_05553_, _05552_, _05274_);
  nor _13882_ (_05554_, _05553_, _05544_);
  and _13883_ (_05555_, _05554_, _05551_);
  or _13884_ (_05556_, _05555_, _05544_);
  nand _13885_ (_05557_, _05556_, _05538_);
  nand _13886_ (_05558_, _05557_, _05536_);
  nand _13887_ (_05559_, _05558_, _05529_);
  or _13888_ (_05560_, _05558_, _05529_);
  and _13889_ (_05561_, _05560_, _05559_);
  and _13890_ (_05562_, _05549_, _05253_);
  nor _13891_ (_05563_, _05562_, _05551_);
  and _13892_ (_05564_, _05563_, _05187_);
  and _13893_ (_05566_, _05564_, _05554_);
  or _13894_ (_05567_, _05556_, _05538_);
  and _13895_ (_05568_, _05567_, _05557_);
  and _13896_ (_05570_, _05568_, _05566_);
  and _13897_ (_05571_, _05570_, _05561_);
  not _13898_ (_05572_, _05528_);
  and _13899_ (_05573_, _05558_, _05572_);
  or _13900_ (_05574_, _05573_, _05527_);
  or _13901_ (_05575_, _05574_, _05571_);
  nand _13902_ (_05576_, _05575_, _05309_);
  nor _13903_ (_05577_, _05115_, _05425_);
  not _13904_ (_05578_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor _13905_ (_05579_, _05120_, _05578_);
  nor _13906_ (_05580_, _05579_, _05577_);
  not _13907_ (_05581_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _13908_ (_05582_, _05125_, _05581_);
  not _13909_ (_05583_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _13910_ (_05584_, _05128_, _05583_);
  nor _13911_ (_05585_, _05584_, _05582_);
  and _13912_ (_05586_, _05585_, _05580_);
  nor _13913_ (_05587_, _05136_, ABINPUT[6]);
  nor _13914_ (_05588_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nor _13915_ (_05589_, _05588_, _05587_);
  and _13916_ (_05590_, _05589_, _05133_);
  not _13917_ (_05591_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _13918_ (_05592_, _05144_, _05591_);
  and _13919_ (_05593_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  nor _13920_ (_05594_, _05593_, _05592_);
  not _13921_ (_05595_, _05594_);
  nor _13922_ (_05596_, _05595_, _05590_);
  and _13923_ (_05597_, _05596_, _05586_);
  and _13924_ (_05598_, _05589_, _05296_);
  not _13925_ (_05599_, _05598_);
  and _13926_ (_05600_, _05300_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _13927_ (_05601_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _13928_ (_05602_, _05601_, _05600_);
  and _13929_ (_05603_, _05602_, _05599_);
  and _13930_ (_05604_, _05603_, _05597_);
  nor _13931_ (_05605_, _05603_, _05597_);
  nor _13932_ (_05606_, _05605_, _05604_);
  not _13933_ (_05607_, _05606_);
  or _13934_ (_05608_, _05607_, _05576_);
  nor _13935_ (_05609_, _05115_, _05441_);
  not _13936_ (_05610_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nor _13937_ (_05611_, _05120_, _05610_);
  nor _13938_ (_05612_, _05611_, _05609_);
  not _13939_ (_05613_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _13940_ (_05614_, _05125_, _05613_);
  and _13941_ (_05615_, _05129_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _13942_ (_05616_, _05615_, _05614_);
  and _13943_ (_05617_, _05616_, _05612_);
  nor _13944_ (_05618_, _05136_, ABINPUT[7]);
  nor _13945_ (_05619_, _05138_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nor _13946_ (_05620_, _05619_, _05618_);
  and _13947_ (_05621_, _05620_, _05133_);
  not _13948_ (_05622_, _05621_);
  and _13949_ (_05623_, _05506_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _13950_ (_05624_, _05146_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor _13951_ (_05625_, _05624_, _05623_);
  and _13952_ (_05626_, _05625_, _05622_);
  and _13953_ (_05627_, _05626_, _05617_);
  and _13954_ (_05628_, _05620_, _05296_);
  not _13955_ (_05629_, _05628_);
  and _13956_ (_05630_, _05300_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  and _13957_ (_05631_, _05303_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _13958_ (_05632_, _05631_, _05630_);
  and _13959_ (_05633_, _05632_, _05629_);
  nor _13960_ (_05634_, _05633_, _05627_);
  and _13961_ (_05635_, _05633_, _05627_);
  nor _13962_ (_05636_, _05635_, _05634_);
  not _13963_ (_05637_, _05636_);
  and _13964_ (_05638_, _05606_, _05307_);
  nor _13965_ (_05639_, _05638_, _05605_);
  nor _13966_ (_05640_, _05639_, _05637_);
  and _13967_ (_05641_, _05639_, _05637_);
  nor _13968_ (_05642_, _05641_, _05640_);
  not _13969_ (_05643_, _05642_);
  or _13970_ (_05644_, _05643_, _05608_);
  nor _13971_ (_05645_, _05640_, _05634_);
  and _13972_ (_05646_, _05645_, _05644_);
  or _13973_ (_05647_, _05646_, _05520_);
  and _13974_ (_05648_, _05647_, _05519_);
  or _13975_ (_05649_, _05648_, _05490_);
  and _13976_ (_05650_, _05290_, _05154_);
  not _13977_ (_05651_, _05650_);
  not _13978_ (_05652_, _05517_);
  and _13979_ (_05653_, _05652_, _05510_);
  nor _13980_ (_05654_, _05520_, _05518_);
  not _13981_ (_05655_, _05633_);
  nor _13982_ (_05656_, _05655_, _05627_);
  not _13983_ (_05658_, _05597_);
  and _13984_ (_05659_, _05603_, _05658_);
  not _13985_ (_05661_, _05306_);
  and _13986_ (_05662_, _05661_, _05150_);
  nor _13987_ (_05663_, _05606_, _05662_);
  nor _13988_ (_05664_, _05663_, _05659_);
  nor _13989_ (_05666_, _05664_, _05636_);
  nor _13990_ (_05667_, _05666_, _05656_);
  and _13991_ (_05668_, _05664_, _05636_);
  nor _13992_ (_05669_, _05668_, _05666_);
  not _13993_ (_05671_, _05669_);
  and _13994_ (_05672_, _05606_, _05662_);
  nor _13995_ (_05673_, _05672_, _05663_);
  not _13996_ (_05674_, _05673_);
  not _13997_ (_05675_, _05309_);
  and _13998_ (_05676_, _05550_, _05253_);
  or _13999_ (_05677_, _05676_, _05554_);
  or _14000_ (_05678_, _05543_, _05274_);
  and _14001_ (_05679_, _05678_, _05677_);
  or _14002_ (_05681_, _05679_, _05538_);
  not _14003_ (_05682_, _05534_);
  or _14004_ (_05683_, _05682_, _05233_);
  and _14005_ (_05684_, _05683_, _05681_);
  nor _14006_ (_05685_, _05684_, _05529_);
  and _14007_ (_05686_, _05684_, _05529_);
  or _14008_ (_05687_, _05686_, _05685_);
  and _14009_ (_05689_, _05679_, _05538_);
  not _14010_ (_05690_, _05689_);
  nand _14011_ (_05692_, _05690_, _05681_);
  and _14012_ (_05693_, _05676_, _05554_);
  not _14013_ (_05694_, _05693_);
  nand _14014_ (_05696_, _05694_, _05677_);
  nor _14015_ (_05697_, _05563_, _05188_);
  and _14016_ (_05699_, _05697_, _05696_);
  and _14017_ (_05700_, _05699_, _05692_);
  and _14018_ (_05702_, _05700_, _05687_);
  not _14019_ (_05703_, _05526_);
  or _14020_ (_05705_, _05703_, _05210_);
  and _14021_ (_05707_, _05703_, _05210_);
  or _14022_ (_05708_, _05684_, _05707_);
  and _14023_ (_05710_, _05708_, _05705_);
  or _14024_ (_05711_, _05710_, _05702_);
  and _14025_ (_05713_, _05711_, _05675_);
  and _14026_ (_05714_, _05713_, _05674_);
  and _14027_ (_05715_, _05714_, _05671_);
  nor _14028_ (_05716_, _05715_, _05667_);
  nor _14029_ (_05717_, _05716_, _05654_);
  nor _14030_ (_05718_, _05717_, _05653_);
  or _14031_ (_05719_, _05718_, _05651_);
  and _14032_ (_05720_, _05627_, _05597_);
  not _14033_ (_05722_, _05720_);
  not _14034_ (_05723_, _05150_);
  and _14035_ (_05725_, _05325_, _05163_);
  and _14036_ (_05726_, _05274_, _05233_);
  nor _14037_ (_05728_, _05726_, _05210_);
  and _14038_ (_05729_, _05728_, _05725_);
  and _14039_ (_05731_, _05729_, _05723_);
  nor _14040_ (_05732_, _05731_, _05722_);
  nor _14041_ (_05734_, _05732_, _05510_);
  nor _14042_ (_05735_, _05734_, _05187_);
  not _14043_ (_05736_, _05735_);
  not _14044_ (_05737_, _05725_);
  nor _14045_ (_05738_, _05510_, _05188_);
  not _14046_ (_05739_, _05738_);
  nor _14047_ (_05740_, _05739_, _05732_);
  nor _14048_ (_05741_, _05740_, _05737_);
  and _14049_ (_05742_, _05741_, _05736_);
  not _14050_ (_05743_, _05729_);
  and _14051_ (_05744_, _05168_, _05325_);
  and _14052_ (_05746_, _05280_, _05744_);
  and _14053_ (_05747_, _05185_, _05181_);
  and _14054_ (_05749_, _05171_, _05290_);
  and _14055_ (_05751_, _05312_, _05185_);
  nor _14056_ (_05752_, _05751_, _05749_);
  nor _14057_ (_05753_, _05752_, _05747_);
  nor _14058_ (_05754_, _05753_, _05746_);
  nor _14059_ (_05755_, _05187_, _05185_);
  not _14060_ (_05756_, _05295_);
  and _14061_ (_05758_, _05187_, _05185_);
  or _14062_ (_05759_, _05758_, _05756_);
  and _14063_ (_05760_, _05759_, _05327_);
  or _14064_ (_05761_, _05760_, _05755_);
  and _14065_ (_05762_, _05171_, _05311_);
  not _14066_ (_05763_, _05762_);
  nor _14067_ (_05764_, _05510_, _05763_);
  nor _14068_ (_05765_, _05314_, _05187_);
  and _14069_ (_05766_, _05168_, _05157_);
  not _14070_ (_05767_, _05185_);
  nand _14071_ (_05768_, _05767_, _05766_);
  and _14072_ (_05769_, _05768_, _05159_);
  and _14073_ (_05770_, _05769_, _05187_);
  nor _14074_ (_05771_, _05770_, _05765_);
  nor _14075_ (_05773_, _05771_, _05764_);
  and _14076_ (_05774_, _05773_, _05761_);
  and _14077_ (_05776_, _05774_, _05754_);
  and _14078_ (_05777_, _05776_, _05743_);
  not _14079_ (_05778_, _05777_);
  nor _14080_ (_05779_, _05778_, _05742_);
  and _14081_ (_05781_, _05779_, _05719_);
  nand _14082_ (_05782_, _05781_, _05649_);
  and _14083_ (_05784_, _05782_, _05488_);
  and _14084_ (_05785_, _05401_, _05375_);
  or _14085_ (_05786_, _05376_, _05785_);
  and _14086_ (_05787_, _05786_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _14087_ (_05788_, _05787_, _05784_);
  and _14088_ (_05789_, _05447_, _05433_);
  not _14089_ (_05790_, _05341_);
  not _14090_ (_05791_, _05336_);
  nor _14091_ (_05792_, _05349_, _05791_);
  and _14092_ (_05793_, _05792_, _05790_);
  and _14093_ (_05794_, _05793_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _14094_ (_05795_, _05794_, _05390_);
  and _14095_ (_05796_, _05795_, _05418_);
  and _14096_ (_05797_, _05796_, _05460_);
  and _14097_ (_05798_, _05797_, _05789_);
  and _14098_ (_05799_, _05798_, _05788_);
  nand _14099_ (_05800_, _05798_, _05375_);
  and _14100_ (_05801_, _05800_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _14101_ (_05802_, _05433_, _05418_);
  and _14102_ (_05803_, _05460_, _05447_);
  and _14103_ (_05804_, _05803_, _05802_);
  and _14104_ (_05805_, _05376_, _05401_);
  and _14105_ (_05806_, _05793_, _05335_);
  and _14106_ (_05807_, _05806_, _05390_);
  and _14107_ (_05808_, _05807_, _05805_);
  and _14108_ (_05809_, _05808_, _05804_);
  or _14109_ (_05810_, _05809_, _05801_);
  or _14110_ (_05811_, _05810_, _05799_);
  nor _14111_ (_05812_, _05633_, _05188_);
  nor _14112_ (_05813_, _05627_, _05187_);
  or _14113_ (_05814_, _05813_, _05812_);
  and _14114_ (_05815_, _05814_, _05320_);
  not _14115_ (_05816_, _05627_);
  or _14116_ (_05817_, _05277_, _05723_);
  or _14117_ (_05818_, _05658_, _05817_);
  nand _14118_ (_05819_, _05818_, _05187_);
  or _14119_ (_05820_, _05597_, _05150_);
  nor _14120_ (_05821_, _05820_, _05284_);
  or _14121_ (_05822_, _05821_, _05187_);
  and _14122_ (_05823_, _05822_, _05819_);
  nand _14123_ (_05824_, _05823_, _05816_);
  or _14124_ (_05825_, _05823_, _05816_);
  and _14125_ (_05826_, _05825_, _05291_);
  and _14126_ (_05827_, _05826_, _05824_);
  nor _14127_ (_05828_, _05827_, _05815_);
  nor _14128_ (_05829_, _05627_, _05176_);
  not _14129_ (_05830_, _05829_);
  and _14130_ (_05831_, _05636_, _05295_);
  not _14131_ (_05832_, _05831_);
  nor _14132_ (_05833_, _05635_, _05327_);
  not _14133_ (_05834_, _05833_);
  and _14134_ (_05835_, _05634_, _05312_);
  and _14135_ (_05836_, _05627_, _05314_);
  nor _14136_ (_05837_, _05836_, _05835_);
  and _14137_ (_05838_, _05837_, _05834_);
  and _14138_ (_05839_, _05838_, _05832_);
  and _14139_ (_05840_, _05839_, _05830_);
  and _14140_ (_05841_, _05840_, _05828_);
  nand _14141_ (_05842_, _05841_, _05809_);
  and _14142_ (_05843_, _05842_, _05110_);
  and _14143_ (_07249_, _05843_, _05811_);
  not _14144_ (_05844_, _05809_);
  nor _14145_ (_05845_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _14146_ (_05846_, _05845_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  not _14147_ (_05847_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _14148_ (_05848_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and _14149_ (_05849_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _14150_ (_05850_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _14151_ (_05851_, _05850_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor _14152_ (_05852_, _05851_, _05849_);
  nor _14153_ (_05853_, _05852_, _05848_);
  or _14154_ (_05854_, _05853_, _05847_);
  and _14155_ (_05855_, _05850_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _14156_ (_05856_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _14157_ (_05857_, _05856_, _05855_);
  nor _14158_ (_05858_, _05857_, _05848_);
  and _14159_ (_05859_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _14160_ (_05860_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _05850_);
  nor _14161_ (_05861_, _05860_, _05859_);
  nand _14162_ (_05862_, _05861_, _05858_);
  or _14163_ (_05863_, _05862_, _05854_);
  and _14164_ (_05864_, _05863_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _14165_ (_05865_, _05864_, _05846_);
  nor _14166_ (_05866_, _05375_, _05365_);
  and _14167_ (_05867_, _05866_, _05485_);
  and _14168_ (_05868_, _05867_, _05804_);
  and _14169_ (_05869_, _05868_, _05795_);
  or _14170_ (_05870_, _05869_, _05865_);
  and _14171_ (_05871_, _05870_, _05844_);
  and _14172_ (_05872_, _05781_, _05649_);
  nand _14173_ (_05873_, _05869_, _05872_);
  and _14174_ (_05874_, _05873_, _05871_);
  and _14175_ (_05875_, _05821_, _05816_);
  and _14176_ (_05876_, _05875_, _05188_);
  nor _14177_ (_05877_, _05722_, _05817_);
  and _14178_ (_05878_, _05877_, _05187_);
  nor _14179_ (_05879_, _05878_, _05876_);
  and _14180_ (_05880_, _05879_, _05510_);
  not _14181_ (_05881_, _05880_);
  not _14182_ (_05882_, _05291_);
  nor _14183_ (_05883_, _05879_, _05510_);
  nor _14184_ (_05884_, _05883_, _05882_);
  and _14185_ (_05885_, _05884_, _05881_);
  and _14186_ (_05886_, _05510_, _05188_);
  not _14187_ (_05887_, _05886_);
  and _14188_ (_05888_, _05517_, _05187_);
  nor _14189_ (_05889_, _05888_, _05321_);
  and _14190_ (_05890_, _05889_, _05887_);
  nor _14191_ (_05891_, _05890_, _05885_);
  and _14192_ (_05892_, _05518_, _05312_);
  and _14193_ (_05893_, _05510_, _05314_);
  nor _14194_ (_05894_, _05893_, _05892_);
  nor _14195_ (_05895_, _05510_, _05176_);
  and _14196_ (_05896_, _05654_, _05295_);
  nor _14197_ (_05897_, _05520_, _05327_);
  or _14198_ (_05898_, _05897_, _05896_);
  nor _14199_ (_05899_, _05898_, _05895_);
  and _14200_ (_05900_, _05899_, _05894_);
  and _14201_ (_05901_, _05900_, _05891_);
  nor _14202_ (_05902_, _05901_, _05844_);
  or _14203_ (_05903_, _05902_, _05874_);
  and _14204_ (_07357_, _05903_, _05110_);
  not _14205_ (_05904_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand _14206_ (_05905_, _05853_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor _14207_ (_05906_, _05861_, _05848_);
  or _14208_ (_05907_, _05906_, _05858_);
  or _14209_ (_05908_, _05907_, _05905_);
  and _14210_ (_05909_, _05908_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _14211_ (_05910_, _05909_, _05904_);
  not _14212_ (_05911_, _05375_);
  and _14213_ (_05912_, _05911_, _05365_);
  and _14214_ (_05913_, _05912_, _05402_);
  and _14215_ (_05914_, _05804_, _05913_);
  and _14216_ (_05915_, _05914_, _05794_);
  or _14217_ (_05916_, _05915_, _05910_);
  and _14218_ (_05917_, _05916_, _05844_);
  nand _14219_ (_05918_, _05915_, _05872_);
  and _14220_ (_05919_, _05918_, _05917_);
  and _14221_ (_05920_, _05543_, _05320_);
  nor _14222_ (_05921_, _05282_, _05275_);
  or _14223_ (_05922_, _05921_, _05187_);
  nand _14224_ (_05923_, _05921_, _05187_);
  and _14225_ (_05924_, _05923_, _05291_);
  and _14226_ (_05925_, _05924_, _05922_);
  nor _14227_ (_05926_, _05925_, _05920_);
  or _14228_ (_05927_, _05553_, _05327_);
  or _14229_ (_05928_, _05553_, _05544_);
  or _14230_ (_05929_, _05928_, _05756_);
  and _14231_ (_05930_, _05929_, _05927_);
  nand _14232_ (_05931_, _05544_, _05312_);
  not _14233_ (_05932_, _05314_);
  or _14234_ (_05933_, _05932_, _05281_);
  and _14235_ (_05934_, _05933_, _05931_);
  or _14236_ (_05935_, _05274_, _05176_);
  and _14237_ (_05936_, _05935_, _05934_);
  and _14238_ (_05937_, _05936_, _05930_);
  and _14239_ (_05938_, _05937_, _05926_);
  nor _14240_ (_05939_, _05938_, _05844_);
  or _14241_ (_05940_, _05939_, _05919_);
  and _14242_ (_07655_, _05940_, _05110_);
  and _14243_ (_05941_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _05848_);
  not _14244_ (_05942_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _14245_ (_05943_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _14246_ (_05944_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _14247_ (_05945_, _05944_, _05943_);
  and _14248_ (_05946_, _05945_, _05942_);
  not _14249_ (_05947_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _14250_ (_05948_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _14251_ (_05949_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor _14252_ (_05950_, _05949_, _05948_);
  and _14253_ (_05951_, _05950_, _05947_);
  nor _14254_ (_05952_, _05951_, _05946_);
  not _14255_ (_05953_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _14256_ (_05954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _14257_ (_05955_, _05954_, _05953_);
  not _14258_ (_05956_, _05955_);
  not _14259_ (_05957_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _14260_ (_05958_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _14261_ (_05959_, _05958_, _05957_);
  not _14262_ (_05960_, _05959_);
  not _14263_ (_05961_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _14264_ (_05962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _14265_ (_05963_, _05962_, _05961_);
  not _14266_ (_05964_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _14267_ (_05965_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _14268_ (_05966_, _05965_, _05964_);
  nor _14269_ (_05967_, _05966_, _05963_);
  and _14270_ (_05968_, _05967_, _05960_);
  and _14271_ (_05969_, _05968_, _05956_);
  nand _14272_ (_05970_, _05969_, _05952_);
  nand _14273_ (_05971_, _05970_, _05941_);
  nand _14274_ (_05972_, _05945_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _14275_ (_05973_, _05950_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _14276_ (_05974_, _05973_);
  and _14277_ (_05975_, _05974_, _05972_);
  and _14278_ (_05976_, _05958_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _14279_ (_05977_, _05962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor _14280_ (_05978_, _05977_, _05976_);
  and _14281_ (_05979_, _05965_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _14282_ (_05980_, _05954_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor _14283_ (_05981_, _05980_, _05979_);
  and _14284_ (_05982_, _05981_, _05978_);
  and _14285_ (_05983_, _05982_, _05975_);
  and _14286_ (_05984_, _05983_, _05848_);
  nand _14287_ (_05985_, _05984_, _05971_);
  and _14288_ (_05986_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _14289_ (_05987_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _05850_);
  nand _14290_ (_05988_, _05987_, _05986_);
  and _14291_ (_05989_, _05988_, _05110_);
  and _14292_ (_07918_, _05989_, _05985_);
  and _14293_ (_05990_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _05110_);
  and _14294_ (_08055_, _05990_, _05986_);
  and _14295_ (_08294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _05110_);
  and _14296_ (_05991_, _05401_, _05389_);
  and _14297_ (_05992_, _05991_, _05376_);
  and _14298_ (_05993_, _05802_, _05461_);
  and _14299_ (_05994_, _05993_, _05992_);
  not _14300_ (_05995_, _05337_);
  and _14301_ (_05996_, _05991_, _05912_);
  and _14302_ (_05997_, _05993_, _05996_);
  nor _14303_ (_05998_, _05997_, _05994_);
  and _14304_ (_05999_, _05992_, _05462_);
  not _14305_ (_06000_, _05999_);
  and _14306_ (_06001_, _05913_, _05993_);
  and _14307_ (_06002_, _05993_, _05403_);
  nor _14308_ (_06003_, _06002_, _06001_);
  and _14309_ (_06004_, _06003_, _06000_);
  and _14310_ (_06005_, _06004_, _05998_);
  or _14311_ (_06006_, _06005_, _05995_);
  or _14312_ (_06007_, _06006_, _05994_);
  and _14313_ (_06008_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor _14314_ (_06009_, _05938_, _06000_);
  not _14315_ (_06010_, _05997_);
  nand _14316_ (_06011_, _06003_, _06010_);
  and _14317_ (_06012_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  or _14318_ (_06014_, _06012_, _06009_);
  and _14319_ (_06015_, _06014_, _05337_);
  or _14320_ (_06016_, _06015_, _06008_);
  and _14321_ (_08933_, _06016_, _05110_);
  not _14322_ (_06017_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _14323_ (_06018_, _06017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not _14324_ (_06019_, _05906_);
  or _14325_ (_06020_, _06019_, _05858_);
  or _14326_ (_06021_, _06020_, _05854_);
  and _14327_ (_06022_, _06021_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _14328_ (_06023_, _06022_, _06018_);
  nor _14329_ (_06024_, _05401_, _05389_);
  and _14330_ (_06025_, _06024_, _05912_);
  and _14331_ (_06026_, _06025_, _05804_);
  and _14332_ (_06027_, _06026_, _05794_);
  or _14333_ (_06028_, _06027_, _06023_);
  and _14334_ (_06029_, _06028_, _05844_);
  nand _14335_ (_06030_, _06027_, _05872_);
  and _14336_ (_06031_, _06030_, _06029_);
  nor _14337_ (_06032_, _05597_, _05187_);
  nor _14338_ (_06033_, _05603_, _05188_);
  or _14339_ (_06034_, _06033_, _06032_);
  and _14340_ (_06035_, _06034_, _05320_);
  nand _14341_ (_06036_, _05817_, _05285_);
  and _14342_ (_06037_, _06036_, _05319_);
  or _14343_ (_06038_, _06037_, _05658_);
  nand _14344_ (_06040_, _06037_, _05658_);
  and _14345_ (_06041_, _06040_, _05291_);
  and _14346_ (_06042_, _06041_, _06038_);
  nor _14347_ (_06043_, _06042_, _06035_);
  nor _14348_ (_06044_, _05597_, _05176_);
  not _14349_ (_06045_, _06044_);
  and _14350_ (_06046_, _05606_, _05295_);
  nor _14351_ (_06047_, _05604_, _05327_);
  nor _14352_ (_06048_, _06047_, _06046_);
  and _14353_ (_06049_, _05605_, _05312_);
  and _14354_ (_06050_, _05597_, _05314_);
  nor _14355_ (_06051_, _06050_, _06049_);
  and _14356_ (_06052_, _06051_, _06048_);
  and _14357_ (_06053_, _06052_, _06045_);
  and _14358_ (_06054_, _06053_, _06043_);
  nor _14359_ (_06055_, _06054_, _05844_);
  or _14360_ (_06056_, _06055_, _06031_);
  and _14361_ (_08980_, _06056_, _05110_);
  and _14362_ (_06057_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _14363_ (_06058_, _06020_, _05905_);
  and _14364_ (_06059_, _06058_, _06057_);
  and _14365_ (_06061_, _05866_, _05402_);
  and _14366_ (_06062_, _06061_, _05804_);
  and _14367_ (_06063_, _06062_, _05794_);
  or _14368_ (_06064_, _06063_, _06059_);
  and _14369_ (_06065_, _06064_, _05844_);
  nand _14370_ (_06066_, _06063_, _05872_);
  and _14371_ (_06067_, _06066_, _06065_);
  nor _14372_ (_06068_, _05210_, _05176_);
  not _14373_ (_06069_, _06068_);
  nand _14374_ (_06070_, _05276_, _05187_);
  nand _14375_ (_06071_, _05283_, _05188_);
  and _14376_ (_06072_, _06071_, _06070_);
  or _14377_ (_06073_, _06072_, _05211_);
  nand _14378_ (_06074_, _06072_, _05211_);
  and _14379_ (_06075_, _06074_, _05291_);
  nand _14380_ (_06076_, _06075_, _06073_);
  nand _14381_ (_06077_, _05529_, _05295_);
  or _14382_ (_06078_, _05528_, _05327_);
  and _14383_ (_06079_, _05527_, _05312_);
  not _14384_ (_06080_, _06079_);
  nor _14385_ (_06081_, _05526_, _05321_);
  and _14386_ (_06082_, _05314_, _05210_);
  nor _14387_ (_06083_, _06082_, _06081_);
  and _14388_ (_06084_, _06083_, _06080_);
  and _14389_ (_06085_, _06084_, _06078_);
  and _14390_ (_06086_, _06085_, _06077_);
  and _14391_ (_06087_, _06086_, _06076_);
  and _14392_ (_06088_, _06087_, _06069_);
  nor _14393_ (_06089_, _06088_, _05844_);
  or _14394_ (_06091_, _06089_, _06067_);
  and _14395_ (_09243_, _06091_, _05110_);
  nor _14396_ (_06092_, _05986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _14397_ (_06093_, _06092_);
  and _14398_ (_06094_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _05850_);
  and _14399_ (_06095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _14400_ (_06096_, _06095_, _06094_);
  and _14401_ (_06097_, _06096_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor _14402_ (_06098_, _06097_, _05848_);
  nor _14403_ (_06099_, _06098_, _05983_);
  nor _14404_ (_06100_, _06099_, _05971_);
  not _14405_ (_06101_, _06100_);
  or _14406_ (_06102_, _06101_, _05968_);
  not _14407_ (_06103_, _05976_);
  nor _14408_ (_06104_, _05979_, _05977_);
  and _14409_ (_06105_, _06104_, _06103_);
  or _14410_ (_06106_, _06098_, _06105_);
  and _14411_ (_06107_, _06106_, _06102_);
  or _14412_ (_06108_, _06107_, _06093_);
  not _14413_ (_06109_, _05952_);
  and _14414_ (_06110_, _06109_, _05941_);
  and _14415_ (_06111_, _05955_, _05941_);
  or _14416_ (_06112_, _06111_, _06110_);
  or _14417_ (_06113_, _06112_, _06099_);
  not _14418_ (_06114_, _05980_);
  and _14419_ (_06115_, _06114_, _05975_);
  nand _14420_ (_06116_, _06099_, _06115_);
  and _14421_ (_06117_, _06116_, _06113_);
  and _14422_ (_06118_, _06117_, _06092_);
  or _14423_ (_06119_, _06118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _14424_ (_06120_, _06119_, _05110_);
  and _14425_ (_10256_, _06120_, _06108_);
  not _14426_ (_06121_, _05433_);
  and _14427_ (_06122_, _05447_, _06121_);
  and _14428_ (_06123_, _06122_, _05797_);
  and _14429_ (_06124_, _06123_, _05867_);
  nand _14430_ (_06125_, _06124_, _05872_);
  or _14431_ (_06126_, _06124_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _14432_ (_06127_, _06121_, _05418_);
  and _14433_ (_06128_, _06127_, _05803_);
  and _14434_ (_06129_, _06128_, _05808_);
  not _14435_ (_06130_, _06129_);
  and _14436_ (_06131_, _06130_, _06126_);
  and _14437_ (_06132_, _06131_, _06125_);
  nor _14438_ (_06134_, _06130_, _05901_);
  or _14439_ (_06135_, _06134_, _06132_);
  and _14440_ (_10306_, _06135_, _05110_);
  and _14441_ (_06136_, _05986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not _14442_ (_06137_, _05986_);
  and _14443_ (_06138_, _06107_, _06137_);
  or _14444_ (_06139_, _06138_, _06092_);
  and _14445_ (_06140_, _06117_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _14446_ (_06141_, _06140_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _14447_ (_06142_, _06141_, _06139_);
  or _14448_ (_06143_, _06142_, _06136_);
  and _14449_ (_10385_, _06143_, _05110_);
  nor _14450_ (_06144_, _05433_, _05418_);
  and _14451_ (_06145_, _06144_, _05803_);
  and _14452_ (_06146_, _05806_, _05389_);
  and _14453_ (_06147_, _06146_, _05867_);
  and _14454_ (_06148_, _06147_, _06145_);
  not _14455_ (_06149_, _06148_);
  and _14456_ (_06150_, _05794_, _05460_);
  nor _14457_ (_06151_, _05418_, _05389_);
  and _14458_ (_06152_, _06151_, _06150_);
  and _14459_ (_06153_, _06152_, _06122_);
  and _14460_ (_06154_, _06153_, _05867_);
  or _14461_ (_06155_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _14462_ (_06156_, _06155_, _06149_);
  nand _14463_ (_06157_, _06154_, _05872_);
  and _14464_ (_06158_, _06157_, _06156_);
  nor _14465_ (_06159_, _06149_, _05901_);
  or _14466_ (_06160_, _06159_, _06158_);
  and _14467_ (_10406_, _06160_, _05110_);
  or _14468_ (_06161_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not _14469_ (_06162_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand _14470_ (_06163_, pc_log_change, _06162_);
  and _14471_ (_06164_, _06163_, _05110_);
  and _14472_ (_10427_, _06164_, _06161_);
  and _14473_ (_06165_, _05913_, _05462_);
  not _14474_ (_06166_, _06165_);
  nor _14475_ (_06167_, _06166_, _05334_);
  not _14476_ (_06168_, _05463_);
  and _14477_ (_06169_, _05996_, _05462_);
  nor _14478_ (_06170_, _05999_, _06169_);
  and _14479_ (_06171_, _06170_, _06168_);
  and _14480_ (_06172_, _06171_, _06166_);
  and _14481_ (_06173_, _05401_, _05365_);
  and _14482_ (_06174_, _05993_, _06173_);
  or _14483_ (_06175_, _06174_, _05995_);
  nor _14484_ (_06176_, _06175_, _06172_);
  nand _14485_ (_06177_, _06176_, _06171_);
  and _14486_ (_06178_, _06177_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or _14487_ (_06179_, _06178_, _06167_);
  or _14488_ (_06180_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and _14489_ (_06182_, _06180_, _05110_);
  and _14490_ (_12614_, _06182_, _06179_);
  not _14491_ (_06183_, _06054_);
  and _14492_ (_06184_, _06165_, _05337_);
  and _14493_ (_06185_, _06184_, _06183_);
  or _14494_ (_06186_, _06172_, _05995_);
  and _14495_ (_06187_, _06186_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nand _14496_ (_06188_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _14497_ (_06189_, _06188_, _06171_);
  or _14498_ (_06190_, _06189_, _06187_);
  or _14499_ (_06191_, _06190_, _06185_);
  and _14500_ (_12886_, _06191_, _05110_);
  and _14501_ (_06193_, _06186_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  not _14502_ (_06194_, _06088_);
  and _14503_ (_06195_, _06184_, _06194_);
  nand _14504_ (_06196_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _14505_ (_06197_, _06196_, _06171_);
  or _14506_ (_06198_, _06197_, _06195_);
  or _14507_ (_06199_, _06198_, _06193_);
  and _14508_ (_12945_, _06199_, _05110_);
  not _14509_ (_06200_, _05474_);
  not _14510_ (_06201_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _14511_ (_06202_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _14512_ (_06203_, _06202_, _06201_);
  nor _14513_ (_06204_, _06203_, _06200_);
  nor _14514_ (_06205_, _06204_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _14515_ (_06206_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  not _14516_ (_06207_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand _14517_ (_06208_, _06205_, _06207_);
  and _14518_ (_06209_, _06208_, _05110_);
  and _14519_ (_13108_, _06209_, _06206_);
  and _14520_ (_06210_, _06186_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or _14521_ (_06211_, _05282_, _05187_);
  or _14522_ (_06212_, _05275_, _05188_);
  and _14523_ (_06213_, _06212_, _06211_);
  or _14524_ (_06214_, _06213_, _05279_);
  nand _14525_ (_06215_, _06213_, _05279_);
  and _14526_ (_06216_, _06215_, _05291_);
  and _14527_ (_06217_, _06216_, _06214_);
  nor _14528_ (_06218_, _05534_, _05321_);
  nor _14529_ (_06219_, _06218_, _06217_);
  and _14530_ (_06220_, _05535_, _05312_);
  and _14531_ (_06221_, _05314_, _05233_);
  nor _14532_ (_06222_, _06221_, _06220_);
  nor _14533_ (_06223_, _05233_, _05176_);
  and _14534_ (_06224_, _05538_, _05295_);
  nor _14535_ (_06225_, _05537_, _05327_);
  or _14536_ (_06226_, _06225_, _06224_);
  nor _14537_ (_06227_, _06226_, _06223_);
  and _14538_ (_06228_, _06227_, _06222_);
  and _14539_ (_06229_, _06228_, _06219_);
  not _14540_ (_06230_, _06229_);
  and _14541_ (_06231_, _06230_, _06184_);
  nand _14542_ (_06232_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _14543_ (_06233_, _06232_, _06171_);
  or _14544_ (_06234_, _06233_, _06231_);
  or _14545_ (_06235_, _06234_, _06210_);
  and _14546_ (_13173_, _06235_, _05110_);
  and _14547_ (_06237_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _14548_ (_06238_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _14549_ (_06239_, \oc8051_top_1.oc8051_decoder1.state [0], _05151_);
  and _14550_ (_06240_, _06239_, _06238_);
  not _14551_ (_06241_, _05475_);
  nor _14552_ (_06242_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _14553_ (_06243_, _06242_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _14554_ (_06244_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _14555_ (_06245_, _06202_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _14556_ (_06246_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and _14557_ (_06247_, _06246_, _06244_);
  not _14558_ (_06248_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  not _14559_ (_06249_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _14560_ (_06250_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _06201_);
  nand _14561_ (_06251_, _06250_, _06249_);
  or _14562_ (_06252_, _06251_, _06248_);
  and _14563_ (_06253_, _06252_, _06247_);
  not _14564_ (_06254_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _14565_ (_06255_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _14566_ (_06256_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], _06255_);
  and _14567_ (_06257_, _06256_, _06201_);
  nand _14568_ (_06258_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _14569_ (_06259_, _06258_, _06254_);
  nor _14570_ (_06260_, _06242_, _06201_);
  nand _14571_ (_06261_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _14572_ (_06262_, _06242_, _06201_);
  nand _14573_ (_06263_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and _14574_ (_06264_, _06263_, _06261_);
  and _14575_ (_06265_, _06264_, _06259_);
  nand _14576_ (_06266_, _06265_, _06253_);
  or _14577_ (_06267_, _06266_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14578_ (_06268_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _14579_ (_06269_, _06268_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  not _14580_ (_06270_, _06269_);
  and _14581_ (_06271_, _06270_, _06267_);
  or _14582_ (_06272_, _06271_, _06241_);
  not _14583_ (_06273_, _05472_);
  nor _14584_ (_06274_, _05474_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _14585_ (_06275_, _06274_, _06273_);
  and _14586_ (_06276_, _06275_, _06272_);
  not _14587_ (_06277_, _06276_);
  nand _14588_ (_06278_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _14589_ (_06279_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _14590_ (_06280_, _06279_, _06278_);
  nand _14591_ (_06281_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand _14592_ (_06282_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and _14593_ (_06283_, _06282_, _06281_);
  nand _14594_ (_06284_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  not _14595_ (_06285_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _14596_ (_06286_, _06251_, _06285_);
  and _14597_ (_06287_, _06286_, _06284_);
  and _14598_ (_06288_, _06287_, _06283_);
  and _14599_ (_06289_, _06288_, _06280_);
  or _14600_ (_06290_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _14601_ (_06291_, _06290_, _06289_);
  and _14602_ (_06292_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  not _14603_ (_06293_, _06292_);
  and _14604_ (_06294_, _06293_, _06291_);
  nand _14605_ (_06295_, _06294_, _05475_);
  nor _14606_ (_06296_, _05474_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _14607_ (_06297_, _06296_, _06273_);
  and _14608_ (_06298_, _06297_, _06295_);
  nand _14609_ (_06300_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand _14610_ (_06301_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _14611_ (_06302_, _06301_, _06300_);
  nand _14612_ (_06303_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand _14613_ (_06304_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _14614_ (_06305_, _06304_, _06303_);
  nand _14615_ (_06306_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  not _14616_ (_06307_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _14617_ (_06308_, _06251_, _06307_);
  and _14618_ (_06309_, _06308_, _06306_);
  and _14619_ (_06310_, _06309_, _06305_);
  and _14620_ (_06311_, _06310_, _06302_);
  or _14621_ (_06312_, _06311_, _06290_);
  and _14622_ (_06313_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _14623_ (_06314_, _06313_);
  and _14624_ (_06315_, _06314_, _06312_);
  nand _14625_ (_06316_, _06315_, _05475_);
  nor _14626_ (_06317_, _05474_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _14627_ (_06318_, _06317_, _06273_);
  and _14628_ (_06319_, _06318_, _06316_);
  not _14629_ (_06320_, _06319_);
  and _14630_ (_06321_, _06320_, _06298_);
  nor _14631_ (_06322_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _14632_ (_06323_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand _14633_ (_06324_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _14634_ (_06325_, _06324_, _06323_);
  nand _14635_ (_06326_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand _14636_ (_06327_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and _14637_ (_06328_, _06327_, _06326_);
  nand _14638_ (_06329_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  not _14639_ (_06330_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or _14640_ (_06331_, _06251_, _06330_);
  and _14641_ (_06332_, _06331_, _06329_);
  and _14642_ (_06333_, _06332_, _06328_);
  nand _14643_ (_06334_, _06333_, _06325_);
  nand _14644_ (_06335_, _06334_, _06322_);
  and _14645_ (_06336_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  not _14646_ (_06337_, _06336_);
  and _14647_ (_06338_, _06337_, _06335_);
  nand _14648_ (_06339_, _06338_, _05475_);
  nor _14649_ (_06340_, _05474_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _14650_ (_06341_, _06340_, _06273_);
  and _14651_ (_06342_, _06341_, _06339_);
  and _14652_ (_06343_, _06342_, _06321_);
  and _14653_ (_06344_, _06343_, _06277_);
  nand _14654_ (_06345_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nand _14655_ (_06346_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _14656_ (_06347_, _06346_, _06345_);
  nand _14657_ (_06348_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand _14658_ (_06349_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and _14659_ (_06350_, _06349_, _06348_);
  nand _14660_ (_06351_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  not _14661_ (_06352_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _14662_ (_06353_, _06251_, _06352_);
  and _14663_ (_06354_, _06353_, _06351_);
  and _14664_ (_06355_, _06354_, _06350_);
  nand _14665_ (_06356_, _06355_, _06347_);
  nand _14666_ (_06357_, _06356_, _06254_);
  nand _14667_ (_06358_, _06357_, _06268_);
  nor _14668_ (_06359_, _06268_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  not _14669_ (_06360_, _06359_);
  and _14670_ (_06362_, _06360_, _06358_);
  or _14671_ (_06363_, _06362_, _06241_);
  nor _14672_ (_06364_, _05474_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _14673_ (_06365_, _06364_, _06273_);
  and _14674_ (_06366_, _06365_, _06363_);
  nand _14675_ (_06367_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand _14676_ (_06368_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and _14677_ (_06369_, _06368_, _06367_);
  not _14678_ (_06370_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _14679_ (_06371_, _06251_, _06370_);
  and _14680_ (_06373_, _06371_, _06369_);
  nand _14681_ (_06374_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _14682_ (_06375_, _06374_, _06254_);
  nand _14683_ (_06376_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand _14684_ (_06377_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _14685_ (_06378_, _06377_, _06376_);
  and _14686_ (_06379_, _06378_, _06375_);
  nand _14687_ (_06380_, _06379_, _06373_);
  or _14688_ (_06381_, _06380_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _14689_ (_06382_, _06268_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  not _14690_ (_06383_, _06382_);
  and _14691_ (_06384_, _06383_, _06381_);
  or _14692_ (_06385_, _06384_, _06241_);
  nor _14693_ (_06386_, _05474_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _14694_ (_06387_, _06386_, _06273_);
  and _14695_ (_06388_, _06387_, _06385_);
  nor _14696_ (_06389_, _06388_, _06366_);
  nand _14697_ (_06390_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nand _14698_ (_06391_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _14699_ (_06392_, _06391_, _06390_);
  nand _14700_ (_06393_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand _14701_ (_06394_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _14702_ (_06395_, _06394_, _06393_);
  nand _14703_ (_06396_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  not _14704_ (_06397_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _14705_ (_06398_, _06251_, _06397_);
  and _14706_ (_06399_, _06398_, _06396_);
  and _14707_ (_06400_, _06399_, _06395_);
  nand _14708_ (_06401_, _06400_, _06392_);
  nand _14709_ (_06402_, _06401_, _06254_);
  nand _14710_ (_06403_, _06402_, _06268_);
  nor _14711_ (_06404_, _06268_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  not _14712_ (_06405_, _06404_);
  and _14713_ (_06406_, _06405_, _06403_);
  or _14714_ (_06407_, _06406_, _06241_);
  nor _14715_ (_06409_, _05474_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _14716_ (_06410_, _06409_, _06273_);
  and _14717_ (_06411_, _06410_, _06407_);
  nand _14718_ (_06412_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  not _14719_ (_06413_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _14720_ (_06414_, _06251_, _06413_);
  and _14721_ (_06415_, _06414_, _06412_);
  nand _14722_ (_06416_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nand _14723_ (_06417_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _14724_ (_06418_, _06417_, _06416_);
  nand _14725_ (_06419_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand _14726_ (_06420_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and _14727_ (_06421_, _06420_, _06419_);
  and _14728_ (_06422_, _06421_, _06418_);
  and _14729_ (_06423_, _06422_, _06415_);
  or _14730_ (_06424_, _06423_, _06290_);
  and _14731_ (_06425_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  not _14732_ (_06426_, _06425_);
  and _14733_ (_06427_, _06426_, _06424_);
  nand _14734_ (_06428_, _06427_, _05475_);
  nor _14735_ (_06429_, _05474_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _14736_ (_06430_, _06429_, _06273_);
  and _14737_ (_06431_, _06430_, _06428_);
  not _14738_ (_06432_, _06431_);
  and _14739_ (_06433_, _06432_, _06411_);
  and _14740_ (_06434_, _06433_, _06389_);
  and _14741_ (_06435_, _06434_, _06344_);
  not _14742_ (_06436_, _06342_);
  and _14743_ (_06437_, _06436_, _06321_);
  and _14744_ (_06438_, _06437_, _06277_);
  and _14745_ (_06439_, _06438_, _06434_);
  nor _14746_ (_06440_, _06439_, _06435_);
  not _14747_ (_06442_, _06440_);
  and _14748_ (_06443_, _06442_, _06240_);
  or _14749_ (_06444_, _06443_, _06237_);
  not _14750_ (_06445_, _06388_);
  nor _14751_ (_06446_, _06411_, _06445_);
  and _14752_ (_06447_, _06446_, _06432_);
  and _14753_ (_06448_, _06447_, _06366_);
  and _14754_ (_06449_, _06448_, _06344_);
  nor _14755_ (_06450_, _06431_, _06411_);
  and _14756_ (_06451_, _06450_, _06389_);
  and _14757_ (_06452_, _06437_, _06276_);
  and _14758_ (_06453_, _06452_, _06451_);
  or _14759_ (_06454_, _06453_, _06449_);
  nor _14760_ (_06455_, _06432_, _06276_);
  and _14761_ (_06456_, _06436_, _06319_);
  and _14762_ (_06457_, _06456_, _06455_);
  and _14763_ (_06458_, _06457_, _06298_);
  and _14764_ (_06459_, _06456_, _06298_);
  and _14765_ (_06460_, _06433_, _06388_);
  and _14766_ (_06461_, _06460_, _06459_);
  or _14767_ (_06462_, _06461_, _06458_);
  and _14768_ (_06463_, _06459_, _06277_);
  and _14769_ (_06464_, _06433_, _06445_);
  and _14770_ (_06465_, _06464_, _06463_);
  or _14771_ (_06466_, _06465_, _06462_);
  or _14772_ (_06467_, _06466_, _06454_);
  and _14773_ (_06468_, _06467_, _05474_);
  or _14774_ (_06469_, _06468_, _06444_);
  and _14775_ (_01001_, _06469_, _05110_);
  and _14776_ (_06470_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _05151_);
  and _14777_ (_06471_, _06470_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _14778_ (_06472_, _05785_, _05486_);
  and _14779_ (_06473_, _05804_, _06472_);
  and _14780_ (_06475_, _06473_, _06146_);
  nor _14781_ (_06476_, _06475_, _06471_);
  not _14782_ (_06477_, _06476_);
  or _14783_ (_06478_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nor _14784_ (_06479_, _05697_, _05696_);
  nor _14785_ (_06480_, _06479_, _05699_);
  nor _14786_ (_06481_, _06480_, _05651_);
  not _14787_ (_06482_, _06481_);
  or _14788_ (_06483_, _05233_, _05169_);
  and _14789_ (_06485_, _05157_, _05163_);
  and _14790_ (_06486_, _06485_, ABINPUT000000[2]);
  and _14791_ (_06487_, _05311_, _05154_);
  and _14792_ (_06488_, _06487_, ABINPUT000[2]);
  nor _14793_ (_06489_, _06488_, _06486_);
  and _14794_ (_06490_, _06489_, _06483_);
  and _14795_ (_06491_, _05281_, _05158_);
  and _14796_ (_06492_, _05280_, _05172_);
  nor _14797_ (_06493_, _06492_, _06491_);
  and _14798_ (_06494_, _06493_, _06490_);
  and _14799_ (_06495_, _06494_, _05934_);
  and _14800_ (_06496_, _06495_, _05930_);
  and _14801_ (_06497_, _06496_, _05926_);
  nor _14802_ (_06498_, _05728_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _14803_ (_06499_, _06498_, _05281_);
  nor _14804_ (_06500_, _06498_, _05281_);
  nor _14805_ (_06501_, _06500_, _06499_);
  nor _14806_ (_06502_, _06501_, _05737_);
  or _14807_ (_06503_, _05549_, _05253_);
  and _14808_ (_06504_, _05928_, _06503_);
  or _14809_ (_06505_, _06504_, _05555_);
  and _14810_ (_06506_, _06505_, _05564_);
  nor _14811_ (_06507_, _06505_, _05564_);
  or _14812_ (_06508_, _06507_, _06506_);
  and _14813_ (_06509_, _06508_, _05489_);
  nor _14814_ (_06510_, _06509_, _06502_);
  and _14815_ (_06511_, _06510_, _06497_);
  and _14816_ (_06512_, _06511_, _06482_);
  nand _14817_ (_06513_, _06512_, _06477_);
  and _14818_ (_06514_, _06513_, _05110_);
  and _14819_ (_01593_, _06514_, _06478_);
  nor _14820_ (_06515_, _05713_, _05674_);
  nor _14821_ (_06516_, _06515_, _05714_);
  nor _14822_ (_06517_, _06516_, _05651_);
  not _14823_ (_06518_, _06517_);
  nor _14824_ (_06519_, _05606_, _05307_);
  or _14825_ (_06520_, _06519_, _05638_);
  and _14826_ (_06521_, _06520_, _05576_);
  nor _14827_ (_06522_, _06521_, _05490_);
  and _14828_ (_06523_, _06522_, _05608_);
  nor _14829_ (_06524_, _05597_, _05159_);
  and _14830_ (_06525_, _06485_, ABINPUT000000[6]);
  nor _14831_ (_06526_, _06525_, _06524_);
  and _14832_ (_06528_, _06526_, _06052_);
  nor _14833_ (_06529_, _05720_, _05510_);
  nor _14834_ (_06530_, _06529_, _05187_);
  and _14835_ (_06531_, _06530_, _05743_);
  nor _14836_ (_06532_, _06531_, _05731_);
  and _14837_ (_06533_, _06532_, _05597_);
  nor _14838_ (_06534_, _06532_, _05597_);
  nor _14839_ (_06535_, _06534_, _06533_);
  nor _14840_ (_06536_, _06535_, _05737_);
  nor _14841_ (_06537_, _05174_, _05150_);
  or _14842_ (_06538_, _05627_, _05169_);
  and _14843_ (_06539_, _06487_, ABINPUT000[6]);
  not _14844_ (_06540_, _06539_);
  nand _14845_ (_06541_, _06540_, _06538_);
  or _14846_ (_06542_, _06541_, _06537_);
  nor _14847_ (_06543_, _06542_, _06536_);
  and _14848_ (_06544_, _06543_, _06528_);
  and _14849_ (_06545_, _06544_, _06043_);
  not _14850_ (_06546_, _06545_);
  nor _14851_ (_06547_, _06546_, _06523_);
  and _14852_ (_06548_, _06547_, _06518_);
  nand _14853_ (_06549_, _06548_, _06477_);
  or _14854_ (_06550_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _14855_ (_06551_, _06550_, _05110_);
  and _14856_ (_01615_, _06551_, _06549_);
  not _14857_ (_06552_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  not _14858_ (_06553_, _06002_);
  and _14859_ (_06554_, _06553_, _05998_);
  nor _14860_ (_06555_, _06554_, _05995_);
  nor _14861_ (_06556_, _06555_, _06552_);
  nand _14862_ (_06557_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _14863_ (_06558_, _06557_, _05998_);
  not _14864_ (_06559_, _05938_);
  and _14865_ (_06560_, _06002_, _05337_);
  and _14866_ (_06561_, _06560_, _06559_);
  or _14867_ (_06562_, _06561_, _06558_);
  or _14868_ (_06563_, _06562_, _06556_);
  and _14869_ (_03222_, _06563_, _05110_);
  nand _14870_ (_06564_, _05647_, _05519_);
  nor _14871_ (_06565_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _14872_ (_06566_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05240_);
  nor _14873_ (_06567_, _06566_, _06565_);
  and _14874_ (_06568_, _06567_, _06564_);
  nor _14875_ (_06569_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _14876_ (_06570_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05264_);
  nor _14877_ (_06571_, _06570_, _06569_);
  and _14878_ (_06572_, _06571_, _06568_);
  nor _14879_ (_06573_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _14880_ (_06574_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05218_);
  nor _14881_ (_06575_, _06574_, _06573_);
  and _14882_ (_06576_, _06575_, _06572_);
  nor _14883_ (_06577_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _14884_ (_06578_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05195_);
  nor _14885_ (_06579_, _06578_, _06577_);
  or _14886_ (_06580_, _06579_, _06576_);
  nand _14887_ (_06581_, _06579_, _06576_);
  and _14888_ (_06582_, _06581_, _05489_);
  nand _14889_ (_06583_, _06582_, _06580_);
  and _14890_ (_06584_, _05877_, _05510_);
  and _14891_ (_06585_, _06584_, _05549_);
  and _14892_ (_06586_, _06585_, _05552_);
  and _14893_ (_06587_, _05534_, _05187_);
  and _14894_ (_06588_, _06587_, _06586_);
  nor _14895_ (_06589_, _05549_, _05510_);
  and _14896_ (_06590_, _06589_, _05875_);
  and _14897_ (_06591_, _06590_, _05543_);
  nor _14898_ (_06592_, _05534_, _05187_);
  and _14899_ (_06593_, _06592_, _06591_);
  nor _14900_ (_06594_, _06593_, _06588_);
  and _14901_ (_06595_, _06594_, _05526_);
  not _14902_ (_06596_, _06595_);
  nor _14903_ (_06597_, _06594_, _05526_);
  nor _14904_ (_06598_, _06597_, _05882_);
  and _14905_ (_06599_, _06598_, _06596_);
  and _14906_ (_06600_, _06485_, ABINPUT000000[12]);
  and _14907_ (_06601_, _06487_, ABINPUT000[12]);
  nor _14908_ (_06602_, _06601_, _06600_);
  nor _14909_ (_06603_, _05321_, _05210_);
  nor _14910_ (_06604_, _05526_, _05159_);
  or _14911_ (_06605_, _06604_, _06603_);
  nor _14912_ (_06606_, _06605_, _05764_);
  and _14913_ (_06607_, _06606_, _06602_);
  not _14914_ (_06608_, _06607_);
  nor _14915_ (_06609_, _06608_, _06599_);
  nand _14916_ (_06610_, _06609_, _06583_);
  not _14917_ (_06611_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _14918_ (_06612_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05151_);
  and _14919_ (_06613_, _06612_, _06611_);
  nand _14920_ (_06615_, _06613_, _06610_);
  not _14921_ (_06616_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _14922_ (_06617_, _06470_, _06616_);
  and _14923_ (_06618_, _05460_, _05448_);
  and _14924_ (_06619_, _06618_, _06127_);
  and _14925_ (_06620_, _06619_, _05992_);
  and _14926_ (_06621_, _06620_, _05806_);
  nor _14927_ (_06622_, _06621_, _06617_);
  not _14928_ (_06623_, _06622_);
  and _14929_ (_06624_, _05460_, _05389_);
  and _14930_ (_06625_, _06624_, _05418_);
  nor _14931_ (_06626_, _05447_, _05433_);
  and _14932_ (_06627_, _06626_, _05794_);
  and _14933_ (_06628_, _06627_, _06625_);
  nor _14934_ (_06629_, _06628_, _05204_);
  nor _14935_ (_06630_, _06629_, _06623_);
  and _14936_ (_06631_, _05866_, _05401_);
  and _14937_ (_06632_, _06631_, _05782_);
  nor _14938_ (_06633_, _06631_, _05204_);
  or _14939_ (_06634_, _06633_, _06632_);
  nand _14940_ (_06635_, _06634_, _06628_);
  and _14941_ (_06636_, _06635_, _06630_);
  not _14942_ (_06637_, _06613_);
  and _14943_ (_06638_, _06622_, _06637_);
  nor _14944_ (_06639_, _05700_, _05687_);
  nor _14945_ (_06640_, _06639_, _05702_);
  nor _14946_ (_06641_, _06640_, _05651_);
  not _14947_ (_06642_, _06641_);
  nor _14948_ (_06643_, _05570_, _05561_);
  or _14949_ (_06644_, _06643_, _05490_);
  nor _14950_ (_06645_, _06644_, _05571_);
  not _14951_ (_06646_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _14952_ (_06647_, _05726_, _06646_);
  nor _14953_ (_06648_, _06647_, _05211_);
  nor _14954_ (_06649_, _05728_, _05737_);
  not _14955_ (_06650_, _06649_);
  nor _14956_ (_06651_, _06650_, _06648_);
  nor _14957_ (_06652_, _05233_, _05174_);
  and _14958_ (_06653_, _06485_, ABINPUT000000[4]);
  and _14959_ (_06654_, _06487_, ABINPUT000[4]);
  nor _14960_ (_06655_, _06654_, _06653_);
  not _14961_ (_06656_, _06655_);
  nor _14962_ (_06657_, _06656_, _06652_);
  or _14963_ (_06658_, _05169_, _05150_);
  nor _14964_ (_06659_, _05210_, _05159_);
  not _14965_ (_06660_, _06659_);
  and _14966_ (_06661_, _06660_, _06658_);
  and _14967_ (_06662_, _06661_, _06657_);
  not _14968_ (_06663_, _06662_);
  nor _14969_ (_06664_, _06663_, _06651_);
  and _14970_ (_06665_, _06664_, _06087_);
  not _14971_ (_06666_, _06665_);
  nor _14972_ (_06667_, _06666_, _06645_);
  and _14973_ (_06668_, _06667_, _06642_);
  nor _14974_ (_06669_, _06668_, _06613_);
  nor _14975_ (_06670_, _06669_, _06638_);
  or _14976_ (_06671_, _06670_, _06636_);
  nand _14977_ (_06672_, _06671_, _06615_);
  and _14978_ (_03832_, _06672_, _05110_);
  and _14979_ (_06673_, _05994_, _05337_);
  nand _14980_ (_06674_, _06673_, _06088_);
  or _14981_ (_06675_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _14982_ (_06676_, _06675_, _05110_);
  and _14983_ (_03950_, _06676_, _06674_);
  nand _14984_ (_06677_, _06673_, _06054_);
  or _14985_ (_06678_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _14986_ (_06679_, _06678_, _05110_);
  and _14987_ (_04296_, _06679_, _06677_);
  nor _14988_ (_06680_, _06010_, _05334_);
  and _14989_ (_06681_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _14990_ (_06682_, _06681_, _05995_);
  or _14991_ (_06683_, _06682_, _06680_);
  or _14992_ (_06685_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _14993_ (_06686_, _06685_, _05110_);
  and _14994_ (_04377_, _06686_, _06683_);
  nand _14995_ (_06687_, _06673_, _05334_);
  or _14996_ (_06688_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _14997_ (_06689_, _06688_, _05110_);
  and _14998_ (_05107_, _06689_, _06687_);
  nand _14999_ (_06690_, _06560_, _06229_);
  or _15000_ (_06691_, _06560_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _15001_ (_06692_, _06691_, _05110_);
  and _15002_ (_05108_, _06692_, _06690_);
  and _15003_ (_06693_, _06579_, _06576_);
  nor _15004_ (_06694_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15005_ (_06695_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05581_);
  nor _15006_ (_06696_, _06695_, _06694_);
  nor _15007_ (_06697_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15008_ (_06698_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05123_);
  nor _15009_ (_06699_, _06698_, _06697_);
  and _15010_ (_06700_, _06699_, _06696_);
  and _15011_ (_06701_, _06700_, _06693_);
  nor _15012_ (_06702_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _15013_ (_06703_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05613_);
  nor _15014_ (_06704_, _06703_, _06702_);
  or _15015_ (_06705_, _06704_, _06701_);
  nand _15016_ (_06706_, _06704_, _06701_);
  and _15017_ (_06707_, _06706_, _05489_);
  nand _15018_ (_06708_, _06707_, _06705_);
  not _15019_ (_06709_, _05510_);
  and _15020_ (_06710_, _05875_, _06709_);
  and _15021_ (_06711_, _06710_, _05550_);
  and _15022_ (_06712_, _06711_, _05543_);
  and _15023_ (_06713_, _06712_, _05682_);
  and _15024_ (_06714_, _06713_, _05703_);
  and _15025_ (_06716_, _06714_, _05661_);
  nor _15026_ (_06717_, _06716_, _05187_);
  and _15027_ (_06718_, _06586_, _05534_);
  and _15028_ (_06719_, _06718_, _05526_);
  and _15029_ (_06720_, _06719_, _05306_);
  nor _15030_ (_06721_, _06720_, _05188_);
  or _15031_ (_06722_, _06721_, _06717_);
  and _15032_ (_06723_, _05603_, _05188_);
  nor _15033_ (_06724_, _06723_, _06033_);
  not _15034_ (_06725_, _06724_);
  nor _15035_ (_06726_, _06725_, _06722_);
  and _15036_ (_06727_, _06726_, _05655_);
  or _15037_ (_06728_, _06726_, _05655_);
  nand _15038_ (_06729_, _06728_, _05291_);
  or _15039_ (_06730_, _06729_, _06727_);
  and _15040_ (_06731_, _06487_, ABINPUT000[15]);
  and _15041_ (_06732_, _05627_, _05187_);
  not _15042_ (_06733_, _06732_);
  and _15043_ (_06734_, _05633_, _05188_);
  nor _15044_ (_06735_, _06734_, _05321_);
  and _15045_ (_06736_, _06735_, _06733_);
  nor _15046_ (_06737_, _05233_, _05763_);
  nor _15047_ (_06738_, _05633_, _05159_);
  and _15048_ (_06739_, _06485_, ABINPUT000000[15]);
  or _15049_ (_06740_, _06739_, _06738_);
  or _15050_ (_06741_, _06740_, _06737_);
  or _15051_ (_06742_, _06741_, _06736_);
  nor _15052_ (_06743_, _06742_, _06731_);
  and _15053_ (_06744_, _06743_, _06730_);
  nand _15054_ (_06745_, _06744_, _06708_);
  and _15055_ (_06746_, _06745_, _06613_);
  and _15056_ (_06747_, _06628_, _05488_);
  nor _15057_ (_06748_, _06747_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  not _15058_ (_06749_, _06748_);
  and _15059_ (_06750_, _06749_, _06638_);
  nand _15060_ (_06751_, _06747_, _05872_);
  and _15061_ (_06752_, _06751_, _06750_);
  and _15062_ (_06753_, _05643_, _05608_);
  not _15063_ (_06754_, _06753_);
  and _15064_ (_06755_, _05644_, _05489_);
  and _15065_ (_06756_, _06755_, _06754_);
  not _15066_ (_06757_, _06756_);
  nor _15067_ (_06758_, _05714_, _05671_);
  nor _15068_ (_06759_, _06758_, _05715_);
  nor _15069_ (_06760_, _06759_, _05651_);
  nor _15070_ (_06761_, _06533_, _05627_);
  and _15071_ (_06762_, _06533_, _05627_);
  nor _15072_ (_06763_, _06762_, _06761_);
  nor _15073_ (_06764_, _06763_, _05737_);
  or _15074_ (_06765_, _05510_, _05169_);
  and _15075_ (_06766_, _06485_, ABINPUT000000[7]);
  and _15076_ (_06767_, _06487_, ABINPUT000[7]);
  nor _15077_ (_06768_, _06767_, _06766_);
  and _15078_ (_06769_, _06768_, _06765_);
  nor _15079_ (_06770_, _05627_, _05159_);
  nor _15080_ (_06771_, _05597_, _05174_);
  nor _15081_ (_06772_, _06771_, _06770_);
  and _15082_ (_06773_, _06772_, _06769_);
  and _15083_ (_06774_, _06773_, _05839_);
  not _15084_ (_06775_, _06774_);
  nor _15085_ (_06776_, _06775_, _06764_);
  and _15086_ (_06777_, _06776_, _05828_);
  not _15087_ (_06778_, _06777_);
  nor _15088_ (_06779_, _06778_, _06760_);
  and _15089_ (_06780_, _06779_, _06757_);
  nor _15090_ (_06781_, _06780_, _06622_);
  or _15091_ (_06783_, _06781_, _06752_);
  and _15092_ (_06784_, _06783_, _06637_);
  or _15093_ (_06785_, _06784_, _06746_);
  and _15094_ (_05109_, _06785_, _05110_);
  or _15095_ (_06786_, _05551_, _05756_);
  and _15096_ (_06787_, _06786_, _05327_);
  or _15097_ (_06788_, _06787_, _05562_);
  nand _15098_ (_06789_, _05551_, _05312_);
  or _15099_ (_06790_, _05932_, _05280_);
  and _15100_ (_06791_, _06790_, _06789_);
  or _15101_ (_06792_, _05549_, _05321_);
  or _15102_ (_06793_, _05882_, _05280_);
  and _15103_ (_06794_, _06793_, _06792_);
  or _15104_ (_06795_, _05253_, _05176_);
  and _15105_ (_06796_, _06795_, _06794_);
  and _15106_ (_06797_, _06796_, _06791_);
  and _15107_ (_06798_, _06797_, _06788_);
  not _15108_ (_06799_, _06798_);
  and _15109_ (_06800_, _06799_, _05463_);
  not _15110_ (_06801_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor _15111_ (_06802_, _05464_, _06801_);
  or _15112_ (_06803_, _06802_, _06800_);
  or _15113_ (_06804_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _15114_ (_06805_, _06804_, _05110_);
  and _15115_ (_05173_, _06805_, _06803_);
  and _15116_ (_06807_, \oc8051_top_1.oc8051_sfr1.wait_data , _05110_);
  and _15117_ (_06808_, _06807_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _15118_ (_06809_, _06445_, _06366_);
  and _15119_ (_06810_, _06809_, _06433_);
  and _15120_ (_06811_, _06459_, _06276_);
  and _15121_ (_06812_, _06811_, _06810_);
  nor _15122_ (_06813_, _06319_, _06298_);
  and _15123_ (_06814_, _06813_, _06436_);
  and _15124_ (_06815_, _06814_, _06277_);
  and _15125_ (_06816_, _06815_, _06434_);
  and _15126_ (_06817_, _06815_, _06810_);
  or _15127_ (_06818_, _06817_, _06816_);
  or _15128_ (_06819_, _06818_, _06812_);
  and _15129_ (_06820_, _06814_, _06276_);
  and _15130_ (_06821_, _06820_, _06464_);
  or _15131_ (_06822_, _06821_, _06819_);
  and _15132_ (_06823_, _06814_, _06460_);
  and _15133_ (_06824_, _06342_, _06276_);
  and _15134_ (_06825_, _06824_, _06321_);
  and _15135_ (_06826_, _06411_, _06388_);
  or _15136_ (_06827_, _06826_, _06431_);
  and _15137_ (_06828_, _06827_, _06825_);
  nor _15138_ (_06829_, _06828_, _06823_);
  and _15139_ (_06830_, _06431_, _06276_);
  or _15140_ (_06831_, _06814_, _06459_);
  and _15141_ (_06832_, _06831_, _06830_);
  and _15142_ (_06833_, _06814_, _06455_);
  nor _15143_ (_06834_, _06833_, _06832_);
  nand _15144_ (_06835_, _06834_, _06829_);
  and _15145_ (_06836_, _06825_, _06434_);
  and _15146_ (_06837_, _06452_, _06434_);
  or _15147_ (_06838_, _06837_, _06836_);
  or _15148_ (_06839_, _06838_, _06454_);
  or _15149_ (_06840_, _06839_, _06835_);
  or _15150_ (_06841_, _06840_, _06822_);
  and _15151_ (_06842_, _05474_, _05110_);
  and _15152_ (_06843_, _06842_, _06841_);
  or _15153_ (_05179_, _06843_, _06808_);
  and _15154_ (_06844_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _15155_ (_06845_, _06810_, _06438_);
  and _15156_ (_06846_, _06845_, _05474_);
  or _15157_ (_06847_, _06846_, _06844_);
  or _15158_ (_06848_, _06847_, _06443_);
  and _15159_ (_05205_, _06848_, _05110_);
  and _15160_ (_06849_, _06448_, _06437_);
  not _15161_ (_06850_, _06849_);
  and _15162_ (_06851_, _06342_, _06319_);
  and _15163_ (_06852_, _06851_, _06298_);
  and _15164_ (_06853_, _06852_, _06451_);
  and _15165_ (_06854_, _06853_, _06277_);
  and _15166_ (_06856_, _06852_, _06277_);
  and _15167_ (_06857_, _06856_, _06447_);
  nor _15168_ (_06858_, _06857_, _06854_);
  nand _15169_ (_06859_, _06858_, _06850_);
  and _15170_ (_06860_, _06859_, _06240_);
  or _15171_ (_06861_, _06860_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _15172_ (_06862_, _06448_, _06438_);
  nor _15173_ (_06863_, _06431_, _06366_);
  and _15174_ (_06864_, _06863_, _06446_);
  and _15175_ (_06865_, _06864_, _06820_);
  and _15176_ (_06866_, _06809_, _06450_);
  and _15177_ (_06867_, _06866_, _06276_);
  or _15178_ (_06868_, _06867_, _06865_);
  or _15179_ (_06869_, _06868_, _06862_);
  or _15180_ (_06870_, _05473_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _15181_ (_06871_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _15182_ (_06872_, \oc8051_top_1.oc8051_decoder1.state [1], _05151_);
  and _15183_ (_06873_, _06872_, _06871_);
  and _15184_ (_06874_, _06868_, _06873_);
  or _15185_ (_06875_, _06874_, _06870_);
  and _15186_ (_06876_, _06875_, _06869_);
  or _15187_ (_06877_, _06876_, _06861_);
  or _15188_ (_06878_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05151_);
  and _15189_ (_06879_, _06878_, _05110_);
  and _15190_ (_05208_, _06879_, _06877_);
  and _15191_ (_06880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _15192_ (_06881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _15193_ (_06882_, _06881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _15194_ (_06883_, _06882_, _06880_);
  or _15195_ (_06884_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not _15196_ (_06885_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _15197_ (_06886_, _06883_, _06885_);
  and _15198_ (_06887_, _06886_, _06884_);
  and _15199_ (_06888_, _06618_, _05802_);
  and _15200_ (_06889_, _05807_, _06472_);
  and _15201_ (_06890_, _06889_, _06888_);
  or _15202_ (_06891_, _06890_, _06887_);
  nand _15203_ (_06892_, _06890_, _06798_);
  and _15204_ (_06893_, _06892_, _06891_);
  and _15205_ (_06894_, _06631_, _05807_);
  and _15206_ (_06895_, _06894_, _06888_);
  or _15207_ (_06896_, _06895_, _06893_);
  not _15208_ (_06897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _15209_ (_06898_, _06895_, _06897_);
  and _15210_ (_06899_, _06898_, _05110_);
  and _15211_ (_05216_, _06899_, _06896_);
  and _15212_ (_06901_, _05999_, _05337_);
  and _15213_ (_06902_, _06183_, _06901_);
  and _15214_ (_06903_, _06174_, _05337_);
  or _15215_ (_06904_, _06903_, _06006_);
  and _15216_ (_06905_, _06904_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or _15217_ (_06906_, _06905_, _06902_);
  and _15218_ (_05289_, _06906_, _05110_);
  and _15219_ (_06907_, _05472_, _05151_);
  and _15220_ (_06908_, _06907_, _06871_);
  not _15221_ (_06909_, _06338_);
  and _15222_ (_06910_, _06315_, _06294_);
  and _15223_ (_06911_, _06910_, _06909_);
  not _15224_ (_06912_, _06362_);
  not _15225_ (_06913_, _06406_);
  and _15226_ (_06914_, _06427_, _06384_);
  and _15227_ (_06915_, _06914_, _06913_);
  and _15228_ (_06916_, _06915_, _06912_);
  and _15229_ (_06917_, _06916_, _06911_);
  not _15230_ (_06918_, _06294_);
  and _15231_ (_06920_, _06315_, _06918_);
  and _15232_ (_06921_, _06920_, _06338_);
  and _15233_ (_06922_, _06915_, _06362_);
  and _15234_ (_06923_, _06922_, _06921_);
  not _15235_ (_06924_, _06427_);
  nor _15236_ (_06925_, _06924_, _06384_);
  and _15237_ (_06926_, _06925_, _06406_);
  and _15238_ (_06927_, _06926_, _06912_);
  not _15239_ (_06928_, _06271_);
  and _15240_ (_06929_, _06920_, _06928_);
  and _15241_ (_06930_, _06929_, _06927_);
  or _15242_ (_06931_, _06930_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _15243_ (_06932_, _06931_, _06923_);
  or _15244_ (_06933_, _06932_, _06917_);
  and _15245_ (_06934_, _06933_, _06908_);
  nor _15246_ (_06935_, _06907_, _06871_);
  or _15247_ (_06936_, _06935_, rst);
  or _15248_ (_05315_, _06936_, _06934_);
  and _15249_ (_06937_, _06807_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and _15250_ (_06938_, _06864_, _06811_);
  and _15251_ (_06939_, _06811_, _06448_);
  or _15252_ (_06940_, _06939_, _06938_);
  and _15253_ (_06941_, _06864_, _06343_);
  or _15254_ (_06942_, _06941_, _06458_);
  or _15255_ (_06943_, _06942_, _06940_);
  or _15256_ (_06944_, _06832_, _06812_);
  or _15257_ (_06945_, _06944_, _06449_);
  or _15258_ (_06946_, _06820_, _06463_);
  and _15259_ (_06947_, _06820_, _06434_);
  or _15260_ (_06948_, _06810_, _06460_);
  or _15261_ (_06949_, _06948_, _06947_);
  and _15262_ (_06950_, _06949_, _06946_);
  or _15263_ (_06951_, _06950_, _06945_);
  or _15264_ (_06952_, _06951_, _06943_);
  and _15265_ (_06953_, _06952_, _06842_);
  or _15266_ (_05331_, _06953_, _06937_);
  not _15267_ (_06954_, _06842_);
  nor _15268_ (_06955_, _06853_, _06849_);
  or _15269_ (_05342_, _06955_, _06954_);
  nor _15270_ (_06956_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _15271_ (_06957_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _05496_);
  nor _15272_ (_06958_, _06957_, _06956_);
  or _15273_ (_06959_, _06958_, _06706_);
  nand _15274_ (_06960_, _06958_, _06706_);
  nand _15275_ (_06962_, _06960_, _06959_);
  nand _15276_ (_06963_, _06962_, _05489_);
  nor _15277_ (_06964_, _06734_, _05812_);
  and _15278_ (_06966_, _06964_, _06726_);
  and _15279_ (_06967_, _06966_, _05517_);
  nor _15280_ (_06968_, _06966_, _05517_);
  nor _15281_ (_06969_, _06968_, _06967_);
  nor _15282_ (_06970_, _06969_, _05882_);
  and _15283_ (_06971_, _06487_, ABINPUT000[16]);
  nor _15284_ (_06972_, _05517_, _05187_);
  nor _15285_ (_06973_, _06972_, _05738_);
  nor _15286_ (_06974_, _06973_, _05321_);
  nor _15287_ (_06975_, _05210_, _05763_);
  nor _15288_ (_06976_, _05517_, _05159_);
  and _15289_ (_06977_, _06485_, ABINPUT000000[16]);
  or _15290_ (_06978_, _06977_, _06976_);
  or _15291_ (_06979_, _06978_, _06975_);
  or _15292_ (_06980_, _06979_, _06974_);
  nor _15293_ (_06981_, _06980_, _06971_);
  not _15294_ (_06982_, _06981_);
  nor _15295_ (_06983_, _06982_, _06970_);
  nand _15296_ (_06984_, _06983_, _06963_);
  and _15297_ (_06985_, _06984_, _06613_);
  and _15298_ (_06986_, _06628_, _05867_);
  nor _15299_ (_06987_, _06986_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _15300_ (_06988_, _06987_);
  and _15301_ (_06989_, _06988_, _06638_);
  not _15302_ (_06990_, _06989_);
  and _15303_ (_06991_, _06986_, _05872_);
  nor _15304_ (_06992_, _06991_, _06990_);
  not _15305_ (_06993_, _05654_);
  and _15306_ (_06994_, _05716_, _06993_);
  nor _15307_ (_06996_, _05716_, _06993_);
  nor _15308_ (_06997_, _06996_, _06994_);
  and _15309_ (_06998_, _06997_, _05650_);
  not _15310_ (_06999_, _06998_);
  nor _15311_ (_07000_, _06993_, _05646_);
  and _15312_ (_07001_, _06993_, _05646_);
  nor _15313_ (_07002_, _07001_, _07000_);
  and _15314_ (_07003_, _07002_, _05489_);
  and _15315_ (_07004_, _05280_, _05766_);
  and _15316_ (_07005_, _06487_, ABINPUT000[8]);
  or _15317_ (_07006_, _07005_, _07004_);
  nor _15318_ (_07007_, _05627_, _05174_);
  nor _15319_ (_07008_, _05510_, _05159_);
  and _15320_ (_07009_, _05187_, _05744_);
  and _15321_ (_07010_, _06485_, ABINPUT000000[8]);
  or _15322_ (_07011_, _07010_, _07009_);
  or _15323_ (_07012_, _07011_, _07008_);
  nor _15324_ (_07013_, _07012_, _07007_);
  nand _15325_ (_07014_, _07013_, _05894_);
  or _15326_ (_07015_, _07014_, _07006_);
  nor _15327_ (_07016_, _06531_, _05732_);
  and _15328_ (_07017_, _07016_, _05510_);
  nor _15329_ (_07018_, _07016_, _05510_);
  nor _15330_ (_07019_, _07018_, _07017_);
  nor _15331_ (_07020_, _07019_, _05737_);
  not _15332_ (_07021_, _07020_);
  nand _15333_ (_07023_, _07021_, _05891_);
  or _15334_ (_07024_, _07023_, _07015_);
  nor _15335_ (_07025_, _07024_, _05898_);
  not _15336_ (_07026_, _07025_);
  nor _15337_ (_07027_, _07026_, _07003_);
  and _15338_ (_07028_, _07027_, _06999_);
  nor _15339_ (_07029_, _07028_, _06622_);
  or _15340_ (_07030_, _07029_, _06992_);
  and _15341_ (_07031_, _07030_, _06637_);
  or _15342_ (_07032_, _07031_, _06985_);
  and _15343_ (_05360_, _07032_, _05110_);
  and _15344_ (_07033_, _06177_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor _15345_ (_07034_, _06798_, _05995_);
  and _15346_ (_07035_, _07034_, _06165_);
  or _15347_ (_07037_, _07035_, _07033_);
  and _15348_ (_05428_, _07037_, _05110_);
  and _15349_ (_07038_, _06813_, _06342_);
  and _15350_ (_07039_, _07038_, _06431_);
  and _15351_ (_07040_, _06460_, _06276_);
  and _15352_ (_07041_, _07040_, _06437_);
  or _15353_ (_07043_, _07041_, _07039_);
  and _15354_ (_07044_, _07038_, _06460_);
  and _15355_ (_07045_, _06452_, _06431_);
  or _15356_ (_07046_, _07045_, _07044_);
  and _15357_ (_07048_, _07038_, _06464_);
  or _15358_ (_07049_, _07048_, _07046_);
  or _15359_ (_07050_, _07049_, _07043_);
  and _15360_ (_07051_, _06810_, _06452_);
  or _15361_ (_07052_, _07051_, _06837_);
  or _15362_ (_07053_, _07052_, _06442_);
  or _15363_ (_07054_, _07053_, _07050_);
  and _15364_ (_07055_, _07054_, _06842_);
  nor _15365_ (_07056_, _06870_, _06440_);
  and _15366_ (_07057_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _15367_ (_07058_, _07057_, _07056_);
  and _15368_ (_07059_, _07058_, _05110_);
  or _15369_ (_05430_, _07059_, _07055_);
  and _15370_ (_07060_, _06807_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _15371_ (_07061_, _07040_, _06459_);
  nor _15372_ (_07062_, _06431_, _06276_);
  and _15373_ (_07063_, _07062_, _06826_);
  and _15374_ (_07064_, _07063_, _06459_);
  or _15375_ (_07065_, _07064_, _07061_);
  not _15376_ (_07066_, _06460_);
  not _15377_ (_07067_, _06298_);
  and _15378_ (_07068_, _06851_, _07067_);
  and _15379_ (_07069_, _07068_, _06277_);
  and _15380_ (_07070_, _06319_, _07067_);
  and _15381_ (_07071_, _07070_, _06436_);
  and _15382_ (_07072_, _07071_, _06277_);
  nor _15383_ (_07073_, _07072_, _07069_);
  nor _15384_ (_07074_, _07073_, _07066_);
  or _15385_ (_07075_, _07074_, _07065_);
  and _15386_ (_07076_, _07069_, _06447_);
  and _15387_ (_07077_, _06451_, _06343_);
  and _15388_ (_07078_, _07069_, _06464_);
  and _15389_ (_07079_, _06456_, _07067_);
  and _15390_ (_07080_, _07079_, _06277_);
  and _15391_ (_07081_, _07080_, _06810_);
  or _15392_ (_07082_, _07081_, _07078_);
  or _15393_ (_07083_, _07082_, _07077_);
  or _15394_ (_07084_, _07083_, _07076_);
  or _15395_ (_07085_, _07084_, _07075_);
  and _15396_ (_07086_, _07080_, _06447_);
  and _15397_ (_07087_, _07068_, _06276_);
  and _15398_ (_07088_, _07087_, _06864_);
  and _15399_ (_07089_, _07080_, _06434_);
  or _15400_ (_07090_, _07089_, _07088_);
  or _15401_ (_07091_, _07090_, _07086_);
  not _15402_ (_07092_, _06834_);
  and _15403_ (_07093_, _06813_, _06448_);
  or _15404_ (_07094_, _07093_, _07092_);
  and _15405_ (_07095_, _07068_, _06455_);
  or _15406_ (_07096_, _07095_, _06457_);
  or _15407_ (_07097_, _06823_, _06465_);
  or _15408_ (_07098_, _07097_, _07096_);
  or _15409_ (_07099_, _07098_, _07094_);
  or _15410_ (_07100_, _07099_, _06822_);
  or _15411_ (_07101_, _07100_, _07091_);
  or _15412_ (_07103_, _07101_, _07085_);
  and _15413_ (_07104_, _07103_, _06842_);
  or _15414_ (_05477_, _07104_, _07060_);
  and _15415_ (_07105_, _06864_, _06814_);
  and _15416_ (_07106_, _07105_, _06276_);
  and _15417_ (_07107_, _06810_, _06276_);
  and _15418_ (_07108_, _07107_, _06851_);
  or _15419_ (_07109_, _06811_, _06452_);
  nand _15420_ (_07110_, _07109_, _06864_);
  not _15421_ (_07111_, _07110_);
  or _15422_ (_07113_, _07111_, _07108_);
  or _15423_ (_07114_, _07113_, _07106_);
  and _15424_ (_07115_, _06831_, _06810_);
  and _15425_ (_07116_, _06459_, _06451_);
  or _15426_ (_07117_, _07116_, _06845_);
  or _15427_ (_07118_, _07117_, _07115_);
  or _15428_ (_07119_, _07118_, _07086_);
  and _15429_ (_07120_, _06864_, _06463_);
  and _15430_ (_07121_, _06941_, _06276_);
  or _15431_ (_07122_, _07121_, _07120_);
  or _15432_ (_07123_, _07122_, _07076_);
  or _15433_ (_07124_, _07123_, _07119_);
  or _15434_ (_07125_, _07124_, _07114_);
  and _15435_ (_07126_, _06851_, _06830_);
  and _15436_ (_07127_, _06455_, _06343_);
  or _15437_ (_07128_, _07127_, _07126_);
  nor _15438_ (_07129_, _07128_, _06462_);
  nand _15439_ (_07130_, _07129_, _06834_);
  and _15440_ (_07131_, _06851_, _07040_);
  and _15441_ (_07132_, _07063_, _06343_);
  or _15442_ (_07133_, _07132_, _06823_);
  or _15443_ (_07134_, _07133_, _07131_);
  and _15444_ (_07135_, _06455_, _06437_);
  or _15445_ (_07136_, _07135_, _06867_);
  and _15446_ (_07137_, _06460_, _06438_);
  and _15447_ (_07138_, _07079_, _06276_);
  and _15448_ (_07139_, _07138_, _06447_);
  or _15449_ (_07140_, _07139_, _07137_);
  or _15450_ (_07141_, _07140_, _07136_);
  or _15451_ (_07142_, _07141_, _07134_);
  or _15452_ (_07143_, _07142_, _07130_);
  or _15453_ (_07144_, _07143_, _07125_);
  and _15454_ (_07145_, _07144_, _05474_);
  and _15455_ (_07146_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and _15456_ (_07147_, _06820_, _06451_);
  and _15457_ (_07148_, _07147_, _06873_);
  or _15458_ (_07149_, _06874_, _06443_);
  or _15459_ (_07150_, _07149_, _07148_);
  or _15460_ (_07151_, _07150_, _07146_);
  or _15461_ (_07152_, _07151_, _07145_);
  and _15462_ (_05513_, _07152_, _05110_);
  not _15463_ (_07153_, _05473_);
  or _15464_ (_07154_, _06362_, _07153_);
  or _15465_ (_07155_, _05473_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _15466_ (_07156_, _07155_, _05110_);
  and _15467_ (_05525_, _07156_, _07154_);
  nor _15468_ (_05565_, _06294_, rst);
  nor _15469_ (_07157_, _05474_, _05492_);
  and _15470_ (_07158_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _15471_ (_07159_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _15472_ (_07160_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _15473_ (_07161_, _07160_, _07159_);
  and _15474_ (_07162_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _15475_ (_07163_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _15476_ (_07164_, _07163_, _07162_);
  and _15477_ (_07165_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  not _15478_ (_07167_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _15479_ (_07168_, _06251_, _07167_);
  nor _15480_ (_07169_, _07168_, _07165_);
  and _15481_ (_07170_, _07169_, _07164_);
  and _15482_ (_07171_, _07170_, _07161_);
  nor _15483_ (_07172_, _07171_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _15484_ (_07173_, _07172_, _07158_);
  nor _15485_ (_07174_, _07173_, _06200_);
  nor _15486_ (_07176_, _07174_, _07157_);
  nor _15487_ (_05569_, _07176_, rst);
  not _15488_ (_07177_, _06471_);
  or _15489_ (_07178_, _06699_, _06693_);
  nand _15490_ (_07179_, _06699_, _06693_);
  and _15491_ (_07180_, _07179_, _05489_);
  nand _15492_ (_07181_, _07180_, _07178_);
  and _15493_ (_07182_, _06588_, _05526_);
  and _15494_ (_07183_, _06593_, _05703_);
  nor _15495_ (_07184_, _07183_, _07182_);
  and _15496_ (_07185_, _07184_, _05306_);
  nor _15497_ (_07186_, _07184_, _05306_);
  nor _15498_ (_07187_, _07186_, _07185_);
  and _15499_ (_07188_, _07187_, _05291_);
  and _15500_ (_07190_, _06487_, ABINPUT000[13]);
  nor _15501_ (_07191_, _05306_, _05187_);
  nor _15502_ (_07192_, _05188_, _05150_);
  or _15503_ (_07193_, _07192_, _07191_);
  and _15504_ (_07194_, _07193_, _05320_);
  and _15505_ (_07195_, _05280_, _05762_);
  nor _15506_ (_07196_, _05306_, _05159_);
  and _15507_ (_07197_, _06485_, ABINPUT000000[13]);
  or _15508_ (_07198_, _07197_, _07196_);
  or _15509_ (_07199_, _07198_, _07195_);
  or _15510_ (_07200_, _07199_, _07194_);
  nor _15511_ (_07201_, _07200_, _07190_);
  not _15512_ (_07202_, _07201_);
  nor _15513_ (_07203_, _07202_, _07188_);
  nand _15514_ (_07204_, _07203_, _07181_);
  or _15515_ (_07205_, _07204_, _07177_);
  and _15516_ (_07206_, _06146_, _05804_);
  and _15517_ (_07207_, _07206_, _06631_);
  not _15518_ (_07208_, _07207_);
  nor _15519_ (_07209_, _05711_, _05309_);
  and _15520_ (_07210_, _05711_, _05309_);
  nor _15521_ (_07211_, _07210_, _07209_);
  and _15522_ (_07212_, _07211_, _05650_);
  not _15523_ (_07213_, _07212_);
  nor _15524_ (_07214_, _05575_, _05309_);
  nor _15525_ (_07215_, _07214_, _05490_);
  and _15526_ (_07216_, _07215_, _05576_);
  nor _15527_ (_07217_, _06649_, _05158_);
  nor _15528_ (_07218_, _07217_, _05150_);
  not _15529_ (_07219_, _07218_);
  and _15530_ (_07220_, _05729_, _05150_);
  or _15531_ (_07221_, _05597_, _05169_);
  nor _15532_ (_07222_, _05210_, _05174_);
  and _15533_ (_07223_, _06485_, ABINPUT000000[5]);
  and _15534_ (_07224_, _06487_, ABINPUT000[5]);
  nor _15535_ (_07225_, _07224_, _07223_);
  not _15536_ (_07226_, _07225_);
  nor _15537_ (_07227_, _07226_, _07222_);
  and _15538_ (_07228_, _07227_, _07221_);
  not _15539_ (_07229_, _07228_);
  nor _15540_ (_07230_, _07229_, _07220_);
  and _15541_ (_07231_, _07230_, _07219_);
  and _15542_ (_07232_, _07231_, _05333_);
  not _15543_ (_07233_, _07232_);
  nor _15544_ (_07234_, _07233_, _07216_);
  and _15545_ (_07235_, _07234_, _07213_);
  nor _15546_ (_07236_, _07235_, _07208_);
  and _15547_ (_07237_, _07208_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _15548_ (_07238_, _07237_, _06471_);
  or _15549_ (_07239_, _07238_, _07236_);
  and _15550_ (_07240_, _07239_, _05110_);
  and _15551_ (_05657_, _07240_, _07205_);
  or _15552_ (_07241_, _06610_, _07177_);
  nand _15553_ (_07242_, _07207_, _06668_);
  or _15554_ (_07243_, _07207_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _15555_ (_07244_, _07243_, _07242_);
  or _15556_ (_07245_, _07244_, _06471_);
  and _15557_ (_07246_, _07245_, _05110_);
  and _15558_ (_05660_, _07246_, _07241_);
  or _15559_ (_07247_, _06745_, _07177_);
  nor _15560_ (_07248_, _07208_, _06780_);
  and _15561_ (_07250_, _07208_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _15562_ (_07251_, _07250_, _06471_);
  or _15563_ (_07252_, _07251_, _07248_);
  and _15564_ (_07253_, _07252_, _05110_);
  and _15565_ (_05665_, _07253_, _07247_);
  not _15566_ (_07254_, _06696_);
  nand _15567_ (_07255_, _07179_, _07254_);
  nor _15568_ (_07256_, _06701_, _05490_);
  nand _15569_ (_07257_, _07256_, _07255_);
  and _15570_ (_07258_, _06722_, _05603_);
  not _15571_ (_07259_, _07258_);
  nor _15572_ (_07260_, _06722_, _05603_);
  nor _15573_ (_07261_, _07260_, _05882_);
  and _15574_ (_07262_, _07261_, _07259_);
  and _15575_ (_07263_, _05281_, _05762_);
  and _15576_ (_07264_, _06487_, ABINPUT000[14]);
  nor _15577_ (_07265_, _07264_, _07263_);
  and _15578_ (_07266_, _05597_, _05187_);
  not _15579_ (_07267_, _07266_);
  nor _15580_ (_07268_, _06723_, _05321_);
  and _15581_ (_07269_, _07268_, _07267_);
  nor _15582_ (_07270_, _05603_, _05159_);
  and _15583_ (_07271_, _06485_, ABINPUT000000[14]);
  or _15584_ (_07272_, _07271_, _07270_);
  nor _15585_ (_07273_, _07272_, _07269_);
  and _15586_ (_07274_, _07273_, _07265_);
  not _15587_ (_07275_, _07274_);
  nor _15588_ (_07276_, _07275_, _07262_);
  nand _15589_ (_07277_, _07276_, _07257_);
  or _15590_ (_07278_, _07277_, _07177_);
  nor _15591_ (_07279_, _07208_, _06548_);
  and _15592_ (_07280_, _07208_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _15593_ (_07281_, _07280_, _06471_);
  or _15594_ (_07282_, _07281_, _07279_);
  and _15595_ (_07283_, _07282_, _05110_);
  and _15596_ (_05670_, _07283_, _07278_);
  or _15597_ (_07284_, _06575_, _06572_);
  nor _15598_ (_07285_, _06576_, _05490_);
  nand _15599_ (_07286_, _07285_, _07284_);
  nor _15600_ (_07287_, _06586_, _05188_);
  nor _15601_ (_07288_, _06591_, _05187_);
  nor _15602_ (_07289_, _07288_, _07287_);
  and _15603_ (_07290_, _07289_, _05534_);
  nor _15604_ (_07291_, _07289_, _05534_);
  nor _15605_ (_07292_, _07291_, _07290_);
  nor _15606_ (_07293_, _07292_, _05882_);
  nor _15607_ (_07294_, _05627_, _05763_);
  nor _15608_ (_07295_, _05534_, _05159_);
  and _15609_ (_07296_, _06485_, ABINPUT000000[11]);
  or _15610_ (_07297_, _07296_, _07295_);
  nor _15611_ (_07298_, _07297_, _07294_);
  nor _15612_ (_07299_, _05321_, _05233_);
  and _15613_ (_07300_, _06487_, ABINPUT000[11]);
  nor _15614_ (_07301_, _07300_, _07299_);
  and _15615_ (_07302_, _07301_, _07298_);
  not _15616_ (_07303_, _07302_);
  nor _15617_ (_07304_, _07303_, _07293_);
  nand _15618_ (_07305_, _07304_, _07286_);
  or _15619_ (_07306_, _07305_, _07177_);
  or _15620_ (_07307_, _07207_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor _15621_ (_07308_, _05699_, _05692_);
  nor _15622_ (_07309_, _07308_, _05700_);
  nor _15623_ (_07310_, _07309_, _05651_);
  and _15624_ (_07311_, _05726_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _15625_ (_07312_, _06500_, _05233_);
  nor _15626_ (_07313_, _07312_, _07311_);
  nor _15627_ (_07314_, _07313_, _05737_);
  not _15628_ (_07315_, _06226_);
  nor _15629_ (_07316_, _05233_, _05159_);
  and _15630_ (_07317_, _06487_, ABINPUT000[3]);
  nor _15631_ (_07318_, _07317_, _07316_);
  or _15632_ (_07319_, _05210_, _05169_);
  and _15633_ (_07320_, _05281_, _05172_);
  and _15634_ (_07321_, _06485_, ABINPUT000000[3]);
  nor _15635_ (_07322_, _07321_, _07320_);
  and _15636_ (_07323_, _07322_, _07319_);
  and _15637_ (_07324_, _07323_, _07318_);
  and _15638_ (_07325_, _07324_, _07315_);
  not _15639_ (_07326_, _07325_);
  nor _15640_ (_07327_, _07326_, _07314_);
  not _15641_ (_07328_, _07327_);
  nor _15642_ (_07329_, _07328_, _07310_);
  nor _15643_ (_07330_, _05568_, _05566_);
  not _15644_ (_07331_, _07330_);
  nor _15645_ (_07332_, _05570_, _05490_);
  and _15646_ (_07333_, _07332_, _07331_);
  and _15647_ (_07334_, _06222_, _06219_);
  not _15648_ (_07335_, _07334_);
  nor _15649_ (_07336_, _07335_, _07333_);
  and _15650_ (_07337_, _07336_, _07329_);
  nand _15651_ (_07338_, _07337_, _07207_);
  and _15652_ (_07339_, _07338_, _07307_);
  or _15653_ (_07340_, _07339_, _06471_);
  and _15654_ (_07341_, _07340_, _05110_);
  and _15655_ (_05680_, _07341_, _07306_);
  or _15656_ (_07342_, _06571_, _06568_);
  nor _15657_ (_07343_, _06572_, _05490_);
  nand _15658_ (_07344_, _07343_, _07342_);
  nor _15659_ (_07345_, _06711_, _05187_);
  nor _15660_ (_07346_, _06585_, _05188_);
  or _15661_ (_07347_, _07346_, _07345_);
  nor _15662_ (_07348_, _07347_, _05543_);
  and _15663_ (_07349_, _07347_, _05543_);
  nor _15664_ (_07350_, _07349_, _07348_);
  nor _15665_ (_07351_, _07350_, _05882_);
  nor _15666_ (_07352_, _05597_, _05763_);
  and _15667_ (_07353_, _05543_, _05158_);
  and _15668_ (_07354_, _06485_, ABINPUT000000[10]);
  or _15669_ (_07355_, _07354_, _07353_);
  nor _15670_ (_07356_, _07355_, _07352_);
  and _15671_ (_07358_, _05320_, _05281_);
  and _15672_ (_07359_, _06487_, ABINPUT000[10]);
  nor _15673_ (_07360_, _07359_, _07358_);
  and _15674_ (_07361_, _07360_, _07356_);
  not _15675_ (_07362_, _07361_);
  nor _15676_ (_07363_, _07362_, _07351_);
  nand _15677_ (_07364_, _07363_, _07344_);
  or _15678_ (_07365_, _07364_, _07177_);
  or _15679_ (_07366_, _07207_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nand _15680_ (_07367_, _07207_, _06512_);
  and _15681_ (_07368_, _07367_, _07366_);
  or _15682_ (_07369_, _07368_, _06471_);
  and _15683_ (_07370_, _07369_, _05110_);
  and _15684_ (_05688_, _07370_, _07365_);
  or _15685_ (_07371_, _06567_, _06564_);
  nor _15686_ (_07372_, _06568_, _05490_);
  nand _15687_ (_07373_, _07372_, _07371_);
  nor _15688_ (_07374_, _06584_, _05876_);
  nor _15689_ (_07375_, _07374_, _05886_);
  nor _15690_ (_07376_, _07375_, _05550_);
  and _15691_ (_07377_, _07375_, _05550_);
  nor _15692_ (_07378_, _07377_, _07376_);
  and _15693_ (_07379_, _07378_, _05291_);
  nor _15694_ (_07380_, _05763_, _05150_);
  nor _15695_ (_07381_, _05549_, _05159_);
  and _15696_ (_07382_, _06485_, ABINPUT000000[9]);
  or _15697_ (_07383_, _07382_, _07381_);
  nor _15698_ (_07384_, _07383_, _07380_);
  and _15699_ (_07385_, _05320_, _05280_);
  and _15700_ (_07386_, _06487_, ABINPUT000[9]);
  nor _15701_ (_07387_, _07386_, _07385_);
  and _15702_ (_07388_, _07387_, _07384_);
  not _15703_ (_07389_, _07388_);
  nor _15704_ (_07390_, _07389_, _07379_);
  nand _15705_ (_07391_, _07390_, _07373_);
  or _15706_ (_07392_, _07391_, _07177_);
  or _15707_ (_07393_, _07207_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nor _15708_ (_07394_, _05563_, _05187_);
  nor _15709_ (_07395_, _07394_, _05564_);
  not _15710_ (_07396_, _07395_);
  nor _15711_ (_07397_, _05489_, _05650_);
  nor _15712_ (_07398_, _07397_, _07396_);
  not _15713_ (_07399_, _07398_);
  and _15714_ (_07400_, _06709_, _05749_);
  not _15715_ (_07401_, _07400_);
  and _15716_ (_07402_, _06794_, _07401_);
  or _15717_ (_07403_, _05274_, _05169_);
  nor _15718_ (_07404_, _05725_, _05158_);
  nor _15719_ (_07405_, _07404_, _05253_);
  not _15720_ (_07406_, _07405_);
  and _15721_ (_07407_, _07406_, _07403_);
  and _15722_ (_07408_, _05187_, _05762_);
  and _15723_ (_07409_, _06485_, ABINPUT000000[1]);
  and _15724_ (_07410_, _06487_, ABINPUT000[1]);
  nor _15725_ (_07411_, _07410_, _07409_);
  not _15726_ (_07412_, _07411_);
  nor _15727_ (_07413_, _07412_, _07408_);
  and _15728_ (_07414_, _07413_, _07407_);
  and _15729_ (_07415_, _07414_, _06791_);
  and _15730_ (_07416_, _07415_, _07402_);
  and _15731_ (_07417_, _07416_, _06788_);
  and _15732_ (_07418_, _07417_, _07399_);
  nand _15733_ (_07419_, _07418_, _07207_);
  and _15734_ (_07420_, _07419_, _07393_);
  or _15735_ (_07421_, _07420_, _06471_);
  and _15736_ (_07422_, _07421_, _05110_);
  and _15737_ (_05691_, _07422_, _07392_);
  and _15738_ (_05695_, _06362_, _05110_);
  and _15739_ (_05698_, _06384_, _05110_);
  and _15740_ (_05701_, _06406_, _05110_);
  nor _15741_ (_05704_, _06427_, rst);
  and _15742_ (_05706_, _06271_, _05110_);
  nor _15743_ (_05709_, _06338_, rst);
  nor _15744_ (_05712_, _06315_, rst);
  nor _15745_ (_07423_, _05474_, _05258_);
  and _15746_ (_07424_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  not _15747_ (_07425_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _15748_ (_07426_, _06251_, _07425_);
  nor _15749_ (_07427_, _07426_, _07424_);
  and _15750_ (_07428_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _15751_ (_07429_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _15752_ (_07430_, _07429_, _07428_);
  and _15753_ (_07431_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _15754_ (_07432_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _15755_ (_07433_, _07432_, _07431_);
  and _15756_ (_07434_, _07433_, _07430_);
  and _15757_ (_07435_, _07434_, _07427_);
  and _15758_ (_07436_, _05474_, _06254_);
  not _15759_ (_07437_, _07436_);
  nor _15760_ (_07438_, _07437_, _07435_);
  nor _15761_ (_07439_, _07438_, _07423_);
  nor _15762_ (_05721_, _07439_, rst);
  nor _15763_ (_07440_, _05474_, _05212_);
  and _15764_ (_07441_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  not _15765_ (_07442_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _15766_ (_07443_, _06251_, _07442_);
  nor _15767_ (_07444_, _07443_, _07441_);
  and _15768_ (_07445_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _15769_ (_07446_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _15770_ (_07447_, _07446_, _07445_);
  and _15771_ (_07448_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _15772_ (_07449_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _15773_ (_07450_, _07449_, _07448_);
  and _15774_ (_07451_, _07450_, _07447_);
  and _15775_ (_07452_, _07451_, _07444_);
  nor _15776_ (_07453_, _07452_, _07437_);
  nor _15777_ (_07454_, _07453_, _07440_);
  nor _15778_ (_05724_, _07454_, rst);
  nor _15779_ (_07455_, _05474_, _05189_);
  and _15780_ (_07456_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  not _15781_ (_07457_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _15782_ (_07458_, _06251_, _07457_);
  nor _15783_ (_07459_, _07458_, _07456_);
  and _15784_ (_07460_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _15785_ (_07461_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _15786_ (_07462_, _07461_, _07460_);
  and _15787_ (_07463_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _15788_ (_07464_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _15789_ (_07465_, _07464_, _07463_);
  and _15790_ (_07466_, _07465_, _07462_);
  and _15791_ (_07467_, _07466_, _07459_);
  nor _15792_ (_07469_, _07467_, _07437_);
  nor _15793_ (_07470_, _07469_, _07455_);
  nor _15794_ (_05727_, _07470_, rst);
  nor _15795_ (_07471_, _05474_, _05111_);
  and _15796_ (_07473_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  not _15797_ (_07474_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _15798_ (_07475_, _06251_, _07474_);
  nor _15799_ (_07477_, _07475_, _07473_);
  and _15800_ (_07478_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _15801_ (_07479_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _15802_ (_07480_, _07479_, _07478_);
  and _15803_ (_07482_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _15804_ (_07483_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _15805_ (_07485_, _07483_, _07482_);
  and _15806_ (_07486_, _07485_, _07480_);
  and _15807_ (_07487_, _07486_, _07477_);
  nor _15808_ (_07489_, _07487_, _07437_);
  nor _15809_ (_07490_, _07489_, _07471_);
  nor _15810_ (_05730_, _07490_, rst);
  nor _15811_ (_07492_, _05474_, _05425_);
  and _15812_ (_07493_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  not _15813_ (_07494_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _15814_ (_07496_, _06251_, _07494_);
  nor _15815_ (_07497_, _07496_, _07493_);
  and _15816_ (_07498_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _15817_ (_07499_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _15818_ (_07500_, _07499_, _07498_);
  and _15819_ (_07501_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _15820_ (_07502_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _15821_ (_07503_, _07502_, _07501_);
  and _15822_ (_07504_, _07503_, _07500_);
  and _15823_ (_07505_, _07504_, _07497_);
  nor _15824_ (_07506_, _07505_, _07437_);
  nor _15825_ (_07507_, _07506_, _07492_);
  nor _15826_ (_05733_, _07507_, rst);
  nor _15827_ (_07508_, _05474_, _05260_);
  and _15828_ (_07509_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _15829_ (_07510_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _15830_ (_07511_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _15831_ (_07512_, _07511_, _07510_);
  and _15832_ (_07513_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  not _15833_ (_07514_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _15834_ (_07515_, _06251_, _07514_);
  nor _15835_ (_07516_, _07515_, _07513_);
  and _15836_ (_07517_, _07516_, _07512_);
  and _15837_ (_07518_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _15838_ (_07519_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _15839_ (_07520_, _07519_, _07518_);
  and _15840_ (_07521_, _07520_, _07517_);
  nor _15841_ (_07522_, _07521_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _15842_ (_07523_, _07522_, _07509_);
  nor _15843_ (_07524_, _07523_, _06200_);
  nor _15844_ (_07525_, _07524_, _07508_);
  nor _15845_ (_05745_, _07525_, rst);
  nor _15846_ (_07526_, _05474_, _05214_);
  and _15847_ (_07527_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _15848_ (_07528_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _15849_ (_07529_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _15850_ (_07530_, _07529_, _07528_);
  and _15851_ (_07531_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  not _15852_ (_07532_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _15853_ (_07533_, _06251_, _07532_);
  nor _15854_ (_07534_, _07533_, _07531_);
  and _15855_ (_07535_, _07534_, _07530_);
  and _15856_ (_07536_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _15857_ (_07537_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _15858_ (_07538_, _07537_, _07536_);
  and _15859_ (_07539_, _07538_, _07535_);
  nor _15860_ (_07540_, _07539_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _15861_ (_07541_, _07540_, _07527_);
  nor _15862_ (_07542_, _07541_, _06200_);
  nor _15863_ (_07543_, _07542_, _07526_);
  nor _15864_ (_05748_, _07543_, rst);
  nor _15865_ (_07544_, _05474_, _05191_);
  and _15866_ (_07545_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _15867_ (_07546_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _15868_ (_07547_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _15869_ (_07548_, _07547_, _07546_);
  and _15870_ (_07549_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _15871_ (_07550_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _15872_ (_07551_, _07550_, _07549_);
  and _15873_ (_07552_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  not _15874_ (_07553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _15875_ (_07554_, _06251_, _07553_);
  nor _15876_ (_07555_, _07554_, _07552_);
  and _15877_ (_07556_, _07555_, _07551_);
  and _15878_ (_07557_, _07556_, _07548_);
  nor _15879_ (_07558_, _07557_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _15880_ (_07559_, _07558_, _07545_);
  nor _15881_ (_07560_, _07559_, _06200_);
  nor _15882_ (_07561_, _07560_, _07544_);
  nor _15883_ (_05750_, _07561_, rst);
  nor _15884_ (_07562_, _05474_, _05610_);
  and _15885_ (_07563_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _15886_ (_07564_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _15887_ (_07565_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _15888_ (_07566_, _07565_, _07564_);
  and _15889_ (_07567_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _15890_ (_07568_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _15891_ (_07569_, _07568_, _07567_);
  and _15892_ (_07570_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  not _15893_ (_07571_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _15894_ (_07572_, _06251_, _07571_);
  nor _15895_ (_07574_, _07572_, _07570_);
  and _15896_ (_07575_, _07574_, _07569_);
  and _15897_ (_07576_, _07575_, _07566_);
  nor _15898_ (_07578_, _07576_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _15899_ (_07579_, _07578_, _07563_);
  nor _15900_ (_07580_, _07579_, _06200_);
  nor _15901_ (_07582_, _07580_, _07562_);
  nor _15902_ (_05757_, _07582_, rst);
  nand _15903_ (_07583_, _07235_, _06477_);
  or _15904_ (_07585_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _15905_ (_07586_, _07585_, _05110_);
  and _15906_ (_05772_, _07586_, _07583_);
  nor _15907_ (_07588_, _07418_, _06476_);
  and _15908_ (_07589_, _06476_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or _15909_ (_07591_, _07589_, _07588_);
  and _15910_ (_05775_, _07591_, _05110_);
  nand _15911_ (_07592_, _06668_, _06477_);
  or _15912_ (_07594_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _15913_ (_07595_, _07594_, _05110_);
  and _15914_ (_05780_, _07595_, _07592_);
  nand _15915_ (_07596_, _06780_, _06477_);
  or _15916_ (_07598_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _15917_ (_07599_, _07598_, _05110_);
  and _15918_ (_05783_, _07599_, _07596_);
  nor _15919_ (_07600_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  not _15920_ (_07601_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _15921_ (_07602_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _07601_);
  nor _15922_ (_07603_, _07602_, _07600_);
  not _15923_ (_07604_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not _15924_ (_07605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _15925_ (_07606_, _06205_, _07605_);
  and _15926_ (_07607_, _07606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _15927_ (_07608_, _07606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _15928_ (_07609_, _07608_, _07607_);
  nor _15929_ (_07610_, _07609_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _15930_ (_07611_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _07601_);
  nor _15931_ (_07612_, _07611_, _07610_);
  nor _15932_ (_07613_, _07612_, _07604_);
  and _15933_ (_07614_, _07612_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _15934_ (_07615_, _07614_, _07613_);
  nor _15935_ (_07616_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _15936_ (_07617_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _07601_);
  nor _15937_ (_07618_, _07617_, _07616_);
  and _15938_ (_07619_, _06205_, _07605_);
  nor _15939_ (_07620_, _07619_, _07606_);
  nor _15940_ (_07621_, _07620_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _15941_ (_07622_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _07601_);
  nor _15942_ (_07623_, _07622_, _07621_);
  nor _15943_ (_07624_, _07623_, _07618_);
  not _15944_ (_07625_, _07624_);
  nor _15945_ (_07626_, _07625_, _07615_);
  not _15946_ (_07627_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _15947_ (_07628_, _07612_, _07627_);
  nor _15948_ (_07629_, _07612_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _15949_ (_07630_, _07629_, _07628_);
  not _15950_ (_07631_, _07630_);
  not _15951_ (_07632_, _07618_);
  and _15952_ (_07633_, _07623_, _07632_);
  and _15953_ (_07634_, _07633_, _07631_);
  nor _15954_ (_07635_, _07634_, _07626_);
  nor _15955_ (_07636_, _07623_, _07632_);
  not _15956_ (_07637_, _07636_);
  not _15957_ (_07638_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _15958_ (_07640_, _07612_, _07638_);
  and _15959_ (_07641_, _07612_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _15960_ (_07642_, _07641_, _07640_);
  nor _15961_ (_07643_, _07642_, _07637_);
  and _15962_ (_07644_, _07623_, _07618_);
  not _15963_ (_07645_, _07644_);
  nor _15964_ (_07646_, _07612_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not _15965_ (_07647_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _15966_ (_07649_, _07612_, _07647_);
  or _15967_ (_07650_, _07649_, _07646_);
  nor _15968_ (_07651_, _07650_, _07645_);
  nor _15969_ (_07652_, _07651_, _07643_);
  and _15970_ (_07654_, _07652_, _07635_);
  and _15971_ (_07656_, _07654_, _07603_);
  and _15972_ (_07657_, _07612_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _15973_ (_07658_, _07657_, _07636_);
  not _15974_ (_07659_, _07612_);
  and _15975_ (_07660_, _07659_, _07636_);
  and _15976_ (_07661_, _07660_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _15977_ (_07662_, _07661_, _07603_);
  or _15978_ (_07663_, _07662_, _07658_);
  and _15979_ (_07664_, _07612_, \oc8051_symbolic_cxrom1.regvalid [8]);
  not _15980_ (_07666_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _15981_ (_07667_, _07612_, _07666_);
  nor _15982_ (_07668_, _07667_, _07664_);
  nor _15983_ (_07669_, _07668_, _07625_);
  and _15984_ (_07670_, _07659_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _15985_ (_07671_, _07612_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _15986_ (_07672_, _07671_, _07670_);
  nor _15987_ (_07673_, _07672_, _07645_);
  not _15988_ (_07674_, _07633_);
  not _15989_ (_07675_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _15990_ (_07676_, _07612_, _07675_);
  nor _15991_ (_07677_, _07612_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _15992_ (_07678_, _07677_, _07676_);
  nor _15993_ (_07679_, _07678_, _07674_);
  or _15994_ (_07680_, _07679_, _07673_);
  or _15995_ (_07681_, _07680_, _07669_);
  nor _15996_ (_07682_, _07681_, _07663_);
  nor _15997_ (_07683_, _07682_, _07656_);
  not _15998_ (_07684_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _15999_ (_07685_, _07603_, _07684_);
  or _16000_ (_07687_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _16001_ (_07688_, _07687_, _07685_);
  and _16002_ (_07690_, _07688_, _07644_);
  not _16003_ (_07691_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _16004_ (_07693_, _07603_, _07691_);
  or _16005_ (_07694_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _16006_ (_07695_, _07694_, _07693_);
  and _16007_ (_07696_, _07695_, _07636_);
  or _16008_ (_07698_, _07696_, _07690_);
  not _16009_ (_07699_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _16010_ (_07701_, _07603_, _07699_);
  or _16011_ (_07702_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _16012_ (_07704_, _07702_, _07701_);
  and _16013_ (_07705_, _07704_, _07633_);
  not _16014_ (_07706_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _16015_ (_07707_, _07603_, _07706_);
  or _16016_ (_07709_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _16017_ (_07710_, _07709_, _07707_);
  and _16018_ (_07711_, _07710_, _07624_);
  or _16019_ (_07712_, _07711_, _07705_);
  or _16020_ (_07714_, _07712_, _07698_);
  and _16021_ (_07715_, _07714_, _07612_);
  not _16022_ (_07716_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _16023_ (_07717_, _07603_, _07716_);
  or _16024_ (_07718_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _16025_ (_07719_, _07718_, _07717_);
  and _16026_ (_07720_, _07719_, _07636_);
  not _16027_ (_07721_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _16028_ (_07722_, _07603_, _07721_);
  or _16029_ (_07723_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _16030_ (_07724_, _07723_, _07722_);
  and _16031_ (_07725_, _07724_, _07644_);
  or _16032_ (_07726_, _07725_, _07720_);
  not _16033_ (_07727_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _16034_ (_07728_, _07603_, _07727_);
  or _16035_ (_07729_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _16036_ (_07730_, _07729_, _07728_);
  and _16037_ (_07731_, _07730_, _07633_);
  not _16038_ (_07732_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand _16039_ (_07733_, _07603_, _07732_);
  or _16040_ (_07734_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _16041_ (_07735_, _07734_, _07733_);
  and _16042_ (_07736_, _07735_, _07624_);
  or _16043_ (_07737_, _07736_, _07731_);
  or _16044_ (_07738_, _07737_, _07726_);
  and _16045_ (_07739_, _07738_, _07659_);
  or _16046_ (_07740_, _07739_, _07715_);
  and _16047_ (_07741_, _07740_, _07683_);
  not _16048_ (_07742_, _07683_);
  and _16049_ (_07743_, _07742_, word_in[7]);
  or _16050_ (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _07743_, _07741_);
  and _16051_ (_07744_, _07632_, _07603_);
  not _16052_ (_07745_, _07744_);
  and _16053_ (_07746_, _07618_, _07603_);
  nor _16054_ (_07747_, _07746_, _07623_);
  and _16055_ (_07748_, _07746_, _07623_);
  nor _16056_ (_07749_, _07748_, _07747_);
  not _16057_ (_07750_, _07749_);
  nor _16058_ (_07751_, _07750_, _07672_);
  nor _16059_ (_07752_, _07748_, _07659_);
  not _16060_ (_07753_, _07623_);
  nor _16061_ (_07754_, _07612_, _07753_);
  and _16062_ (_07755_, _07746_, _07754_);
  nor _16063_ (_07756_, _07755_, _07752_);
  nor _16064_ (_07757_, _07756_, _07749_);
  and _16065_ (_07759_, _07757_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16066_ (_07760_, _07756_, _07750_);
  and _16067_ (_07761_, _07760_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _16068_ (_07762_, _07761_, _07759_);
  nor _16069_ (_07763_, _07762_, _07751_);
  nor _16070_ (_07764_, _07763_, _07745_);
  not _16071_ (_07765_, _07764_);
  not _16072_ (_07766_, _07746_);
  nor _16073_ (_07767_, _07750_, _07678_);
  and _16074_ (_07768_, _07760_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _16075_ (_07769_, _07768_, _07767_);
  or _16076_ (_07770_, _07769_, _07766_);
  nand _16077_ (_07771_, _07755_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16078_ (_07772_, _07771_, _07770_);
  and _16079_ (_07773_, _07772_, _07765_);
  not _16080_ (_07774_, _07603_);
  and _16081_ (_07775_, _07618_, _07774_);
  not _16082_ (_07776_, _07775_);
  nor _16083_ (_07777_, _07750_, _07650_);
  and _16084_ (_07778_, _07757_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _16085_ (_07779_, _07760_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or _16086_ (_07780_, _07779_, _07778_);
  nor _16087_ (_07781_, _07780_, _07777_);
  nor _16088_ (_07782_, _07781_, _07776_);
  nor _16089_ (_07783_, _07618_, _07603_);
  not _16090_ (_07784_, _07783_);
  nor _16091_ (_07785_, _07750_, _07630_);
  and _16092_ (_07786_, _07757_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16093_ (_07787_, _07760_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16094_ (_07788_, _07787_, _07786_);
  nor _16095_ (_07789_, _07788_, _07785_);
  nor _16096_ (_07790_, _07789_, _07784_);
  nor _16097_ (_07791_, _07790_, _07782_);
  and _16098_ (_07793_, _07791_, _07773_);
  or _16099_ (_07794_, _07746_, _07783_);
  not _16100_ (_07796_, _07794_);
  not _16101_ (_07797_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _16102_ (_07799_, _07603_, _07797_);
  or _16103_ (_07800_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _16104_ (_07801_, _07800_, _07799_);
  and _16105_ (_07802_, _07801_, _07796_);
  not _16106_ (_07804_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _16107_ (_07805_, _07603_, _07804_);
  or _16108_ (_07806_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _16109_ (_07808_, _07806_, _07805_);
  and _16110_ (_07809_, _07808_, _07794_);
  or _16111_ (_07810_, _07809_, _07802_);
  and _16112_ (_07811_, _07810_, _07757_);
  and _16113_ (_07813_, _07749_, _07612_);
  not _16114_ (_07814_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _16115_ (_07815_, _07603_, _07814_);
  or _16116_ (_07816_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _16117_ (_07818_, _07816_, _07815_);
  and _16118_ (_07819_, _07818_, _07796_);
  not _16119_ (_07820_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _16120_ (_07821_, _07603_, _07820_);
  or _16121_ (_07823_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _16122_ (_07824_, _07823_, _07821_);
  and _16123_ (_07825_, _07824_, _07794_);
  or _16124_ (_07826_, _07825_, _07819_);
  and _16125_ (_07827_, _07826_, _07813_);
  or _16126_ (_07828_, _07827_, _07811_);
  not _16127_ (_07829_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _16128_ (_07830_, _07603_, _07829_);
  or _16129_ (_07831_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _16130_ (_07832_, _07831_, _07830_);
  and _16131_ (_07833_, _07832_, _07794_);
  not _16132_ (_07834_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _16133_ (_07835_, _07603_, _07834_);
  or _16134_ (_07836_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _16135_ (_07837_, _07836_, _07835_);
  and _16136_ (_07838_, _07837_, _07796_);
  or _16137_ (_07839_, _07838_, _07833_);
  and _16138_ (_07840_, _07839_, _07760_);
  and _16139_ (_07841_, _07749_, _07659_);
  not _16140_ (_07842_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _16141_ (_07843_, _07603_, _07842_);
  or _16142_ (_07844_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _16143_ (_07845_, _07844_, _07843_);
  and _16144_ (_07846_, _07845_, _07794_);
  not _16145_ (_07847_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand _16146_ (_07848_, _07603_, _07847_);
  or _16147_ (_07849_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _16148_ (_07850_, _07849_, _07848_);
  and _16149_ (_07851_, _07850_, _07796_);
  or _16150_ (_07852_, _07851_, _07846_);
  and _16151_ (_07853_, _07852_, _07841_);
  or _16152_ (_07854_, _07853_, _07840_);
  nor _16153_ (_07855_, _07854_, _07828_);
  nor _16154_ (_07856_, _07855_, _07793_);
  and _16155_ (_07857_, _07793_, word_in[15]);
  or _16156_ (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _07857_, _07856_);
  nor _16157_ (_07858_, _07644_, _07624_);
  not _16158_ (_07859_, _07858_);
  nor _16159_ (_07860_, _07859_, _07630_);
  and _16160_ (_07861_, _07644_, _07612_);
  nor _16161_ (_07862_, _07644_, _07612_);
  nor _16162_ (_07863_, _07862_, _07861_);
  and _16163_ (_07865_, _07863_, _07859_);
  and _16164_ (_07866_, _07865_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _16165_ (_07868_, _07863_, _07858_);
  and _16166_ (_07869_, _07868_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16167_ (_07870_, _07869_, _07866_);
  nor _16168_ (_07871_, _07870_, _07860_);
  nor _16169_ (_07872_, _07871_, _07766_);
  and _16170_ (_07873_, _07868_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not _16171_ (_07874_, _07873_);
  nor _16172_ (_07875_, _07859_, _07650_);
  and _16173_ (_07876_, _07865_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16174_ (_07877_, _07876_, _07875_);
  and _16175_ (_07879_, _07877_, _07874_);
  nor _16176_ (_07880_, _07879_, _07745_);
  nor _16177_ (_07881_, _07880_, _07872_);
  and _16178_ (_07882_, _07868_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not _16179_ (_07883_, _07882_);
  nor _16180_ (_07884_, _07859_, _07672_);
  and _16181_ (_07885_, _07865_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _16182_ (_07886_, _07885_, _07884_);
  and _16183_ (_07887_, _07886_, _07883_);
  nor _16184_ (_07888_, _07887_, _07784_);
  nor _16185_ (_07889_, _07859_, _07678_);
  and _16186_ (_07890_, _07865_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16187_ (_07891_, _07868_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _16188_ (_07892_, _07891_, _07890_);
  nor _16189_ (_07893_, _07892_, _07889_);
  nor _16190_ (_07894_, _07893_, _07776_);
  nor _16191_ (_07895_, _07894_, _07888_);
  and _16192_ (_07896_, _07895_, _07881_);
  and _16193_ (_07897_, _07896_, word_in[23]);
  and _16194_ (_07898_, _07730_, _07636_);
  and _16195_ (_07899_, _07719_, _07624_);
  or _16196_ (_07901_, _07899_, _07898_);
  and _16197_ (_07902_, _07724_, _07633_);
  and _16198_ (_07903_, _07735_, _07644_);
  or _16199_ (_07904_, _07903_, _07902_);
  or _16200_ (_07905_, _07904_, _07901_);
  or _16201_ (_07906_, _07905_, _07863_);
  not _16202_ (_07907_, _07863_);
  and _16203_ (_07908_, _07688_, _07633_);
  and _16204_ (_07909_, _07710_, _07659_);
  or _16205_ (_07910_, _07909_, _07908_);
  and _16206_ (_07912_, _07704_, _07636_);
  and _16207_ (_07913_, _07695_, _07624_);
  or _16208_ (_07914_, _07913_, _07912_);
  or _16209_ (_07916_, _07914_, _07910_);
  or _16210_ (_07917_, _07916_, _07907_);
  nand _16211_ (_07920_, _07917_, _07906_);
  nor _16212_ (_07921_, _07920_, _07896_);
  or _16213_ (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _07921_, _07897_);
  and _16214_ (_07923_, _07748_, _07612_);
  and _16215_ (_07925_, _07923_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _16216_ (_07926_, _07784_, _07623_);
  not _16217_ (_07927_, _07926_);
  nand _16218_ (_07929_, _07784_, _07623_);
  and _16219_ (_07930_, _07929_, _07927_);
  not _16220_ (_07931_, _07930_);
  nor _16221_ (_07933_, _07672_, _07931_);
  nor _16222_ (_07935_, _07929_, _07612_);
  and _16223_ (_07936_, _07929_, _07612_);
  nor _16224_ (_07937_, _07936_, _07935_);
  nor _16225_ (_07938_, _07937_, _07930_);
  and _16226_ (_07939_, _07938_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _16227_ (_07940_, _07939_, _07933_);
  nor _16228_ (_07941_, _07940_, _07766_);
  nor _16229_ (_07942_, _07678_, _07931_);
  and _16230_ (_07943_, _07938_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16231_ (_07944_, _07937_, _07931_);
  and _16232_ (_07945_, _07944_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _16233_ (_07946_, _07945_, _07943_);
  nor _16234_ (_07947_, _07946_, _07942_);
  nor _16235_ (_07948_, _07947_, _07745_);
  or _16236_ (_07949_, _07948_, _07941_);
  nor _16237_ (_07950_, _07949_, _07925_);
  and _16238_ (_07951_, _07930_, _07631_);
  and _16239_ (_07952_, _07944_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _16240_ (_07953_, _07938_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _16241_ (_07954_, _07953_, _07952_);
  nor _16242_ (_07955_, _07954_, _07951_);
  nor _16243_ (_07956_, _07955_, _07776_);
  nor _16244_ (_07957_, _07931_, _07650_);
  and _16245_ (_07958_, _07938_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16246_ (_07959_, _07958_, _07957_);
  nor _16247_ (_07960_, _07959_, _07784_);
  and _16248_ (_07961_, _07926_, _07640_);
  or _16249_ (_07962_, _07961_, _07960_);
  nor _16250_ (_07963_, _07962_, _07956_);
  and _16251_ (_07964_, _07963_, _07950_);
  and _16252_ (_07965_, _07808_, _07796_);
  and _16253_ (_07966_, _07801_, _07794_);
  or _16254_ (_07967_, _07966_, _07965_);
  and _16255_ (_07968_, _07967_, _07938_);
  and _16256_ (_07969_, _07832_, _07796_);
  and _16257_ (_07970_, _07837_, _07794_);
  or _16258_ (_07971_, _07970_, _07969_);
  and _16259_ (_07972_, _07971_, _07944_);
  and _16260_ (_07973_, _07930_, _07659_);
  and _16261_ (_07974_, _07845_, _07796_);
  and _16262_ (_07975_, _07850_, _07794_);
  or _16263_ (_07976_, _07975_, _07974_);
  and _16264_ (_07977_, _07976_, _07973_);
  and _16265_ (_07978_, _07824_, _07796_);
  and _16266_ (_07979_, _07818_, _07794_);
  or _16267_ (_07980_, _07979_, _07978_);
  and _16268_ (_07981_, _07936_, _07927_);
  and _16269_ (_07982_, _07981_, _07980_);
  or _16270_ (_07983_, _07982_, _07977_);
  or _16271_ (_07984_, _07983_, _07972_);
  nor _16272_ (_07985_, _07984_, _07968_);
  nor _16273_ (_07986_, _07985_, _07964_);
  and _16274_ (_07987_, _07964_, word_in[31]);
  or _16275_ (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _07987_, _07986_);
  and _16276_ (_07988_, _07612_, _07623_);
  nor _16277_ (_07989_, _07861_, _07647_);
  or _16278_ (_07990_, _07989_, _07988_);
  and _16279_ (_06013_, _07990_, _05110_);
  and _16280_ (_07992_, _07858_, _07612_);
  and _16281_ (_07993_, _07896_, _05110_);
  and _16282_ (_07995_, _07993_, _07744_);
  and _16283_ (_07996_, _07995_, _07992_);
  not _16284_ (_07998_, _07996_);
  and _16285_ (_07999_, _07793_, _05110_);
  and _16286_ (_08001_, _07999_, _07775_);
  and _16287_ (_08002_, _08001_, _07813_);
  and _16288_ (_08004_, _07656_, _05110_);
  and _16289_ (_08005_, _08004_, _07618_);
  nor _16290_ (_08007_, _07683_, rst);
  and _16291_ (_08008_, _08007_, _07988_);
  and _16292_ (_08010_, _08008_, _08005_);
  and _16293_ (_08011_, _08007_, word_in[7]);
  and _16294_ (_08013_, _08011_, _08010_);
  nor _16295_ (_08014_, _08010_, _07684_);
  nor _16296_ (_08015_, _08014_, _08013_);
  nor _16297_ (_08016_, _08015_, _08002_);
  and _16298_ (_08017_, _08002_, word_in[15]);
  or _16299_ (_08018_, _08017_, _08016_);
  and _16300_ (_08019_, _08018_, _07998_);
  and _16301_ (_08020_, _07988_, _07783_);
  and _16302_ (_08021_, _07964_, _05110_);
  and _16303_ (_08022_, _08021_, _08020_);
  and _16304_ (_08023_, _07993_, word_in[23]);
  and _16305_ (_08024_, _08023_, _07996_);
  or _16306_ (_08025_, _08024_, _08022_);
  or _16307_ (_08026_, _08025_, _08019_);
  not _16308_ (_08027_, _08022_);
  and _16309_ (_08028_, _08021_, word_in[31]);
  or _16310_ (_08029_, _08028_, _08027_);
  and _16311_ (_06039_, _08029_, _08026_);
  or _16312_ (_08030_, _07944_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _16313_ (_06060_, _08030_, _05110_);
  and _16314_ (_08031_, _07624_, _07659_);
  or _16315_ (_08032_, _08031_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _16316_ (_08033_, _08032_, _07861_);
  and _16317_ (_06090_, _08033_, _05110_);
  nor _16318_ (_08034_, _08031_, _07923_);
  or _16319_ (_08035_, _07745_, _07623_);
  nor _16320_ (_08036_, _08035_, _07612_);
  and _16321_ (_08037_, _07775_, _07973_);
  nor _16322_ (_08038_, _08037_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _16323_ (_08039_, _08038_, _08036_);
  nand _16324_ (_08040_, _08039_, _08034_);
  and _16325_ (_06133_, _08040_, _05110_);
  not _16326_ (_08041_, _07760_);
  and _16327_ (_08042_, _07746_, _07973_);
  or _16328_ (_08043_, _08042_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _16329_ (_08044_, _08043_, _08041_);
  and _16330_ (_08045_, _07624_, _07640_);
  or _16331_ (_08046_, _08045_, _08037_);
  or _16332_ (_08047_, _08046_, _08044_);
  and _16333_ (_08048_, _08047_, _08034_);
  and _16334_ (_08049_, _08043_, _07923_);
  or _16335_ (_08050_, _08049_, _08031_);
  or _16336_ (_08051_, _08050_, _08048_);
  and _16337_ (_06181_, _08051_, _05110_);
  not _16338_ (_08052_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _16339_ (_08053_, _06001_, _05337_);
  nor _16340_ (_08054_, _08053_, _08052_);
  not _16341_ (_08056_, _08053_);
  nor _16342_ (_08057_, _08056_, _06088_);
  or _16343_ (_08058_, _08057_, _08054_);
  and _16344_ (_06192_, _08058_, _05110_);
  and _16345_ (_08059_, _07754_, _07783_);
  or _16346_ (_08060_, _08059_, _08042_);
  or _16347_ (_08061_, _08060_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _16348_ (_08062_, _08061_, _08041_);
  and _16349_ (_08063_, _07926_, _07659_);
  or _16350_ (_08064_, _08063_, _07923_);
  and _16351_ (_08065_, _08064_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _16352_ (_08066_, _08065_, _08036_);
  or _16353_ (_08067_, _08066_, _08062_);
  or _16354_ (_08068_, _08067_, _08037_);
  and _16355_ (_06236_, _08068_, _05110_);
  nor _16356_ (_08069_, _08063_, _07973_);
  not _16357_ (_08070_, _07862_);
  or _16358_ (_08071_, _08070_, _08060_);
  and _16359_ (_08072_, _08071_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _16360_ (_08073_, _08037_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _16361_ (_08074_, _07744_, _07754_);
  and _16362_ (_08075_, _08031_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _16363_ (_08076_, _08075_, _08074_);
  or _16364_ (_08078_, _08076_, _08073_);
  or _16365_ (_08079_, _08078_, _08072_);
  and _16366_ (_08081_, _08079_, _08069_);
  and _16367_ (_08082_, _08063_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _16368_ (_08083_, _08036_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _16369_ (_08085_, _08083_, _08037_);
  or _16370_ (_08086_, _08085_, _08082_);
  or _16371_ (_08087_, _08086_, _08059_);
  or _16372_ (_08088_, _08087_, _08042_);
  or _16373_ (_08090_, _08088_, _08081_);
  and _16374_ (_06299_, _08090_, _05110_);
  or _16375_ (_08092_, _07752_, _07935_);
  and _16376_ (_08093_, _07644_, _07659_);
  or _16377_ (_08095_, _07752_, _08093_);
  and _16378_ (_08096_, _07775_, _07754_);
  or _16379_ (_08097_, _08096_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _16380_ (_08099_, _08097_, _08095_);
  and _16381_ (_08100_, _08060_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _16382_ (_08101_, _08100_, _08074_);
  or _16383_ (_08102_, _08101_, _08099_);
  and _16384_ (_08104_, _08102_, _08092_);
  and _16385_ (_08105_, _08097_, _07923_);
  and _16386_ (_08106_, _07670_, _07747_);
  or _16387_ (_08107_, _08106_, _08042_);
  or _16388_ (_08108_, _08107_, _08059_);
  or _16389_ (_08109_, _08108_, _08105_);
  or _16390_ (_08110_, _08109_, _08104_);
  and _16391_ (_06361_, _08110_, _05110_);
  not _16392_ (_08111_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor _16393_ (_08112_, _08053_, _08111_);
  nor _16394_ (_08113_, _08056_, _06229_);
  or _16395_ (_08114_, _08113_, _08112_);
  and _16396_ (_06372_, _08114_, _05110_);
  and _16397_ (_08115_, _08053_, _06559_);
  not _16398_ (_08116_, _06903_);
  or _16399_ (_08117_, _08116_, _06555_);
  and _16400_ (_08118_, _08117_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _16401_ (_08119_, _08118_, _08115_);
  and _16402_ (_06408_, _08119_, _05110_);
  or _16403_ (_08120_, _07748_, _07612_);
  or _16404_ (_08121_, _07755_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _16405_ (_08122_, _08121_, _08120_);
  and _16406_ (_08123_, _07973_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _16407_ (_08124_, _08063_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _16408_ (_08125_, _08124_, _08059_);
  or _16409_ (_08126_, _08125_, _08123_);
  or _16410_ (_08127_, _08126_, _08096_);
  or _16411_ (_08128_, _08127_, _08074_);
  or _16412_ (_08129_, _08128_, _08122_);
  and _16413_ (_06441_, _08129_, _05110_);
  nor _16414_ (_08130_, _06628_, _05591_);
  and _16415_ (_08131_, _06625_, _05794_);
  and _16416_ (_08132_, _08131_, _06626_);
  and _16417_ (_08133_, _05912_, _05485_);
  and _16418_ (_08134_, _08133_, _05782_);
  nor _16419_ (_08135_, _08133_, _05591_);
  or _16420_ (_08136_, _08135_, _08134_);
  nand _16421_ (_08137_, _08136_, _08132_);
  nand _16422_ (_08138_, _08137_, _06622_);
  or _16423_ (_08139_, _08138_, _08130_);
  and _16424_ (_08140_, _06623_, _06548_);
  nor _16425_ (_08141_, _08140_, _06613_);
  nand _16426_ (_08142_, _08141_, _08139_);
  nand _16427_ (_08143_, _07277_, _06613_);
  nand _16428_ (_08144_, _08143_, _08142_);
  and _16429_ (_06474_, _08144_, _05110_);
  nor _16430_ (_08145_, _07418_, _06622_);
  nor _16431_ (_08146_, _08145_, _06613_);
  and _16432_ (_08147_, _08132_, _05805_);
  nand _16433_ (_08148_, _08147_, _05872_);
  nor _16434_ (_08149_, _08147_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  not _16435_ (_08150_, _08149_);
  and _16436_ (_08151_, _08150_, _06638_);
  nand _16437_ (_08152_, _08151_, _08148_);
  nand _16438_ (_08153_, _08152_, _08146_);
  or _16439_ (_08154_, _07391_, _06637_);
  and _16440_ (_08155_, _08154_, _08153_);
  and _16441_ (_06484_, _08155_, _05110_);
  and _16442_ (_08156_, _07926_, _07612_);
  or _16443_ (_08157_, _08156_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16444_ (_08158_, _08157_, _07612_);
  or _16445_ (_08159_, _08031_, _07660_);
  and _16446_ (_08160_, _08159_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _16447_ (_08161_, _08059_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _16448_ (_08162_, _08074_, _07755_);
  or _16449_ (_08163_, _08162_, _08161_);
  or _16450_ (_08164_, _08163_, _08160_);
  or _16451_ (_08165_, _08164_, _08096_);
  or _16452_ (_08166_, _08165_, _08158_);
  and _16453_ (_06527_, _08166_, _05110_);
  and _16454_ (_08167_, _07752_, _07927_);
  nor _16455_ (_08168_, _08035_, _07659_);
  or _16456_ (_08169_, _08168_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16457_ (_08170_, _08169_, _08167_);
  or _16458_ (_08172_, _08170_, _08156_);
  and _16459_ (_08173_, _07862_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16460_ (_08174_, _08169_, _07923_);
  or _16461_ (_08176_, _08174_, _08093_);
  or _16462_ (_08177_, _08176_, _08173_);
  or _16463_ (_08178_, _08177_, _08172_);
  and _16464_ (_06614_, _08178_, _05110_);
  not _16465_ (_08179_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor _16466_ (_08180_, _08053_, _08179_);
  nor _16467_ (_08181_, _08056_, _05334_);
  or _16468_ (_08182_, _08181_, _08180_);
  and _16469_ (_06684_, _08182_, _05110_);
  and _16470_ (_08183_, _07752_, _07625_);
  or _16471_ (_08184_, _08183_, _07923_);
  and _16472_ (_08186_, _07796_, _07973_);
  and _16473_ (_08187_, _08186_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _16474_ (_08188_, _08156_, _07755_);
  and _16475_ (_08189_, _08188_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16476_ (_08190_, _07775_, _07936_);
  and _16477_ (_08191_, _08063_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _16478_ (_08192_, _08191_, _08190_);
  and _16479_ (_08193_, _07841_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand _16480_ (_08194_, _08035_, _07747_);
  and _16481_ (_08195_, _08194_, _07657_);
  or _16482_ (_08196_, _08195_, _08193_);
  or _16483_ (_08197_, _08196_, _08192_);
  or _16484_ (_08198_, _08197_, _08189_);
  or _16485_ (_08199_, _08198_, _08187_);
  and _16486_ (_08200_, _08199_, _08184_);
  or _16487_ (_08201_, _08189_, _08168_);
  or _16488_ (_08202_, _08201_, _08200_);
  and _16489_ (_08203_, _08202_, _08167_);
  and _16490_ (_08204_, _08199_, _07923_);
  or _16491_ (_08205_, _08204_, _07755_);
  not _16492_ (_08206_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _16493_ (_08207_, _08120_, _08206_);
  or _16494_ (_08208_, _08207_, _08156_);
  or _16495_ (_08209_, _08208_, _08205_);
  or _16496_ (_08210_, _08209_, _08203_);
  and _16497_ (_06715_, _08210_, _05110_);
  and _16498_ (_08211_, _07746_, _07936_);
  and _16499_ (_08212_, _07988_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _16500_ (_08213_, _08212_, _08211_);
  or _16501_ (_08214_, _08186_, _07755_);
  and _16502_ (_08215_, _08214_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _16503_ (_08216_, _07841_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _16504_ (_08217_, _07926_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _16505_ (_08218_, _08217_, _08156_);
  or _16506_ (_08219_, _08218_, _08216_);
  or _16507_ (_08220_, _08219_, _08215_);
  or _16508_ (_08221_, _08220_, _08168_);
  or _16509_ (_08222_, _08221_, _08190_);
  or _16510_ (_08223_, _08222_, _08213_);
  and _16511_ (_06806_, _08223_, _05110_);
  not _16512_ (_08224_, _05841_);
  and _16513_ (_08225_, _06184_, _08224_);
  not _16514_ (_08226_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor _16515_ (_08227_, _06184_, _08226_);
  or _16516_ (_08228_, _08227_, _08225_);
  and _16517_ (_06855_, _08228_, _05110_);
  or _16518_ (_08229_, _07926_, _07659_);
  and _16519_ (_08230_, _08229_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _16520_ (_08231_, _07988_, _07784_);
  and _16521_ (_08232_, _08231_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _16522_ (_08233_, _08232_, _07981_);
  or _16523_ (_08234_, _08233_, _08230_);
  and _16524_ (_06900_, _08234_, _05110_);
  nor _16525_ (_08235_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _16526_ (_08236_, _08235_);
  nor _16527_ (_08237_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _16528_ (_08238_, _08237_, _08236_);
  and _16529_ (_08239_, _08238_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not _16530_ (_08240_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor _16531_ (_08241_, _08238_, _08240_);
  or _16532_ (_08242_, _08241_, _08239_);
  and _16533_ (_08243_, _06152_, _05789_);
  or _16534_ (_08244_, _08243_, _08242_);
  and _16535_ (_08245_, _06472_, _05782_);
  or _16536_ (_08246_, _06472_, _08240_);
  nand _16537_ (_08248_, _08246_, _08243_);
  or _16538_ (_08249_, _08248_, _08245_);
  and _16539_ (_08251_, _08249_, _08244_);
  and _16540_ (_08252_, _05803_, _05434_);
  and _16541_ (_08253_, _08252_, _05808_);
  or _16542_ (_08254_, _08253_, _08251_);
  nand _16543_ (_08255_, _08253_, _06229_);
  and _16544_ (_08256_, _08255_, _05110_);
  and _16545_ (_06961_, _08256_, _08254_);
  and _16546_ (_08257_, _07206_, _05867_);
  or _16547_ (_08258_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _16548_ (_08259_, _08258_, _05110_);
  nand _16549_ (_08260_, _08257_, _05334_);
  and _16550_ (_06965_, _08260_, _08259_);
  or _16551_ (_08261_, _07992_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _16552_ (_06995_, _08261_, _05110_);
  and _16553_ (_08262_, _05806_, _05403_);
  and _16554_ (_08263_, _08252_, _08262_);
  and _16555_ (_08264_, _08243_, _08133_);
  nand _16556_ (_08265_, _08264_, _05872_);
  or _16557_ (_08266_, _08264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _16558_ (_08267_, _08266_, _08265_);
  or _16559_ (_08268_, _08267_, _08263_);
  nand _16560_ (_08269_, _08253_, _06054_);
  and _16561_ (_08270_, _08269_, _05110_);
  and _16562_ (_07022_, _08270_, _08268_);
  and _16563_ (_08272_, _06173_, _05911_);
  and _16564_ (_08273_, _05807_, _08272_);
  and _16565_ (_08274_, _08273_, _08252_);
  and _16566_ (_08276_, _08274_, _08236_);
  and _16567_ (_08277_, _08276_, _06799_);
  and _16568_ (_08278_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _16569_ (_08280_, _08278_, _08235_);
  and _16570_ (_08281_, _08236_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _16571_ (_08282_, _08281_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _16572_ (_08283_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _16573_ (_08285_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _16574_ (_08286_, _08285_, _08283_);
  and _16575_ (_08287_, _08286_, _08282_);
  nor _16576_ (_08288_, _08287_, _08280_);
  not _16577_ (_08290_, _08288_);
  and _16578_ (_08291_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _16579_ (_08292_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _16580_ (_08293_, _08292_, _08291_);
  nor _16581_ (_08296_, _08293_, _08274_);
  and _16582_ (_08297_, _08274_, _08235_);
  and _16583_ (_08298_, _08297_, _06559_);
  or _16584_ (_08300_, _08298_, _08296_);
  or _16585_ (_08301_, _08300_, _08277_);
  and _16586_ (_07036_, _08301_, _05110_);
  and _16587_ (_08302_, _07305_, _06613_);
  nor _16588_ (_08303_, _07337_, _06622_);
  and _16589_ (_08304_, _08132_, _06472_);
  nand _16590_ (_08305_, _08304_, _05872_);
  nor _16591_ (_08306_, _08304_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not _16592_ (_08307_, _08306_);
  and _16593_ (_08308_, _08307_, _06638_);
  and _16594_ (_08309_, _08308_, _08305_);
  or _16595_ (_08310_, _08309_, _08303_);
  and _16596_ (_08311_, _08310_, _06637_);
  or _16597_ (_08312_, _08311_, _08302_);
  and _16598_ (_07042_, _08312_, _05110_);
  and _16599_ (_08313_, _08243_, _05488_);
  nand _16600_ (_08314_, _08313_, _05872_);
  or _16601_ (_08315_, _08313_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _16602_ (_08316_, _08315_, _08314_);
  or _16603_ (_08317_, _08316_, _08263_);
  nand _16604_ (_08318_, _08253_, _05841_);
  and _16605_ (_08319_, _08318_, _05110_);
  and _16606_ (_07047_, _08319_, _08317_);
  nor _16607_ (_08320_, _05901_, _05465_);
  not _16608_ (_08321_, _06174_);
  and _16609_ (_08322_, _08321_, _06170_);
  and _16610_ (_08323_, _08322_, _06168_);
  or _16611_ (_08324_, _08323_, _05995_);
  not _16612_ (_08325_, _06001_);
  nand _16613_ (_08326_, _08325_, _06170_);
  nand _16614_ (_08327_, _08326_, _05337_);
  nand _16615_ (_08328_, _08327_, _06554_);
  or _16616_ (_08329_, _08328_, _08324_);
  and _16617_ (_08330_, _08329_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  or _16618_ (_08331_, _08330_, _08320_);
  and _16619_ (_07102_, _08331_, _05110_);
  or _16620_ (_08332_, _07813_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _16621_ (_07112_, _08332_, _05110_);
  nor _16622_ (_08333_, _06229_, _06010_);
  not _16623_ (_08334_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor _16624_ (_08335_, _05997_, _08334_);
  or _16625_ (_08336_, _08335_, _05995_);
  or _16626_ (_08337_, _08336_, _08333_);
  or _16627_ (_08338_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _16628_ (_08339_, _08338_, _05110_);
  and _16629_ (_07166_, _08339_, _08337_);
  and _16630_ (_08340_, _08282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  or _16631_ (_08341_, _08340_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _16632_ (_08342_, _08340_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _16633_ (_08343_, _08342_, rst);
  nand _16634_ (_08344_, _08343_, _08341_);
  nor _16635_ (_07175_, _08344_, _08274_);
  or _16636_ (_08345_, _08282_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _16637_ (_08346_, _08340_, rst);
  nand _16638_ (_08347_, _08346_, _08345_);
  nor _16639_ (_07189_, _08347_, _08274_);
  and _16640_ (_08348_, _07999_, _07923_);
  not _16641_ (_08349_, _08348_);
  not _16642_ (_08350_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _16643_ (_08351_, _08007_, _07618_);
  nor _16644_ (_08352_, _08351_, _08004_);
  and _16645_ (_08353_, _08007_, _07623_);
  and _16646_ (_08354_, _08007_, _07612_);
  nor _16647_ (_08355_, _08354_, _08353_);
  and _16648_ (_08356_, _08355_, _08007_);
  and _16649_ (_08357_, _08356_, _08352_);
  nor _16650_ (_08358_, _08357_, _08350_);
  and _16651_ (_08359_, _08357_, word_in[0]);
  or _16652_ (_08360_, _08359_, _08358_);
  and _16653_ (_08361_, _08360_, _08349_);
  and _16654_ (_08362_, _08348_, word_in[8]);
  or _16655_ (_08363_, _08362_, _08361_);
  and _16656_ (_08364_, _07988_, _07775_);
  and _16657_ (_08365_, _07993_, _08364_);
  not _16658_ (_08366_, _08365_);
  and _16659_ (_08367_, _08366_, _08363_);
  and _16660_ (_08368_, _07988_, _07744_);
  and _16661_ (_08369_, _08021_, _08368_);
  and _16662_ (_08370_, _07993_, word_in[16]);
  and _16663_ (_08371_, _08370_, _08364_);
  or _16664_ (_08372_, _08371_, _08369_);
  or _16665_ (_08373_, _08372_, _08367_);
  not _16666_ (_08375_, _08369_);
  or _16667_ (_08376_, _08375_, word_in[24]);
  and _16668_ (_07468_, _08376_, _08373_);
  or _16669_ (_08378_, _08357_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  not _16670_ (_08379_, word_in[1]);
  nand _16671_ (_08381_, _08357_, _08379_);
  and _16672_ (_08383_, _08381_, _08349_);
  and _16673_ (_08384_, _08383_, _08378_);
  and _16674_ (_08385_, _07923_, word_in[9]);
  and _16675_ (_08387_, _08385_, _07999_);
  or _16676_ (_08388_, _08387_, _08365_);
  or _16677_ (_08390_, _08388_, _08384_);
  nor _16678_ (_08391_, _08366_, word_in[17]);
  nor _16679_ (_08393_, _08391_, _08369_);
  and _16680_ (_08394_, _08393_, _08390_);
  and _16681_ (_08395_, _08021_, word_in[25]);
  and _16682_ (_08397_, _08395_, _08369_);
  or _16683_ (_07472_, _08397_, _08394_);
  not _16684_ (_08398_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _16685_ (_08400_, _08357_, _08398_);
  and _16686_ (_08401_, _08007_, word_in[2]);
  and _16687_ (_08402_, _08401_, _08357_);
  or _16688_ (_08403_, _08402_, _08400_);
  or _16689_ (_08404_, _08403_, _08348_);
  or _16690_ (_08405_, _08349_, word_in[10]);
  and _16691_ (_08406_, _08405_, _08404_);
  or _16692_ (_08407_, _08406_, _08365_);
  nor _16693_ (_08408_, _08366_, word_in[18]);
  nor _16694_ (_08409_, _08408_, _08369_);
  and _16695_ (_08410_, _08409_, _08407_);
  and _16696_ (_08411_, _08021_, word_in[26]);
  and _16697_ (_08412_, _08411_, _08369_);
  or _16698_ (_07476_, _08412_, _08410_);
  not _16699_ (_08413_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _16700_ (_08414_, _08357_, _08413_);
  and _16701_ (_08415_, _08007_, word_in[3]);
  and _16702_ (_08416_, _08415_, _08357_);
  or _16703_ (_08417_, _08416_, _08414_);
  or _16704_ (_08418_, _08417_, _08348_);
  or _16705_ (_08419_, _08349_, word_in[11]);
  and _16706_ (_08420_, _08419_, _08418_);
  or _16707_ (_08421_, _08420_, _08365_);
  nor _16708_ (_08422_, _08366_, word_in[19]);
  nor _16709_ (_08423_, _08422_, _08369_);
  and _16710_ (_08424_, _08423_, _08421_);
  and _16711_ (_08425_, _08021_, word_in[27]);
  and _16712_ (_08426_, _08425_, _08369_);
  or _16713_ (_07481_, _08426_, _08424_);
  not _16714_ (_08427_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _16715_ (_08428_, _08357_, _08427_);
  and _16716_ (_08429_, _08007_, word_in[4]);
  and _16717_ (_08430_, _08429_, _08357_);
  or _16718_ (_08431_, _08430_, _08428_);
  and _16719_ (_08432_, _08431_, _08349_);
  and _16720_ (_08433_, _08348_, word_in[12]);
  or _16721_ (_08434_, _08433_, _08432_);
  or _16722_ (_08435_, _08434_, _08365_);
  nor _16723_ (_08436_, _08366_, word_in[20]);
  nor _16724_ (_08437_, _08436_, _08369_);
  and _16725_ (_08438_, _08437_, _08435_);
  and _16726_ (_08439_, _08021_, word_in[28]);
  and _16727_ (_08440_, _08439_, _08369_);
  or _16728_ (_07484_, _08440_, _08438_);
  not _16729_ (_08441_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _16730_ (_08442_, _08357_, _08441_);
  and _16731_ (_08443_, _08007_, word_in[5]);
  and _16732_ (_08444_, _08443_, _08357_);
  or _16733_ (_08445_, _08444_, _08442_);
  or _16734_ (_08446_, _08445_, _08348_);
  or _16735_ (_08447_, _08349_, word_in[13]);
  and _16736_ (_08448_, _08447_, _08446_);
  or _16737_ (_08449_, _08448_, _08365_);
  nor _16738_ (_08450_, _08366_, word_in[21]);
  nor _16739_ (_08451_, _08450_, _08369_);
  and _16740_ (_08452_, _08451_, _08449_);
  and _16741_ (_08453_, _08021_, word_in[29]);
  and _16742_ (_08454_, _08453_, _08369_);
  or _16743_ (_07488_, _08454_, _08452_);
  not _16744_ (_08455_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _16745_ (_08456_, _08357_, _08455_);
  and _16746_ (_08457_, _08007_, word_in[6]);
  and _16747_ (_08458_, _08457_, _08357_);
  or _16748_ (_08459_, _08458_, _08456_);
  or _16749_ (_08460_, _08459_, _08348_);
  or _16750_ (_08461_, _08349_, word_in[14]);
  and _16751_ (_08462_, _08461_, _08460_);
  or _16752_ (_08463_, _08462_, _08365_);
  nor _16753_ (_08464_, _08366_, word_in[22]);
  nor _16754_ (_08466_, _08464_, _08369_);
  and _16755_ (_08467_, _08466_, _08463_);
  and _16756_ (_08469_, _08021_, word_in[30]);
  and _16757_ (_08470_, _08469_, _08369_);
  or _16758_ (_07491_, _08470_, _08467_);
  and _16759_ (_08471_, _08369_, word_in[31]);
  nor _16760_ (_08473_, _08357_, _07829_);
  and _16761_ (_08474_, _08357_, word_in[7]);
  or _16762_ (_08476_, _08474_, _08473_);
  and _16763_ (_08478_, _08476_, _08349_);
  and _16764_ (_08480_, _08348_, word_in[15]);
  or _16765_ (_08481_, _08480_, _08478_);
  or _16766_ (_08483_, _08481_, _08365_);
  nor _16767_ (_08484_, _08366_, word_in[23]);
  nor _16768_ (_08486_, _08484_, _08369_);
  and _16769_ (_08487_, _08486_, _08483_);
  or _16770_ (_07495_, _08487_, _08471_);
  and _16771_ (_08488_, _08021_, _08364_);
  not _16772_ (_08489_, _08488_);
  and _16773_ (_08490_, _07993_, _07746_);
  and _16774_ (_08491_, _08490_, _07868_);
  and _16775_ (_08492_, _08491_, _08370_);
  and _16776_ (_08493_, _07999_, _07783_);
  and _16777_ (_08494_, _08493_, _07760_);
  and _16778_ (_08495_, _08007_, word_in[0]);
  and _16779_ (_08496_, _08004_, _07632_);
  and _16780_ (_08497_, _08496_, _08355_);
  and _16781_ (_08498_, _08497_, _08495_);
  not _16782_ (_08499_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor _16783_ (_08500_, _08497_, _08499_);
  or _16784_ (_08501_, _08500_, _08498_);
  or _16785_ (_08502_, _08501_, _08494_);
  not _16786_ (_08503_, _08491_);
  not _16787_ (_08504_, _08494_);
  or _16788_ (_08505_, _08504_, word_in[8]);
  and _16789_ (_08506_, _08505_, _08503_);
  and _16790_ (_08507_, _08506_, _08502_);
  or _16791_ (_08508_, _08507_, _08492_);
  and _16792_ (_08509_, _08508_, _08489_);
  and _16793_ (_08510_, _08488_, word_in[24]);
  or _16794_ (_07573_, _08510_, _08509_);
  and _16795_ (_08511_, _07993_, word_in[17]);
  and _16796_ (_08512_, _08491_, _08511_);
  and _16797_ (_08513_, _08007_, word_in[1]);
  and _16798_ (_08514_, _08497_, _08513_);
  not _16799_ (_08515_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _16800_ (_08516_, _08497_, _08515_);
  nor _16801_ (_08517_, _08516_, _08514_);
  nor _16802_ (_08518_, _08517_, _08494_);
  and _16803_ (_08519_, _08494_, word_in[9]);
  or _16804_ (_08520_, _08519_, _08518_);
  and _16805_ (_08521_, _08520_, _08503_);
  or _16806_ (_08522_, _08521_, _08512_);
  and _16807_ (_08523_, _08522_, _08489_);
  and _16808_ (_08524_, _08488_, word_in[25]);
  or _16809_ (_07577_, _08524_, _08523_);
  and _16810_ (_08525_, _07993_, word_in[18]);
  and _16811_ (_08526_, _08491_, _08525_);
  and _16812_ (_08527_, _08497_, _08401_);
  not _16813_ (_08528_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _16814_ (_08529_, _08497_, _08528_);
  or _16815_ (_08530_, _08529_, _08527_);
  or _16816_ (_08531_, _08530_, _08494_);
  or _16817_ (_08532_, _08504_, word_in[10]);
  and _16818_ (_08533_, _08532_, _08503_);
  and _16819_ (_08534_, _08533_, _08531_);
  or _16820_ (_08535_, _08534_, _08526_);
  and _16821_ (_08536_, _08535_, _08489_);
  and _16822_ (_08537_, _08488_, word_in[26]);
  or _16823_ (_07581_, _08537_, _08536_);
  not _16824_ (_08538_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _16825_ (_08539_, _08497_, _08538_);
  and _16826_ (_08540_, _08497_, _08415_);
  or _16827_ (_08541_, _08540_, _08539_);
  or _16828_ (_08542_, _08541_, _08494_);
  or _16829_ (_08543_, _08504_, word_in[11]);
  and _16830_ (_08544_, _08543_, _08542_);
  or _16831_ (_08545_, _08544_, _08491_);
  and _16832_ (_08546_, _07993_, word_in[19]);
  or _16833_ (_08547_, _08503_, _08546_);
  and _16834_ (_08548_, _08547_, _08489_);
  and _16835_ (_08549_, _08548_, _08545_);
  and _16836_ (_08551_, _08488_, word_in[27]);
  or _16837_ (_07584_, _08551_, _08549_);
  not _16838_ (_08553_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _16839_ (_08554_, _08497_, _08553_);
  and _16840_ (_08555_, _08497_, _08429_);
  or _16841_ (_08557_, _08555_, _08554_);
  or _16842_ (_08558_, _08557_, _08494_);
  or _16843_ (_08560_, _08504_, word_in[12]);
  and _16844_ (_08561_, _08560_, _08558_);
  or _16845_ (_08563_, _08561_, _08491_);
  and _16846_ (_08564_, _07993_, word_in[20]);
  or _16847_ (_08565_, _08503_, _08564_);
  and _16848_ (_08567_, _08565_, _08489_);
  and _16849_ (_08569_, _08567_, _08563_);
  and _16850_ (_08570_, _08488_, word_in[28]);
  or _16851_ (_07587_, _08570_, _08569_);
  and _16852_ (_08572_, _07993_, word_in[21]);
  and _16853_ (_08573_, _08491_, _08572_);
  and _16854_ (_08574_, _08497_, _08443_);
  not _16855_ (_08575_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _16856_ (_08576_, _08497_, _08575_);
  nor _16857_ (_08577_, _08576_, _08574_);
  nor _16858_ (_08578_, _08577_, _08494_);
  and _16859_ (_08579_, _08494_, word_in[13]);
  or _16860_ (_08580_, _08579_, _08578_);
  and _16861_ (_08581_, _08580_, _08503_);
  or _16862_ (_08582_, _08581_, _08573_);
  and _16863_ (_08583_, _08582_, _08489_);
  and _16864_ (_08584_, _08488_, word_in[29]);
  or _16865_ (_07590_, _08584_, _08583_);
  not _16866_ (_08585_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _16867_ (_08586_, _08497_, _08585_);
  and _16868_ (_08587_, _08497_, _08457_);
  or _16869_ (_08588_, _08587_, _08586_);
  or _16870_ (_08589_, _08588_, _08494_);
  or _16871_ (_08590_, _08504_, word_in[14]);
  and _16872_ (_08591_, _08590_, _08589_);
  or _16873_ (_08592_, _08591_, _08491_);
  and _16874_ (_08593_, _07993_, word_in[22]);
  or _16875_ (_08594_, _08503_, _08593_);
  and _16876_ (_08595_, _08594_, _08489_);
  and _16877_ (_08596_, _08595_, _08592_);
  and _16878_ (_08597_, _08488_, word_in[30]);
  or _16879_ (_07593_, _08597_, _08596_);
  and _16880_ (_08598_, _08491_, _08023_);
  and _16881_ (_08599_, _08497_, _08011_);
  nor _16882_ (_08600_, _08497_, _07732_);
  or _16883_ (_08601_, _08600_, _08599_);
  or _16884_ (_08602_, _08601_, _08494_);
  or _16885_ (_08603_, _08504_, word_in[15]);
  and _16886_ (_08604_, _08603_, _08503_);
  and _16887_ (_08605_, _08604_, _08602_);
  or _16888_ (_08606_, _08605_, _08598_);
  and _16889_ (_08607_, _08606_, _08489_);
  and _16890_ (_08608_, _08488_, word_in[31]);
  or _16891_ (_07597_, _08608_, _08607_);
  and _16892_ (_08609_, _06559_, _05464_);
  and _16893_ (_08610_, _08329_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  or _16894_ (_08611_, _08610_, _08609_);
  and _16895_ (_07639_, _08611_, _05110_);
  not _16896_ (_08612_, _06004_);
  nand _16897_ (_08613_, _05998_, _05337_);
  or _16898_ (_08614_, _08613_, _08322_);
  or _16899_ (_08615_, _08614_, _08612_);
  and _16900_ (_08616_, _08615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and _16901_ (_08617_, _06169_, _05337_);
  and _16902_ (_08618_, _08617_, _06194_);
  or _16903_ (_08619_, _08618_, _08616_);
  and _16904_ (_07648_, _08619_, _05110_);
  and _16905_ (_08620_, _08614_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _16906_ (_08621_, _08617_, _06559_);
  nand _16907_ (_08622_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor _16908_ (_08623_, _08622_, _06004_);
  or _16909_ (_08624_, _08623_, _08621_);
  or _16910_ (_08625_, _08624_, _08620_);
  and _16911_ (_07653_, _08625_, _05110_);
  not _16912_ (_08626_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor _16913_ (_08627_, _05464_, _08626_);
  nor _16914_ (_08628_, _06088_, _05465_);
  or _16915_ (_08629_, _08628_, _08627_);
  and _16916_ (_07665_, _08629_, _05110_);
  and _16917_ (_08630_, _07999_, _07744_);
  and _16918_ (_08631_, _08630_, _07760_);
  not _16919_ (_08632_, _08004_);
  and _16920_ (_08633_, _08351_, _08632_);
  and _16921_ (_08634_, _08633_, _08355_);
  and _16922_ (_08635_, _08634_, _08495_);
  not _16923_ (_08637_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor _16924_ (_08638_, _08634_, _08637_);
  or _16925_ (_08639_, _08638_, _08635_);
  or _16926_ (_08641_, _08639_, _08631_);
  and _16927_ (_08642_, _07993_, _07783_);
  and _16928_ (_08643_, _08642_, _07868_);
  not _16929_ (_08644_, _08643_);
  not _16930_ (_08646_, _08631_);
  or _16931_ (_08647_, _08646_, word_in[8]);
  and _16932_ (_08648_, _08647_, _08644_);
  and _16933_ (_08649_, _08648_, _08641_);
  and _16934_ (_08651_, _08021_, _07746_);
  and _16935_ (_08652_, _08651_, _07944_);
  and _16936_ (_08653_, _08643_, _08370_);
  or _16937_ (_08654_, _08653_, _08652_);
  or _16938_ (_08655_, _08654_, _08649_);
  not _16939_ (_08656_, _08652_);
  or _16940_ (_08657_, _08656_, word_in[24]);
  and _16941_ (_07686_, _08657_, _08655_);
  and _16942_ (_08658_, _08634_, _08513_);
  not _16943_ (_08659_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _16944_ (_08660_, _08634_, _08659_);
  or _16945_ (_08661_, _08660_, _08658_);
  or _16946_ (_08662_, _08661_, _08631_);
  or _16947_ (_08663_, _08646_, word_in[9]);
  and _16948_ (_08664_, _08663_, _08644_);
  and _16949_ (_08665_, _08664_, _08662_);
  and _16950_ (_08666_, _08643_, _08511_);
  or _16951_ (_08667_, _08666_, _08652_);
  or _16952_ (_08668_, _08667_, _08665_);
  or _16953_ (_08669_, _08656_, word_in[25]);
  and _16954_ (_07689_, _08669_, _08668_);
  and _16955_ (_08670_, _08634_, _08401_);
  not _16956_ (_08671_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _16957_ (_08672_, _08634_, _08671_);
  or _16958_ (_08673_, _08672_, _08670_);
  or _16959_ (_08674_, _08673_, _08631_);
  or _16960_ (_08675_, _08646_, word_in[10]);
  and _16961_ (_08676_, _08675_, _08644_);
  and _16962_ (_08677_, _08676_, _08674_);
  and _16963_ (_08678_, _08643_, _08525_);
  or _16964_ (_08679_, _08678_, _08652_);
  or _16965_ (_08680_, _08679_, _08677_);
  or _16966_ (_08681_, _08656_, word_in[26]);
  and _16967_ (_07692_, _08681_, _08680_);
  and _16968_ (_08682_, _08634_, _08415_);
  not _16969_ (_08683_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _16970_ (_08684_, _08634_, _08683_);
  or _16971_ (_08685_, _08684_, _08682_);
  or _16972_ (_08686_, _08685_, _08631_);
  or _16973_ (_08687_, _08646_, word_in[11]);
  and _16974_ (_08688_, _08687_, _08644_);
  and _16975_ (_08689_, _08688_, _08686_);
  and _16976_ (_08690_, _08643_, _08546_);
  or _16977_ (_08691_, _08690_, _08652_);
  or _16978_ (_08692_, _08691_, _08689_);
  or _16979_ (_08693_, _08656_, word_in[27]);
  and _16980_ (_07697_, _08693_, _08692_);
  and _16981_ (_08694_, _08643_, _08564_);
  and _16982_ (_08695_, _08634_, _08429_);
  not _16983_ (_08696_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _16984_ (_08697_, _08634_, _08696_);
  nor _16985_ (_08698_, _08697_, _08695_);
  nor _16986_ (_08699_, _08698_, _08631_);
  and _16987_ (_08700_, _08631_, word_in[12]);
  or _16988_ (_08701_, _08700_, _08699_);
  and _16989_ (_08702_, _08701_, _08644_);
  or _16990_ (_08703_, _08702_, _08694_);
  and _16991_ (_08704_, _08703_, _08656_);
  and _16992_ (_08705_, _08652_, word_in[28]);
  or _16993_ (_07700_, _08705_, _08704_);
  and _16994_ (_08706_, _08643_, _08572_);
  and _16995_ (_08707_, _08634_, _08443_);
  not _16996_ (_08708_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _16997_ (_08709_, _08634_, _08708_);
  or _16998_ (_08710_, _08709_, _08707_);
  or _16999_ (_08711_, _08710_, _08631_);
  or _17000_ (_08712_, _08646_, word_in[13]);
  and _17001_ (_08713_, _08712_, _08644_);
  and _17002_ (_08714_, _08713_, _08711_);
  or _17003_ (_08715_, _08714_, _08706_);
  and _17004_ (_08716_, _08715_, _08656_);
  and _17005_ (_08717_, _08652_, word_in[29]);
  or _17006_ (_07703_, _08717_, _08716_);
  not _17007_ (_08718_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _17008_ (_08719_, _08634_, _08718_);
  and _17009_ (_08720_, _08634_, _08457_);
  or _17010_ (_08721_, _08720_, _08719_);
  or _17011_ (_08722_, _08721_, _08631_);
  or _17012_ (_08723_, _08646_, word_in[14]);
  and _17013_ (_08724_, _08723_, _08722_);
  or _17014_ (_08725_, _08724_, _08643_);
  nor _17015_ (_08726_, _08644_, _08593_);
  nor _17016_ (_08727_, _08726_, _08652_);
  and _17017_ (_08728_, _08727_, _08725_);
  and _17018_ (_08729_, _08652_, word_in[30]);
  or _17019_ (_07708_, _08729_, _08728_);
  and _17020_ (_08730_, _08643_, _08023_);
  and _17021_ (_08731_, _08634_, _08011_);
  nor _17022_ (_08732_, _08634_, _07834_);
  or _17023_ (_08733_, _08732_, _08731_);
  or _17024_ (_08734_, _08733_, _08631_);
  or _17025_ (_08735_, _08646_, word_in[15]);
  and _17026_ (_08736_, _08735_, _08644_);
  and _17027_ (_08737_, _08736_, _08734_);
  or _17028_ (_08738_, _08737_, _08730_);
  and _17029_ (_08739_, _08738_, _08656_);
  and _17030_ (_08740_, _08652_, word_in[31]);
  or _17031_ (_07713_, _08740_, _08739_);
  not _17032_ (_08741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not _17033_ (_08742_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor _17034_ (_08743_, _08235_, _08742_);
  and _17035_ (_08745_, _08743_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and _17036_ (_08746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _17037_ (_08748_, _08746_, _08236_);
  nor _17038_ (_08749_, _08748_, _08745_);
  or _17039_ (_08750_, _08749_, _08741_);
  and _17040_ (_08751_, _08750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _17041_ (_08752_, _08745_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _17042_ (_08753_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _17043_ (_08754_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _17044_ (_08755_, _08754_, _08753_);
  and _17045_ (_08756_, _08755_, _08752_);
  or _17046_ (_08757_, _08756_, _08751_);
  and _17047_ (_07758_, _08757_, _05110_);
  and _17048_ (_08758_, _08021_, _08063_);
  not _17049_ (_08759_, _08758_);
  and _17050_ (_08760_, _07995_, _07868_);
  and _17051_ (_08761_, _08760_, _08370_);
  and _17052_ (_08762_, _08001_, _07760_);
  and _17053_ (_08763_, _08355_, _08005_);
  and _17054_ (_08764_, _08763_, _08495_);
  not _17055_ (_08765_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor _17056_ (_08766_, _08763_, _08765_);
  or _17057_ (_08767_, _08766_, _08764_);
  or _17058_ (_08768_, _08767_, _08762_);
  not _17059_ (_08769_, _08760_);
  not _17060_ (_08770_, _08762_);
  or _17061_ (_08771_, _08770_, word_in[8]);
  and _17062_ (_08772_, _08771_, _08769_);
  and _17063_ (_08773_, _08772_, _08768_);
  or _17064_ (_08774_, _08773_, _08761_);
  and _17065_ (_08775_, _08774_, _08759_);
  and _17066_ (_08776_, _08758_, word_in[24]);
  or _17067_ (_07792_, _08776_, _08775_);
  and _17068_ (_08777_, _08760_, _08511_);
  and _17069_ (_08778_, _08763_, _08513_);
  not _17070_ (_08779_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _17071_ (_08780_, _08763_, _08779_);
  or _17072_ (_08781_, _08780_, _08778_);
  or _17073_ (_08782_, _08781_, _08762_);
  or _17074_ (_08783_, _08770_, word_in[9]);
  and _17075_ (_08784_, _08783_, _08769_);
  and _17076_ (_08785_, _08784_, _08782_);
  or _17077_ (_08786_, _08785_, _08777_);
  and _17078_ (_08787_, _08786_, _08759_);
  and _17079_ (_08788_, _08758_, word_in[25]);
  or _17080_ (_07795_, _08788_, _08787_);
  and _17081_ (_08789_, _08760_, _08525_);
  and _17082_ (_08790_, _08763_, _08401_);
  not _17083_ (_08791_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _17084_ (_08792_, _08763_, _08791_);
  or _17085_ (_08793_, _08792_, _08790_);
  or _17086_ (_08794_, _08793_, _08762_);
  or _17087_ (_08795_, _08770_, word_in[10]);
  and _17088_ (_08796_, _08795_, _08769_);
  and _17089_ (_08797_, _08796_, _08794_);
  or _17090_ (_08798_, _08797_, _08789_);
  and _17091_ (_08799_, _08798_, _08759_);
  and _17092_ (_08800_, _08758_, word_in[26]);
  or _17093_ (_07798_, _08800_, _08799_);
  and _17094_ (_08801_, _08760_, _08546_);
  and _17095_ (_08802_, _08763_, _08415_);
  not _17096_ (_08803_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _17097_ (_08804_, _08763_, _08803_);
  or _17098_ (_08805_, _08804_, _08802_);
  or _17099_ (_08806_, _08805_, _08762_);
  or _17100_ (_08807_, _08770_, word_in[11]);
  and _17101_ (_08808_, _08807_, _08769_);
  and _17102_ (_08809_, _08808_, _08806_);
  or _17103_ (_08810_, _08809_, _08801_);
  and _17104_ (_08811_, _08810_, _08759_);
  and _17105_ (_08812_, _08758_, word_in[27]);
  or _17106_ (_07803_, _08812_, _08811_);
  and _17107_ (_08813_, _08760_, _08564_);
  and _17108_ (_08814_, _08763_, _08429_);
  not _17109_ (_08815_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _17110_ (_08816_, _08763_, _08815_);
  or _17111_ (_08817_, _08816_, _08814_);
  or _17112_ (_08818_, _08817_, _08762_);
  or _17113_ (_08819_, _08770_, word_in[12]);
  and _17114_ (_08820_, _08819_, _08769_);
  and _17115_ (_08821_, _08820_, _08818_);
  or _17116_ (_08822_, _08821_, _08813_);
  and _17117_ (_08824_, _08822_, _08759_);
  and _17118_ (_08825_, _08758_, word_in[28]);
  or _17119_ (_07807_, _08825_, _08824_);
  and _17120_ (_08827_, _08760_, _08572_);
  and _17121_ (_08828_, _08763_, _08443_);
  not _17122_ (_08830_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _17123_ (_08831_, _08763_, _08830_);
  or _17124_ (_08833_, _08831_, _08828_);
  or _17125_ (_08834_, _08833_, _08762_);
  or _17126_ (_08836_, _08770_, word_in[13]);
  and _17127_ (_08837_, _08836_, _08769_);
  and _17128_ (_08838_, _08837_, _08834_);
  or _17129_ (_08840_, _08838_, _08827_);
  and _17130_ (_08841_, _08840_, _08759_);
  and _17131_ (_08842_, _08758_, word_in[29]);
  or _17132_ (_07812_, _08842_, _08841_);
  and _17133_ (_08844_, _08758_, word_in[30]);
  and _17134_ (_08845_, _08763_, _08457_);
  not _17135_ (_08847_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _17136_ (_08848_, _08763_, _08847_);
  nor _17137_ (_08849_, _08848_, _08845_);
  nor _17138_ (_08850_, _08849_, _08762_);
  and _17139_ (_08851_, _08762_, word_in[14]);
  or _17140_ (_08852_, _08851_, _08850_);
  or _17141_ (_08853_, _08852_, _08760_);
  or _17142_ (_08854_, _08769_, _08593_);
  and _17143_ (_08855_, _08854_, _08759_);
  and _17144_ (_08856_, _08855_, _08853_);
  or _17145_ (_07817_, _08856_, _08844_);
  and _17146_ (_08857_, _08758_, word_in[31]);
  and _17147_ (_08858_, _08763_, _08011_);
  nor _17148_ (_08859_, _08763_, _07716_);
  nor _17149_ (_08860_, _08859_, _08858_);
  nor _17150_ (_08861_, _08860_, _08762_);
  and _17151_ (_08862_, _08762_, word_in[15]);
  or _17152_ (_08863_, _08862_, _08861_);
  or _17153_ (_08864_, _08863_, _08760_);
  or _17154_ (_08865_, _08769_, _08023_);
  and _17155_ (_08866_, _08865_, _08759_);
  and _17156_ (_08867_, _08866_, _08864_);
  or _17157_ (_07822_, _08867_, _08857_);
  nand _17158_ (_08868_, _06890_, _06054_);
  and _17159_ (_08869_, _06061_, _05806_);
  and _17160_ (_08870_, _08869_, _06888_);
  not _17161_ (_08871_, _08870_);
  not _17162_ (_08872_, _06883_);
  and _17163_ (_08873_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _17164_ (_08874_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _17165_ (_08875_, _08874_, _08873_);
  or _17166_ (_08876_, _08875_, _06890_);
  and _17167_ (_08877_, _08876_, _08871_);
  and _17168_ (_08878_, _08877_, _08868_);
  and _17169_ (_08879_, _08870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _17170_ (_08880_, _08879_, _08878_);
  and _17171_ (_07864_, _08880_, _05110_);
  nand _17172_ (_08881_, _07337_, _06477_);
  or _17173_ (_08882_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _17174_ (_08883_, _08882_, _05110_);
  and _17175_ (_07867_, _08883_, _08881_);
  nor _17176_ (_08884_, _06890_, _08872_);
  or _17177_ (_08885_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  not _17178_ (_08886_, _08884_);
  or _17179_ (_08887_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _17180_ (_08888_, _08887_, _08885_);
  or _17181_ (_08889_, _08888_, _08870_);
  nand _17182_ (_08890_, _08870_, _06229_);
  and _17183_ (_08891_, _08890_, _05110_);
  and _17184_ (_07878_, _08891_, _08889_);
  nand _17185_ (_08892_, _08870_, _06054_);
  or _17186_ (_08893_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or _17187_ (_08894_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _17188_ (_08895_, _08894_, _08893_);
  or _17189_ (_08896_, _08895_, _08870_);
  and _17190_ (_08897_, _08896_, _05110_);
  and _17191_ (_07900_, _08897_, _08892_);
  and _17192_ (_08898_, _08021_, _07930_);
  and _17193_ (_08899_, _08898_, _07937_);
  and _17194_ (_08900_, _08899_, _07744_);
  not _17195_ (_08901_, _08900_);
  and _17196_ (_08902_, _07993_, _08037_);
  not _17197_ (_08903_, _08902_);
  and _17198_ (_08904_, _07999_, _08042_);
  not _17199_ (_08905_, _08904_);
  not _17200_ (_08907_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _17201_ (_08908_, _08007_, _07754_);
  and _17202_ (_08910_, _08908_, _08352_);
  nor _17203_ (_08911_, _08910_, _08907_);
  and _17204_ (_08912_, _08910_, word_in[0]);
  or _17205_ (_08914_, _08912_, _08911_);
  and _17206_ (_08915_, _08914_, _08905_);
  and _17207_ (_08917_, _08904_, word_in[8]);
  or _17208_ (_08918_, _08917_, _08915_);
  and _17209_ (_08919_, _08918_, _08903_);
  and _17210_ (_08921_, _08902_, word_in[16]);
  or _17211_ (_08922_, _08921_, _08919_);
  and _17212_ (_08924_, _08922_, _08901_);
  and _17213_ (_08925_, _08021_, word_in[24]);
  and _17214_ (_08927_, _08900_, _08925_);
  or _17215_ (_07911_, _08927_, _08924_);
  or _17216_ (_08928_, _08903_, word_in[17]);
  not _17217_ (_08929_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _17218_ (_08930_, _08910_, _08929_);
  and _17219_ (_08931_, _08910_, word_in[1]);
  or _17220_ (_08932_, _08931_, _08930_);
  or _17221_ (_08934_, _08932_, _08904_);
  or _17222_ (_08935_, _08905_, word_in[9]);
  and _17223_ (_08936_, _08935_, _08934_);
  or _17224_ (_08937_, _08936_, _08902_);
  and _17225_ (_08938_, _08937_, _08928_);
  or _17226_ (_08939_, _08938_, _08900_);
  or _17227_ (_08940_, _08901_, _08395_);
  and _17228_ (_07915_, _08940_, _08939_);
  not _17229_ (_08941_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _17230_ (_08942_, _08910_, _08941_);
  and _17231_ (_08943_, _08910_, word_in[2]);
  or _17232_ (_08944_, _08943_, _08942_);
  and _17233_ (_08945_, _08944_, _08905_);
  and _17234_ (_08946_, _08904_, word_in[10]);
  or _17235_ (_08947_, _08946_, _08945_);
  and _17236_ (_08948_, _08947_, _08903_);
  and _17237_ (_08949_, _08902_, word_in[18]);
  or _17238_ (_08950_, _08949_, _08900_);
  or _17239_ (_08951_, _08950_, _08948_);
  or _17240_ (_08952_, _08901_, _08411_);
  and _17241_ (_07919_, _08952_, _08951_);
  not _17242_ (_08953_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _17243_ (_08954_, _08910_, _08953_);
  and _17244_ (_08955_, _08910_, word_in[3]);
  or _17245_ (_08956_, _08955_, _08954_);
  and _17246_ (_08957_, _08956_, _08905_);
  and _17247_ (_08958_, _08904_, word_in[11]);
  or _17248_ (_08959_, _08958_, _08957_);
  and _17249_ (_08960_, _08959_, _08903_);
  and _17250_ (_08961_, _08902_, word_in[19]);
  or _17251_ (_08962_, _08961_, _08960_);
  and _17252_ (_08963_, _08962_, _08901_);
  and _17253_ (_08964_, _08900_, _08425_);
  or _17254_ (_07922_, _08964_, _08963_);
  not _17255_ (_08965_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _17256_ (_08966_, _08910_, _08965_);
  and _17257_ (_08967_, _08910_, word_in[4]);
  or _17258_ (_08968_, _08967_, _08966_);
  or _17259_ (_08969_, _08968_, _08904_);
  or _17260_ (_08970_, _08905_, word_in[12]);
  and _17261_ (_08971_, _08970_, _08969_);
  or _17262_ (_08972_, _08971_, _08902_);
  or _17263_ (_08973_, _08903_, word_in[20]);
  and _17264_ (_08974_, _08973_, _08972_);
  or _17265_ (_08975_, _08974_, _08900_);
  or _17266_ (_08976_, _08901_, _08439_);
  and _17267_ (_07924_, _08976_, _08975_);
  not _17268_ (_08977_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _17269_ (_08978_, _08910_, _08977_);
  and _17270_ (_08979_, _08910_, word_in[5]);
  or _17271_ (_08981_, _08979_, _08978_);
  or _17272_ (_08982_, _08981_, _08904_);
  or _17273_ (_08983_, _08905_, word_in[13]);
  and _17274_ (_08984_, _08983_, _08982_);
  or _17275_ (_08985_, _08984_, _08902_);
  nor _17276_ (_08986_, _08903_, word_in[21]);
  nor _17277_ (_08987_, _08986_, _08900_);
  and _17278_ (_08988_, _08987_, _08985_);
  and _17279_ (_08989_, _08900_, _08453_);
  or _17280_ (_07928_, _08989_, _08988_);
  not _17281_ (_08990_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _17282_ (_08991_, _08910_, _08990_);
  and _17283_ (_08992_, _08910_, word_in[6]);
  or _17284_ (_08993_, _08992_, _08991_);
  and _17285_ (_08994_, _08993_, _08905_);
  and _17286_ (_08995_, _08904_, word_in[14]);
  or _17287_ (_08996_, _08995_, _08994_);
  and _17288_ (_08997_, _08996_, _08903_);
  and _17289_ (_08998_, _08902_, word_in[22]);
  or _17290_ (_08999_, _08998_, _08900_);
  or _17291_ (_09000_, _08999_, _08997_);
  or _17292_ (_09001_, _08901_, _08469_);
  and _17293_ (_07932_, _09001_, _09000_);
  nor _17294_ (_09002_, _08910_, _07842_);
  and _17295_ (_09003_, _08910_, word_in[7]);
  or _17296_ (_09004_, _09003_, _09002_);
  and _17297_ (_09005_, _09004_, _08905_);
  and _17298_ (_09006_, _08904_, word_in[15]);
  or _17299_ (_09007_, _09006_, _09005_);
  and _17300_ (_09008_, _09007_, _08903_);
  and _17301_ (_09009_, _08902_, _08023_);
  or _17302_ (_09010_, _09009_, _08900_);
  or _17303_ (_09011_, _09010_, _09008_);
  or _17304_ (_09012_, _08901_, _08028_);
  and _17305_ (_07934_, _09012_, _09011_);
  and _17306_ (_09013_, _08899_, _07775_);
  not _17307_ (_09014_, _09013_);
  and _17308_ (_09015_, _07993_, _07858_);
  and _17309_ (_09016_, _09015_, _07907_);
  and _17310_ (_09017_, _09016_, _07746_);
  not _17311_ (_09018_, _09017_);
  or _17312_ (_09019_, _09018_, _08370_);
  and _17313_ (_09020_, _08493_, _07841_);
  not _17314_ (_09021_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _17315_ (_09022_, _08908_, _08496_);
  nor _17316_ (_09023_, _09022_, _09021_);
  and _17317_ (_09024_, _09022_, word_in[0]);
  or _17318_ (_09025_, _09024_, _09023_);
  or _17319_ (_09026_, _09025_, _09020_);
  not _17320_ (_09027_, _09020_);
  or _17321_ (_09028_, _09027_, word_in[8]);
  and _17322_ (_09029_, _09028_, _09026_);
  or _17323_ (_09030_, _09029_, _09017_);
  and _17324_ (_09031_, _09030_, _09019_);
  and _17325_ (_09032_, _09031_, _09014_);
  and _17326_ (_09033_, _09013_, word_in[24]);
  or _17327_ (_07991_, _09033_, _09032_);
  and _17328_ (_09034_, _09022_, word_in[1]);
  not _17329_ (_09035_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _17330_ (_09036_, _09022_, _09035_);
  nor _17331_ (_09037_, _09036_, _09034_);
  nor _17332_ (_09038_, _09037_, _09020_);
  and _17333_ (_09039_, _09020_, word_in[9]);
  or _17334_ (_09040_, _09039_, _09038_);
  and _17335_ (_09041_, _09040_, _09018_);
  and _17336_ (_09042_, _09017_, _08511_);
  or _17337_ (_09043_, _09042_, _09013_);
  or _17338_ (_09044_, _09043_, _09041_);
  or _17339_ (_09045_, _09014_, word_in[25]);
  and _17340_ (_07994_, _09045_, _09044_);
  and _17341_ (_09046_, _09017_, _08525_);
  and _17342_ (_09047_, _09022_, word_in[2]);
  not _17343_ (_09048_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _17344_ (_09049_, _09022_, _09048_);
  nor _17345_ (_09050_, _09049_, _09047_);
  nor _17346_ (_09051_, _09050_, _09020_);
  and _17347_ (_09052_, _09020_, word_in[10]);
  or _17348_ (_09053_, _09052_, _09051_);
  and _17349_ (_09054_, _09053_, _09018_);
  or _17350_ (_09055_, _09054_, _09046_);
  and _17351_ (_09056_, _09055_, _09014_);
  and _17352_ (_09057_, _09013_, word_in[26]);
  or _17353_ (_07997_, _09057_, _09056_);
  or _17354_ (_09058_, _09018_, _08546_);
  not _17355_ (_09059_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _17356_ (_09060_, _09022_, _09059_);
  and _17357_ (_09061_, _09022_, word_in[3]);
  or _17358_ (_09062_, _09061_, _09060_);
  or _17359_ (_09063_, _09062_, _09020_);
  or _17360_ (_09064_, _09027_, word_in[11]);
  and _17361_ (_09065_, _09064_, _09063_);
  or _17362_ (_09066_, _09065_, _09017_);
  and _17363_ (_09067_, _09066_, _09058_);
  or _17364_ (_09068_, _09067_, _09013_);
  or _17365_ (_09069_, _09014_, word_in[27]);
  and _17366_ (_08000_, _09069_, _09068_);
  and _17367_ (_09070_, _09022_, word_in[4]);
  not _17368_ (_09071_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _17369_ (_09072_, _09022_, _09071_);
  nor _17370_ (_09073_, _09072_, _09070_);
  nor _17371_ (_09074_, _09073_, _09020_);
  and _17372_ (_09075_, _09020_, word_in[12]);
  or _17373_ (_09076_, _09075_, _09074_);
  and _17374_ (_09077_, _09076_, _09018_);
  and _17375_ (_09078_, _09017_, _08564_);
  or _17376_ (_09079_, _09078_, _09013_);
  or _17377_ (_09080_, _09079_, _09077_);
  or _17378_ (_09081_, _09014_, word_in[28]);
  and _17379_ (_08003_, _09081_, _09080_);
  not _17380_ (_09082_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _17381_ (_09083_, _09022_, _09082_);
  and _17382_ (_09084_, _09022_, word_in[5]);
  nor _17383_ (_09085_, _09084_, _09083_);
  nor _17384_ (_09086_, _09085_, _09020_);
  and _17385_ (_09087_, _09020_, word_in[13]);
  or _17386_ (_09088_, _09087_, _09086_);
  and _17387_ (_09089_, _09088_, _09018_);
  and _17388_ (_09090_, _09017_, _08572_);
  or _17389_ (_09091_, _09090_, _09013_);
  or _17390_ (_09092_, _09091_, _09089_);
  or _17391_ (_09093_, _09014_, word_in[29]);
  and _17392_ (_08006_, _09093_, _09092_);
  and _17393_ (_09094_, _09022_, word_in[6]);
  not _17394_ (_09095_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _17395_ (_09096_, _09022_, _09095_);
  nor _17396_ (_09097_, _09096_, _09094_);
  nor _17397_ (_09098_, _09097_, _09020_);
  and _17398_ (_09099_, _09020_, word_in[14]);
  or _17399_ (_09100_, _09099_, _09098_);
  and _17400_ (_09101_, _09100_, _09018_);
  and _17401_ (_09102_, _09017_, _08593_);
  or _17402_ (_09103_, _09102_, _09013_);
  or _17403_ (_09104_, _09103_, _09101_);
  or _17404_ (_09105_, _09014_, word_in[30]);
  and _17405_ (_08009_, _09105_, _09104_);
  and _17406_ (_09106_, _09017_, _08023_);
  and _17407_ (_09107_, _09022_, word_in[7]);
  nor _17408_ (_09108_, _09022_, _07727_);
  nor _17409_ (_09109_, _09108_, _09107_);
  nor _17410_ (_09110_, _09109_, _09020_);
  and _17411_ (_09111_, _09020_, word_in[15]);
  or _17412_ (_09112_, _09111_, _09110_);
  and _17413_ (_09113_, _09112_, _09018_);
  or _17414_ (_09114_, _09113_, _09106_);
  and _17415_ (_09115_, _09114_, _09014_);
  and _17416_ (_09116_, _09013_, word_in[31]);
  or _17417_ (_08012_, _09116_, _09115_);
  and _17418_ (_09117_, _08630_, _07841_);
  not _17419_ (_09118_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _17420_ (_09119_, _08633_, _07754_);
  nor _17421_ (_09120_, _09119_, _09118_);
  and _17422_ (_09121_, _09119_, _08495_);
  or _17423_ (_09122_, _09121_, _09120_);
  or _17424_ (_09123_, _09122_, _09117_);
  and _17425_ (_09124_, _09016_, _07783_);
  not _17426_ (_09125_, _09124_);
  not _17427_ (_09126_, _09117_);
  or _17428_ (_09127_, _09126_, word_in[8]);
  and _17429_ (_09128_, _09127_, _09125_);
  and _17430_ (_09129_, _09128_, _09123_);
  and _17431_ (_09130_, _08899_, _07746_);
  and _17432_ (_09131_, _09124_, _08370_);
  or _17433_ (_09132_, _09131_, _09130_);
  or _17434_ (_09133_, _09132_, _09129_);
  not _17435_ (_09134_, _09130_);
  or _17436_ (_09135_, _09134_, word_in[24]);
  and _17437_ (_08077_, _09135_, _09133_);
  not _17438_ (_09136_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _17439_ (_09137_, _09119_, _09136_);
  and _17440_ (_09138_, _09119_, _08513_);
  nor _17441_ (_09139_, _09138_, _09137_);
  nor _17442_ (_09140_, _09139_, _09117_);
  and _17443_ (_09141_, _09117_, word_in[9]);
  or _17444_ (_09142_, _09141_, _09140_);
  and _17445_ (_09143_, _09142_, _09125_);
  and _17446_ (_09144_, _09124_, _08511_);
  or _17447_ (_09145_, _09144_, _09130_);
  or _17448_ (_09146_, _09145_, _09143_);
  or _17449_ (_09147_, _09134_, word_in[25]);
  and _17450_ (_08080_, _09147_, _09146_);
  not _17451_ (_09148_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _17452_ (_09149_, _09119_, _09148_);
  and _17453_ (_09150_, _09119_, _08401_);
  or _17454_ (_09151_, _09150_, _09149_);
  or _17455_ (_09152_, _09151_, _09117_);
  or _17456_ (_09153_, _09126_, word_in[10]);
  and _17457_ (_09154_, _09153_, _09125_);
  and _17458_ (_09155_, _09154_, _09152_);
  and _17459_ (_09156_, _09124_, _08525_);
  or _17460_ (_09157_, _09156_, _09130_);
  or _17461_ (_09158_, _09157_, _09155_);
  or _17462_ (_09159_, _09134_, word_in[26]);
  and _17463_ (_08084_, _09159_, _09158_);
  not _17464_ (_09160_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _17465_ (_09161_, _09119_, _09160_);
  and _17466_ (_09162_, _09119_, _08415_);
  or _17467_ (_09163_, _09162_, _09161_);
  or _17468_ (_09164_, _09163_, _09117_);
  or _17469_ (_09165_, _09126_, word_in[11]);
  and _17470_ (_09166_, _09165_, _09125_);
  and _17471_ (_09167_, _09166_, _09164_);
  and _17472_ (_09168_, _09124_, _08546_);
  or _17473_ (_09169_, _09168_, _09130_);
  or _17474_ (_09170_, _09169_, _09167_);
  or _17475_ (_09171_, _09134_, word_in[27]);
  and _17476_ (_08089_, _09171_, _09170_);
  not _17477_ (_09172_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _17478_ (_09173_, _09119_, _09172_);
  and _17479_ (_09174_, _09119_, _08429_);
  or _17480_ (_09175_, _09174_, _09173_);
  or _17481_ (_09176_, _09175_, _09117_);
  or _17482_ (_09177_, _09126_, word_in[12]);
  and _17483_ (_09178_, _09177_, _09125_);
  and _17484_ (_09179_, _09178_, _09176_);
  and _17485_ (_09180_, _09124_, _08564_);
  or _17486_ (_09181_, _09180_, _09130_);
  or _17487_ (_09182_, _09181_, _09179_);
  or _17488_ (_09183_, _09134_, word_in[28]);
  and _17489_ (_08091_, _09183_, _09182_);
  not _17490_ (_09184_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _17491_ (_09185_, _09119_, _09184_);
  and _17492_ (_09186_, _09119_, _08443_);
  or _17493_ (_09187_, _09186_, _09185_);
  or _17494_ (_09188_, _09187_, _09117_);
  or _17495_ (_09189_, _09126_, word_in[13]);
  and _17496_ (_09190_, _09189_, _09125_);
  and _17497_ (_09191_, _09190_, _09188_);
  and _17498_ (_09192_, _09124_, _08572_);
  or _17499_ (_09193_, _09192_, _09130_);
  or _17500_ (_09194_, _09193_, _09191_);
  or _17501_ (_09195_, _09134_, word_in[29]);
  and _17502_ (_08094_, _09195_, _09194_);
  or _17503_ (_09196_, _09125_, _08593_);
  not _17504_ (_09197_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _17505_ (_09198_, _09119_, _09197_);
  and _17506_ (_09199_, _09119_, _08457_);
  or _17507_ (_09200_, _09199_, _09198_);
  or _17508_ (_09201_, _09200_, _09117_);
  or _17509_ (_09202_, _09126_, word_in[14]);
  and _17510_ (_09203_, _09202_, _09201_);
  or _17511_ (_09204_, _09203_, _09124_);
  and _17512_ (_09205_, _09204_, _09196_);
  or _17513_ (_09206_, _09205_, _09130_);
  or _17514_ (_09207_, _09134_, word_in[30]);
  and _17515_ (_08098_, _09207_, _09206_);
  or _17516_ (_09208_, _09125_, _08023_);
  nor _17517_ (_09209_, _09119_, _07847_);
  and _17518_ (_09210_, _09119_, _08011_);
  or _17519_ (_09211_, _09210_, _09209_);
  or _17520_ (_09212_, _09211_, _09117_);
  or _17521_ (_09213_, _09126_, word_in[15]);
  and _17522_ (_09214_, _09213_, _09212_);
  or _17523_ (_09215_, _09214_, _09124_);
  and _17524_ (_09216_, _09215_, _09208_);
  or _17525_ (_09217_, _09216_, _09130_);
  or _17526_ (_09218_, _09134_, word_in[31]);
  and _17527_ (_08103_, _09218_, _09217_);
  and _17528_ (_09219_, _09016_, _07744_);
  not _17529_ (_09220_, _09219_);
  and _17530_ (_09221_, _08001_, _07841_);
  not _17531_ (_09222_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _17532_ (_09223_, _08908_, _08005_);
  nor _17533_ (_09224_, _09223_, _09222_);
  and _17534_ (_09225_, _09223_, word_in[0]);
  nor _17535_ (_09226_, _09225_, _09224_);
  nor _17536_ (_09227_, _09226_, _09221_);
  and _17537_ (_09228_, _09221_, word_in[8]);
  or _17538_ (_09229_, _09228_, _09227_);
  and _17539_ (_09230_, _09229_, _09220_);
  and _17540_ (_09232_, _08021_, _08059_);
  and _17541_ (_09233_, _09219_, _08370_);
  or _17542_ (_09235_, _09233_, _09232_);
  or _17543_ (_09236_, _09235_, _09230_);
  not _17544_ (_09237_, _09232_);
  or _17545_ (_09238_, _09237_, _08925_);
  and _17546_ (_08171_, _09238_, _09236_);
  not _17547_ (_09239_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _17548_ (_09240_, _09223_, _09239_);
  and _17549_ (_09241_, _09223_, word_in[1]);
  nor _17550_ (_09242_, _09241_, _09240_);
  nor _17551_ (_09244_, _09242_, _09221_);
  and _17552_ (_09245_, _09221_, word_in[9]);
  or _17553_ (_09246_, _09245_, _09244_);
  and _17554_ (_09247_, _09246_, _09220_);
  and _17555_ (_09248_, _09219_, _08511_);
  or _17556_ (_09249_, _09248_, _09232_);
  or _17557_ (_09250_, _09249_, _09247_);
  or _17558_ (_09251_, _09237_, _08395_);
  and _17559_ (_08175_, _09251_, _09250_);
  not _17560_ (_09252_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _17561_ (_09253_, _09223_, _09252_);
  and _17562_ (_09254_, _09223_, word_in[2]);
  nor _17563_ (_09255_, _09254_, _09253_);
  nor _17564_ (_09256_, _09255_, _09221_);
  and _17565_ (_09257_, _09221_, word_in[10]);
  or _17566_ (_09258_, _09257_, _09256_);
  and _17567_ (_09259_, _09258_, _09220_);
  and _17568_ (_09260_, _09219_, _08525_);
  or _17569_ (_09261_, _09260_, _09232_);
  or _17570_ (_09262_, _09261_, _09259_);
  or _17571_ (_09263_, _09237_, _08411_);
  and _17572_ (_13444_, _09263_, _09262_);
  not _17573_ (_09264_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _17574_ (_09265_, _09223_, _09264_);
  and _17575_ (_09266_, _09223_, word_in[3]);
  nor _17576_ (_09267_, _09266_, _09265_);
  nor _17577_ (_09268_, _09267_, _09221_);
  and _17578_ (_09269_, _09221_, word_in[11]);
  or _17579_ (_09270_, _09269_, _09268_);
  and _17580_ (_09271_, _09270_, _09220_);
  and _17581_ (_09272_, _09219_, _08546_);
  or _17582_ (_09273_, _09272_, _09232_);
  or _17583_ (_09274_, _09273_, _09271_);
  or _17584_ (_09275_, _09237_, _08425_);
  and _17585_ (_13445_, _09275_, _09274_);
  not _17586_ (_09276_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _17587_ (_09277_, _09223_, _09276_);
  and _17588_ (_09278_, _09223_, word_in[4]);
  nor _17589_ (_09279_, _09278_, _09277_);
  nor _17590_ (_09280_, _09279_, _09221_);
  and _17591_ (_09281_, _09221_, word_in[12]);
  or _17592_ (_09282_, _09281_, _09280_);
  and _17593_ (_09283_, _09282_, _09220_);
  and _17594_ (_09284_, _09219_, _08564_);
  or _17595_ (_09285_, _09284_, _09232_);
  or _17596_ (_09286_, _09285_, _09283_);
  or _17597_ (_09287_, _09237_, _08439_);
  and _17598_ (_13446_, _09287_, _09286_);
  not _17599_ (_09288_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _17600_ (_09289_, _09223_, _09288_);
  and _17601_ (_09290_, _09223_, word_in[5]);
  nor _17602_ (_09291_, _09290_, _09289_);
  nor _17603_ (_09292_, _09291_, _09221_);
  and _17604_ (_09293_, _09221_, word_in[13]);
  or _17605_ (_09294_, _09293_, _09292_);
  and _17606_ (_09295_, _09294_, _09220_);
  and _17607_ (_09296_, _09219_, _08572_);
  or _17608_ (_09297_, _09296_, _09232_);
  or _17609_ (_09298_, _09297_, _09295_);
  or _17610_ (_09299_, _09237_, _08453_);
  and _17611_ (_13447_, _09299_, _09298_);
  not _17612_ (_09300_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _17613_ (_09301_, _09223_, _09300_);
  and _17614_ (_09302_, _09223_, word_in[6]);
  nor _17615_ (_09303_, _09302_, _09301_);
  nor _17616_ (_09304_, _09303_, _09221_);
  and _17617_ (_09305_, _09221_, word_in[14]);
  or _17618_ (_09306_, _09305_, _09304_);
  and _17619_ (_09307_, _09306_, _09220_);
  and _17620_ (_09308_, _09219_, _08593_);
  or _17621_ (_09309_, _09308_, _09232_);
  or _17622_ (_09310_, _09309_, _09307_);
  or _17623_ (_09311_, _09237_, _08469_);
  and _17624_ (_13448_, _09311_, _09310_);
  nor _17625_ (_09312_, _09223_, _07721_);
  and _17626_ (_09313_, _09223_, word_in[7]);
  nor _17627_ (_09314_, _09313_, _09312_);
  nor _17628_ (_09315_, _09314_, _09221_);
  and _17629_ (_09316_, _09221_, word_in[15]);
  or _17630_ (_09317_, _09316_, _09315_);
  and _17631_ (_09318_, _09317_, _09220_);
  and _17632_ (_09319_, _09219_, _08023_);
  or _17633_ (_09320_, _09319_, _09232_);
  or _17634_ (_09321_, _09320_, _09318_);
  or _17635_ (_09322_, _09237_, _08028_);
  and _17636_ (_08185_, _09322_, _09321_);
  nor _17637_ (_09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and _17638_ (_09324_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _17639_ (_09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _05110_);
  and _17640_ (_09326_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or _17641_ (_08247_, _09326_, _09324_);
  nor _17642_ (_09327_, _08342_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and _17643_ (_09328_, _08342_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _17644_ (_09329_, _09328_, _09327_);
  nand _17645_ (_09330_, _09329_, _05110_);
  nor _17646_ (_08250_, _09330_, _08274_);
  and _17647_ (_09331_, _07993_, _08096_);
  not _17648_ (_09332_, _09331_);
  and _17649_ (_09333_, _07999_, _07755_);
  not _17650_ (_09334_, _09333_);
  not _17651_ (_09335_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _17652_ (_09336_, _08354_, _07753_);
  and _17653_ (_09337_, _09336_, _08352_);
  nor _17654_ (_09338_, _09337_, _09335_);
  and _17655_ (_09339_, _09337_, _08495_);
  or _17656_ (_09340_, _09339_, _09338_);
  and _17657_ (_09341_, _09340_, _09334_);
  and _17658_ (_09342_, _09333_, word_in[8]);
  or _17659_ (_09343_, _09342_, _09341_);
  and _17660_ (_09344_, _09343_, _09332_);
  and _17661_ (_09345_, _08021_, _08074_);
  and _17662_ (_09346_, _09331_, word_in[16]);
  or _17663_ (_09347_, _09346_, _09345_);
  or _17664_ (_09348_, _09347_, _09344_);
  not _17665_ (_09349_, _09345_);
  or _17666_ (_09350_, _09349_, _08925_);
  and _17667_ (_13449_, _09350_, _09348_);
  not _17668_ (_09351_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _17669_ (_09352_, _09337_, _09351_);
  and _17670_ (_09353_, _09337_, _08513_);
  or _17671_ (_09354_, _09353_, _09352_);
  and _17672_ (_09355_, _09354_, _09334_);
  and _17673_ (_09356_, _09333_, word_in[9]);
  or _17674_ (_09357_, _09356_, _09355_);
  and _17675_ (_09358_, _09357_, _09332_);
  and _17676_ (_09359_, _09331_, word_in[17]);
  or _17677_ (_09360_, _09359_, _09358_);
  and _17678_ (_09361_, _09360_, _09349_);
  and _17679_ (_09362_, _09345_, word_in[25]);
  or _17680_ (_08271_, _09362_, _09361_);
  not _17681_ (_09363_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _17682_ (_09364_, _09337_, _09363_);
  and _17683_ (_09365_, _09337_, _08401_);
  or _17684_ (_09366_, _09365_, _09364_);
  and _17685_ (_09367_, _09366_, _09334_);
  and _17686_ (_09368_, _09333_, word_in[10]);
  or _17687_ (_09369_, _09368_, _09367_);
  and _17688_ (_09370_, _09369_, _09332_);
  and _17689_ (_09371_, _09331_, word_in[18]);
  or _17690_ (_09372_, _09371_, _09370_);
  and _17691_ (_09373_, _09372_, _09349_);
  and _17692_ (_09374_, _09345_, word_in[26]);
  or _17693_ (_08275_, _09374_, _09373_);
  not _17694_ (_09375_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _17695_ (_09376_, _09337_, _09375_);
  and _17696_ (_09377_, _09337_, _08415_);
  or _17697_ (_09378_, _09377_, _09376_);
  and _17698_ (_09379_, _09378_, _09334_);
  and _17699_ (_09380_, _09333_, word_in[11]);
  or _17700_ (_09381_, _09380_, _09379_);
  and _17701_ (_09382_, _09381_, _09332_);
  and _17702_ (_09383_, _09331_, word_in[19]);
  or _17703_ (_09384_, _09383_, _09345_);
  or _17704_ (_09385_, _09384_, _09382_);
  or _17705_ (_09386_, _09349_, _08425_);
  and _17706_ (_08279_, _09386_, _09385_);
  not _17707_ (_09387_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _17708_ (_09388_, _09337_, _09387_);
  and _17709_ (_09389_, _09337_, _08429_);
  or _17710_ (_09390_, _09389_, _09388_);
  and _17711_ (_09391_, _09390_, _09334_);
  and _17712_ (_09392_, _09333_, word_in[12]);
  or _17713_ (_09393_, _09392_, _09391_);
  and _17714_ (_09394_, _09393_, _09332_);
  and _17715_ (_09395_, _09331_, word_in[20]);
  or _17716_ (_09396_, _09395_, _09345_);
  or _17717_ (_09397_, _09396_, _09394_);
  or _17718_ (_09398_, _09349_, _08439_);
  and _17719_ (_08284_, _09398_, _09397_);
  not _17720_ (_09399_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _17721_ (_09400_, _09337_, _09399_);
  and _17722_ (_09401_, _09337_, _08443_);
  or _17723_ (_09402_, _09401_, _09400_);
  and _17724_ (_09403_, _09402_, _09334_);
  and _17725_ (_09404_, _09333_, word_in[13]);
  or _17726_ (_09405_, _09404_, _09403_);
  and _17727_ (_09406_, _09405_, _09332_);
  and _17728_ (_09407_, _09331_, word_in[21]);
  or _17729_ (_09408_, _09407_, _09406_);
  and _17730_ (_09409_, _09408_, _09349_);
  and _17731_ (_09410_, _09345_, word_in[29]);
  or _17732_ (_08289_, _09410_, _09409_);
  not _17733_ (_09411_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _17734_ (_09412_, _09337_, _09411_);
  and _17735_ (_09413_, _09337_, _08457_);
  or _17736_ (_09414_, _09413_, _09412_);
  and _17737_ (_09415_, _09414_, _09334_);
  and _17738_ (_09416_, _09333_, word_in[14]);
  or _17739_ (_09417_, _09416_, _09415_);
  and _17740_ (_09418_, _09417_, _09332_);
  and _17741_ (_09419_, _09331_, word_in[22]);
  or _17742_ (_09420_, _09419_, _09418_);
  and _17743_ (_09421_, _09420_, _09349_);
  and _17744_ (_09422_, _09345_, word_in[30]);
  or _17745_ (_08295_, _09422_, _09421_);
  and _17746_ (_09423_, _09331_, word_in[23]);
  nor _17747_ (_09424_, _09337_, _07804_);
  and _17748_ (_09425_, _09337_, _08011_);
  or _17749_ (_09426_, _09425_, _09424_);
  and _17750_ (_09427_, _09426_, _09334_);
  and _17751_ (_09428_, _09333_, word_in[15]);
  or _17752_ (_09429_, _09428_, _09427_);
  and _17753_ (_09430_, _09429_, _09332_);
  or _17754_ (_09431_, _09430_, _09423_);
  and _17755_ (_09432_, _09431_, _09349_);
  and _17756_ (_09433_, _09345_, word_in[31]);
  or _17757_ (_08299_, _09433_, _09432_);
  and _17758_ (_09434_, _08490_, _07865_);
  and _17759_ (_09435_, _08493_, _07757_);
  not _17760_ (_09436_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _17761_ (_09437_, _09336_, _08496_);
  nor _17762_ (_09438_, _09437_, _09436_);
  and _17763_ (_09439_, _09437_, _08495_);
  or _17764_ (_09440_, _09439_, _09438_);
  or _17765_ (_09441_, _09440_, _09435_);
  not _17766_ (_09442_, _09435_);
  or _17767_ (_09443_, _09442_, word_in[8]);
  and _17768_ (_09444_, _09443_, _09441_);
  or _17769_ (_09445_, _09444_, _09434_);
  and _17770_ (_09446_, _08021_, _07938_);
  and _17771_ (_09447_, _09446_, _07775_);
  not _17772_ (_09448_, _09434_);
  nor _17773_ (_09449_, _09448_, _08370_);
  nor _17774_ (_09450_, _09449_, _09447_);
  and _17775_ (_09451_, _09450_, _09445_);
  and _17776_ (_09452_, _09447_, _08925_);
  or _17777_ (_08374_, _09452_, _09451_);
  not _17778_ (_09453_, _09447_);
  and _17779_ (_09454_, _09434_, _08511_);
  and _17780_ (_09455_, _09437_, _08513_);
  not _17781_ (_09456_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _17782_ (_09457_, _09437_, _09456_);
  or _17783_ (_09458_, _09457_, _09455_);
  or _17784_ (_09459_, _09458_, _09435_);
  or _17785_ (_09460_, _09442_, word_in[9]);
  and _17786_ (_09461_, _09460_, _09448_);
  and _17787_ (_09462_, _09461_, _09459_);
  or _17788_ (_09463_, _09462_, _09454_);
  and _17789_ (_09464_, _09463_, _09453_);
  and _17790_ (_09465_, _09447_, word_in[25]);
  or _17791_ (_08377_, _09465_, _09464_);
  or _17792_ (_09466_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not _17793_ (_09467_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand _17794_ (_09468_, _06205_, _09467_);
  and _17795_ (_09469_, _09468_, _05110_);
  and _17796_ (_08380_, _09469_, _09466_);
  and _17797_ (_09470_, _09437_, _08401_);
  not _17798_ (_09471_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _17799_ (_09472_, _09437_, _09471_);
  or _17800_ (_09473_, _09472_, _09470_);
  or _17801_ (_09474_, _09473_, _09435_);
  or _17802_ (_09475_, _09442_, word_in[10]);
  and _17803_ (_09476_, _09475_, _09448_);
  and _17804_ (_09477_, _09476_, _09474_);
  and _17805_ (_09478_, _09434_, _08525_);
  or _17806_ (_09479_, _09478_, _09447_);
  or _17807_ (_09480_, _09479_, _09477_);
  or _17808_ (_09481_, _09453_, _08411_);
  and _17809_ (_08382_, _09481_, _09480_);
  not _17810_ (_09482_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _17811_ (_09483_, _09437_, _09482_);
  and _17812_ (_09484_, _09437_, _08415_);
  or _17813_ (_09485_, _09484_, _09483_);
  or _17814_ (_09486_, _09485_, _09435_);
  or _17815_ (_09487_, _09442_, word_in[11]);
  and _17816_ (_09488_, _09487_, _09486_);
  or _17817_ (_09489_, _09488_, _09434_);
  nor _17818_ (_09490_, _09448_, _08546_);
  nor _17819_ (_09491_, _09490_, _09447_);
  and _17820_ (_09492_, _09491_, _09489_);
  and _17821_ (_09493_, _09447_, _08425_);
  or _17822_ (_08386_, _09493_, _09492_);
  not _17823_ (_09494_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _17824_ (_09495_, _09437_, _09494_);
  and _17825_ (_09496_, _09437_, _08429_);
  or _17826_ (_09497_, _09496_, _09495_);
  or _17827_ (_09498_, _09497_, _09435_);
  or _17828_ (_09499_, _09442_, word_in[12]);
  and _17829_ (_09500_, _09499_, _09498_);
  or _17830_ (_09501_, _09500_, _09434_);
  nor _17831_ (_09502_, _09448_, _08564_);
  nor _17832_ (_09503_, _09502_, _09447_);
  and _17833_ (_09504_, _09503_, _09501_);
  and _17834_ (_09505_, _09447_, _08439_);
  or _17835_ (_08389_, _09505_, _09504_);
  not _17836_ (_09506_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _17837_ (_09507_, _09437_, _09506_);
  and _17838_ (_09508_, _09437_, _08443_);
  or _17839_ (_09509_, _09508_, _09507_);
  or _17840_ (_09510_, _09509_, _09435_);
  or _17841_ (_09511_, _09442_, word_in[13]);
  and _17842_ (_09512_, _09511_, _09510_);
  or _17843_ (_09513_, _09512_, _09434_);
  nor _17844_ (_09514_, _09448_, _08572_);
  nor _17845_ (_09515_, _09514_, _09447_);
  and _17846_ (_09516_, _09515_, _09513_);
  and _17847_ (_09517_, _09447_, _08453_);
  or _17848_ (_08392_, _09517_, _09516_);
  not _17849_ (_09518_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _17850_ (_09519_, _09437_, _09518_);
  and _17851_ (_09520_, _09437_, _08457_);
  or _17852_ (_09521_, _09520_, _09519_);
  or _17853_ (_09522_, _09521_, _09435_);
  or _17854_ (_09523_, _09442_, word_in[14]);
  and _17855_ (_09524_, _09523_, _09522_);
  or _17856_ (_09525_, _09524_, _09434_);
  nor _17857_ (_09526_, _09448_, _08593_);
  nor _17858_ (_09527_, _09526_, _09447_);
  and _17859_ (_09528_, _09527_, _09525_);
  and _17860_ (_09529_, _09447_, _08469_);
  or _17861_ (_08396_, _09529_, _09528_);
  nor _17862_ (_09530_, _09437_, _07706_);
  and _17863_ (_09531_, _09437_, _08011_);
  or _17864_ (_09532_, _09531_, _09530_);
  or _17865_ (_09533_, _09532_, _09435_);
  or _17866_ (_09534_, _09442_, word_in[15]);
  and _17867_ (_09535_, _09534_, _09533_);
  or _17868_ (_09536_, _09535_, _09434_);
  nor _17869_ (_09537_, _09448_, _08023_);
  nor _17870_ (_09538_, _09537_, _09447_);
  and _17871_ (_09539_, _09538_, _09536_);
  and _17872_ (_09540_, _09447_, _08028_);
  or _17873_ (_08399_, _09540_, _09539_);
  and _17874_ (_09541_, _08642_, _07865_);
  and _17875_ (_09542_, _08630_, _07757_);
  not _17876_ (_09543_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _17877_ (_09544_, _09336_, _08633_);
  nor _17878_ (_09545_, _09544_, _09543_);
  and _17879_ (_09546_, _09544_, _08495_);
  or _17880_ (_09547_, _09546_, _09545_);
  or _17881_ (_09548_, _09547_, _09542_);
  not _17882_ (_09549_, _09542_);
  or _17883_ (_09550_, _09549_, word_in[8]);
  and _17884_ (_09551_, _09550_, _09548_);
  or _17885_ (_09552_, _09551_, _09541_);
  and _17886_ (_09553_, _09446_, _07746_);
  not _17887_ (_09554_, _09541_);
  nor _17888_ (_09555_, _09554_, _08370_);
  nor _17889_ (_09556_, _09555_, _09553_);
  and _17890_ (_09557_, _09556_, _09552_);
  and _17891_ (_09558_, _09553_, _08925_);
  or _17892_ (_08465_, _09558_, _09557_);
  not _17893_ (_09559_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _17894_ (_09560_, _09544_, _09559_);
  and _17895_ (_09561_, _09544_, _08513_);
  or _17896_ (_09562_, _09561_, _09560_);
  or _17897_ (_09563_, _09562_, _09542_);
  or _17898_ (_09564_, _09549_, word_in[9]);
  and _17899_ (_09565_, _09564_, _09563_);
  or _17900_ (_09566_, _09565_, _09541_);
  nor _17901_ (_09567_, _09554_, _08511_);
  nor _17902_ (_09568_, _09567_, _09553_);
  and _17903_ (_09569_, _09568_, _09566_);
  and _17904_ (_09570_, _09553_, _08395_);
  or _17905_ (_08468_, _09570_, _09569_);
  and _17906_ (_09571_, _09544_, _08401_);
  not _17907_ (_09572_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _17908_ (_09573_, _09544_, _09572_);
  or _17909_ (_09574_, _09573_, _09571_);
  or _17910_ (_09575_, _09574_, _09542_);
  or _17911_ (_09576_, _09549_, word_in[10]);
  and _17912_ (_09577_, _09576_, _09554_);
  and _17913_ (_09578_, _09577_, _09575_);
  and _17914_ (_09579_, _09541_, _08525_);
  or _17915_ (_09580_, _09579_, _09553_);
  or _17916_ (_09581_, _09580_, _09578_);
  not _17917_ (_09582_, _09553_);
  or _17918_ (_09583_, _09582_, _08411_);
  and _17919_ (_08472_, _09583_, _09581_);
  and _17920_ (_09584_, _09544_, _08415_);
  not _17921_ (_09585_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _17922_ (_09586_, _09544_, _09585_);
  or _17923_ (_09587_, _09586_, _09584_);
  or _17924_ (_09588_, _09587_, _09542_);
  or _17925_ (_09589_, _09549_, word_in[11]);
  and _17926_ (_09590_, _09589_, _09554_);
  and _17927_ (_09591_, _09590_, _09588_);
  and _17928_ (_09592_, _09541_, _08546_);
  or _17929_ (_09593_, _09592_, _09553_);
  or _17930_ (_09594_, _09593_, _09591_);
  or _17931_ (_09595_, _09582_, _08425_);
  and _17932_ (_08475_, _09595_, _09594_);
  and _17933_ (_09596_, _09541_, _08564_);
  and _17934_ (_09597_, _09544_, _08429_);
  not _17935_ (_09598_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _17936_ (_09599_, _09544_, _09598_);
  or _17937_ (_09600_, _09599_, _09597_);
  or _17938_ (_09601_, _09600_, _09542_);
  or _17939_ (_09602_, _09549_, word_in[12]);
  and _17940_ (_09603_, _09602_, _09554_);
  and _17941_ (_09604_, _09603_, _09601_);
  or _17942_ (_09605_, _09604_, _09596_);
  and _17943_ (_09606_, _09605_, _09582_);
  and _17944_ (_09607_, _09553_, word_in[28]);
  or _17945_ (_08477_, _09607_, _09606_);
  not _17946_ (_09608_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _17947_ (_09609_, _09544_, _09608_);
  and _17948_ (_09610_, _09544_, _08443_);
  or _17949_ (_09611_, _09610_, _09609_);
  or _17950_ (_09612_, _09611_, _09542_);
  or _17951_ (_09613_, _09549_, word_in[13]);
  and _17952_ (_09614_, _09613_, _09612_);
  or _17953_ (_09615_, _09614_, _09541_);
  nor _17954_ (_09616_, _09554_, _08572_);
  nor _17955_ (_09617_, _09616_, _09553_);
  and _17956_ (_09618_, _09617_, _09615_);
  and _17957_ (_09619_, _09553_, _08453_);
  or _17958_ (_08479_, _09619_, _09618_);
  and _17959_ (_09620_, _09544_, _08457_);
  not _17960_ (_09621_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _17961_ (_09622_, _09544_, _09621_);
  or _17962_ (_09623_, _09622_, _09620_);
  or _17963_ (_09624_, _09623_, _09542_);
  or _17964_ (_09625_, _09549_, word_in[14]);
  and _17965_ (_09626_, _09625_, _09554_);
  and _17966_ (_09627_, _09626_, _09624_);
  and _17967_ (_09628_, _09541_, _08593_);
  or _17968_ (_09630_, _09628_, _09553_);
  or _17969_ (_09631_, _09630_, _09627_);
  or _17970_ (_09632_, _09582_, _08469_);
  and _17971_ (_08482_, _09632_, _09631_);
  and _17972_ (_09634_, _09541_, _08023_);
  and _17973_ (_09635_, _09544_, _08011_);
  nor _17974_ (_09637_, _09544_, _07797_);
  nor _17975_ (_09638_, _09637_, _09635_);
  nor _17976_ (_09640_, _09638_, _09542_);
  and _17977_ (_09641_, _09542_, word_in[15]);
  or _17978_ (_09642_, _09641_, _09640_);
  and _17979_ (_09643_, _09642_, _09554_);
  or _17980_ (_09644_, _09643_, _09634_);
  and _17981_ (_09645_, _09644_, _09582_);
  and _17982_ (_09646_, _09553_, word_in[31]);
  or _17983_ (_08485_, _09646_, _09645_);
  and _17984_ (_09647_, _07995_, _07865_);
  and _17985_ (_09648_, _08001_, _07757_);
  not _17986_ (_09649_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _17987_ (_09650_, _09336_, _08005_);
  nor _17988_ (_09651_, _09650_, _09649_);
  and _17989_ (_09652_, _09650_, _08495_);
  or _17990_ (_09653_, _09652_, _09651_);
  or _17991_ (_09654_, _09653_, _09648_);
  not _17992_ (_09655_, _09648_);
  or _17993_ (_09656_, _09655_, word_in[8]);
  and _17994_ (_09657_, _09656_, _09654_);
  or _17995_ (_09658_, _09657_, _09647_);
  and _17996_ (_09659_, _08021_, _08156_);
  not _17997_ (_09660_, _09659_);
  not _17998_ (_09661_, _09647_);
  or _17999_ (_09662_, _09661_, _08370_);
  and _18000_ (_09663_, _09662_, _09660_);
  and _18001_ (_09664_, _09663_, _09658_);
  and _18002_ (_09665_, _09659_, word_in[24]);
  or _18003_ (_08550_, _09665_, _09664_);
  and _18004_ (_09666_, _09659_, word_in[25]);
  not _18005_ (_09667_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _18006_ (_09668_, _09650_, _09667_);
  and _18007_ (_09669_, _09650_, _08513_);
  or _18008_ (_09670_, _09669_, _09668_);
  or _18009_ (_09671_, _09670_, _09648_);
  or _18010_ (_09672_, _09655_, word_in[9]);
  and _18011_ (_09673_, _09672_, _09671_);
  or _18012_ (_09674_, _09673_, _09647_);
  or _18013_ (_09675_, _09661_, _08511_);
  and _18014_ (_09676_, _09675_, _09660_);
  and _18015_ (_09677_, _09676_, _09674_);
  or _18016_ (_08552_, _09677_, _09666_);
  and _18017_ (_09678_, _09647_, _08525_);
  and _18018_ (_09679_, _09650_, _08401_);
  not _18019_ (_09680_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _18020_ (_09681_, _09650_, _09680_);
  or _18021_ (_09682_, _09681_, _09679_);
  or _18022_ (_09683_, _09682_, _09648_);
  or _18023_ (_09684_, _09655_, word_in[10]);
  and _18024_ (_09685_, _09684_, _09661_);
  and _18025_ (_09686_, _09685_, _09683_);
  or _18026_ (_09687_, _09686_, _09678_);
  and _18027_ (_09688_, _09687_, _09660_);
  and _18028_ (_09689_, _09659_, word_in[26]);
  or _18029_ (_08556_, _09689_, _09688_);
  and _18030_ (_09690_, _09647_, _08546_);
  and _18031_ (_09691_, _09650_, _08415_);
  not _18032_ (_09692_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _18033_ (_09693_, _09650_, _09692_);
  or _18034_ (_09694_, _09693_, _09691_);
  or _18035_ (_09695_, _09694_, _09648_);
  or _18036_ (_09696_, _09655_, word_in[11]);
  and _18037_ (_09697_, _09696_, _09661_);
  and _18038_ (_09698_, _09697_, _09695_);
  or _18039_ (_09699_, _09698_, _09690_);
  and _18040_ (_09700_, _09699_, _09660_);
  and _18041_ (_09701_, _09659_, word_in[27]);
  or _18042_ (_08559_, _09701_, _09700_);
  and _18043_ (_09702_, _09659_, word_in[28]);
  not _18044_ (_09703_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _18045_ (_09704_, _09650_, _09703_);
  and _18046_ (_09705_, _09650_, _08429_);
  or _18047_ (_09706_, _09705_, _09704_);
  or _18048_ (_09707_, _09706_, _09648_);
  or _18049_ (_09708_, _09655_, word_in[12]);
  and _18050_ (_09709_, _09708_, _09707_);
  or _18051_ (_09710_, _09709_, _09647_);
  or _18052_ (_09711_, _09661_, _08564_);
  and _18053_ (_09712_, _09711_, _09660_);
  and _18054_ (_09713_, _09712_, _09710_);
  or _18055_ (_08562_, _09713_, _09702_);
  and _18056_ (_09714_, _09647_, _08572_);
  and _18057_ (_09715_, _09650_, _08443_);
  not _18058_ (_09716_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _18059_ (_09717_, _09650_, _09716_);
  or _18060_ (_09718_, _09717_, _09715_);
  or _18061_ (_09719_, _09718_, _09648_);
  or _18062_ (_09720_, _09655_, word_in[13]);
  and _18063_ (_09721_, _09720_, _09661_);
  and _18064_ (_09722_, _09721_, _09719_);
  or _18065_ (_09723_, _09722_, _09714_);
  and _18066_ (_09724_, _09723_, _09660_);
  and _18067_ (_09725_, _09659_, word_in[29]);
  or _18068_ (_08566_, _09725_, _09724_);
  and _18069_ (_09726_, _09647_, _08593_);
  and _18070_ (_09727_, _09650_, _08457_);
  not _18071_ (_09728_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _18072_ (_09729_, _09650_, _09728_);
  or _18073_ (_09730_, _09729_, _09727_);
  or _18074_ (_09731_, _09730_, _09648_);
  or _18075_ (_09732_, _09655_, word_in[14]);
  and _18076_ (_09733_, _09732_, _09661_);
  and _18077_ (_09734_, _09733_, _09731_);
  or _18078_ (_09735_, _09734_, _09726_);
  and _18079_ (_09736_, _09735_, _09660_);
  and _18080_ (_09738_, _09659_, word_in[30]);
  or _18081_ (_08568_, _09738_, _09736_);
  and _18082_ (_09739_, _09659_, word_in[31]);
  nor _18083_ (_09740_, _09650_, _07691_);
  and _18084_ (_09741_, _09650_, _08011_);
  or _18085_ (_09742_, _09741_, _09740_);
  or _18086_ (_09743_, _09742_, _09648_);
  or _18087_ (_09744_, _09655_, word_in[15]);
  and _18088_ (_09745_, _09744_, _09743_);
  or _18089_ (_09746_, _09745_, _09647_);
  or _18090_ (_09747_, _09661_, _08023_);
  and _18091_ (_09748_, _09747_, _09660_);
  and _18092_ (_09749_, _09748_, _09746_);
  or _18093_ (_08571_, _09749_, _09739_);
  and _18094_ (_09750_, _07993_, _08190_);
  not _18095_ (_09751_, _09750_);
  and _18096_ (_09752_, _07999_, _08211_);
  not _18097_ (_09753_, _09752_);
  not _18098_ (_09754_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _18099_ (_09755_, _08352_, _08008_);
  nor _18100_ (_09756_, _09755_, _09754_);
  and _18101_ (_09757_, _09755_, word_in[0]);
  or _18102_ (_09758_, _09757_, _09756_);
  and _18103_ (_09759_, _09758_, _09753_);
  and _18104_ (_09760_, _09752_, word_in[8]);
  or _18105_ (_09761_, _09760_, _09759_);
  and _18106_ (_09762_, _09761_, _09751_);
  not _18107_ (_09763_, _07937_);
  and _18108_ (_09764_, _08898_, _09763_);
  and _18109_ (_09765_, _09764_, _07744_);
  and _18110_ (_09766_, _09750_, word_in[16]);
  or _18111_ (_09767_, _09766_, _09765_);
  or _18112_ (_09768_, _09767_, _09762_);
  not _18113_ (_09769_, _09765_);
  or _18114_ (_09770_, _09769_, _08925_);
  and _18115_ (_08636_, _09770_, _09768_);
  not _18116_ (_09771_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _18117_ (_09772_, _09755_, _09771_);
  and _18118_ (_09773_, _09755_, word_in[1]);
  or _18119_ (_09774_, _09773_, _09772_);
  and _18120_ (_09775_, _09774_, _09753_);
  and _18121_ (_09776_, _09752_, word_in[9]);
  or _18122_ (_09777_, _09776_, _09775_);
  and _18123_ (_09778_, _09777_, _09751_);
  and _18124_ (_09779_, _09750_, word_in[17]);
  or _18125_ (_09780_, _09779_, _09765_);
  or _18126_ (_09781_, _09780_, _09778_);
  or _18127_ (_09782_, _09769_, _08395_);
  and _18128_ (_08640_, _09782_, _09781_);
  not _18129_ (_09783_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _18130_ (_09784_, _09755_, _09783_);
  and _18131_ (_09785_, _09755_, word_in[2]);
  or _18132_ (_09786_, _09785_, _09784_);
  and _18133_ (_09787_, _09786_, _09753_);
  and _18134_ (_09788_, _09752_, word_in[10]);
  or _18135_ (_09789_, _09788_, _09787_);
  and _18136_ (_09790_, _09789_, _09751_);
  and _18137_ (_09791_, _09750_, word_in[18]);
  or _18138_ (_09792_, _09791_, _09765_);
  or _18139_ (_09793_, _09792_, _09790_);
  or _18140_ (_09794_, _09769_, _08411_);
  and _18141_ (_08645_, _09794_, _09793_);
  not _18142_ (_09795_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _18143_ (_09796_, _09755_, _09795_);
  and _18144_ (_09797_, _09755_, word_in[3]);
  or _18145_ (_09798_, _09797_, _09796_);
  and _18146_ (_09799_, _09798_, _09753_);
  and _18147_ (_09800_, _09752_, word_in[11]);
  or _18148_ (_09801_, _09800_, _09799_);
  and _18149_ (_09802_, _09801_, _09751_);
  and _18150_ (_09803_, _09750_, word_in[19]);
  or _18151_ (_09804_, _09803_, _09765_);
  or _18152_ (_09805_, _09804_, _09802_);
  or _18153_ (_09806_, _09769_, _08425_);
  and _18154_ (_08650_, _09806_, _09805_);
  not _18155_ (_09807_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _18156_ (_09808_, _09755_, _09807_);
  and _18157_ (_09809_, _09755_, word_in[4]);
  or _18158_ (_09810_, _09809_, _09808_);
  and _18159_ (_09811_, _09810_, _09753_);
  and _18160_ (_09812_, _09752_, word_in[12]);
  or _18161_ (_09813_, _09812_, _09811_);
  and _18162_ (_09814_, _09813_, _09751_);
  and _18163_ (_09815_, _09750_, word_in[20]);
  or _18164_ (_09816_, _09815_, _09765_);
  or _18165_ (_09817_, _09816_, _09814_);
  or _18166_ (_09818_, _09769_, _08439_);
  and _18167_ (_13433_, _09818_, _09817_);
  not _18168_ (_09819_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _18169_ (_09820_, _09755_, _09819_);
  and _18170_ (_09821_, _09755_, word_in[5]);
  or _18171_ (_09822_, _09821_, _09820_);
  and _18172_ (_09823_, _09822_, _09753_);
  and _18173_ (_09824_, _09752_, word_in[13]);
  or _18174_ (_09825_, _09824_, _09823_);
  and _18175_ (_09826_, _09825_, _09751_);
  and _18176_ (_09827_, _09750_, word_in[21]);
  or _18177_ (_09828_, _09827_, _09765_);
  or _18178_ (_09829_, _09828_, _09826_);
  or _18179_ (_09830_, _09769_, _08453_);
  and _18180_ (_13434_, _09830_, _09829_);
  not _18181_ (_09831_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _18182_ (_09832_, _09755_, _09831_);
  and _18183_ (_09833_, _09755_, word_in[6]);
  or _18184_ (_09834_, _09833_, _09832_);
  and _18185_ (_09835_, _09834_, _09753_);
  and _18186_ (_09836_, _09752_, word_in[14]);
  or _18187_ (_09837_, _09836_, _09835_);
  and _18188_ (_09838_, _09837_, _09751_);
  and _18189_ (_09839_, _09750_, word_in[22]);
  or _18190_ (_09840_, _09839_, _09765_);
  or _18191_ (_09841_, _09840_, _09838_);
  or _18192_ (_09842_, _09769_, _08469_);
  and _18193_ (_13435_, _09842_, _09841_);
  nor _18194_ (_09844_, _09755_, _07820_);
  and _18195_ (_09845_, _09755_, word_in[7]);
  or _18196_ (_09846_, _09845_, _09844_);
  and _18197_ (_09847_, _09846_, _09753_);
  and _18198_ (_09848_, _09752_, word_in[15]);
  or _18199_ (_09849_, _09848_, _09847_);
  and _18200_ (_09850_, _09849_, _09751_);
  and _18201_ (_09851_, _09750_, _08023_);
  or _18202_ (_09852_, _09851_, _09765_);
  or _18203_ (_09853_, _09852_, _09850_);
  or _18204_ (_09854_, _09769_, _08028_);
  and _18205_ (_13436_, _09854_, _09853_);
  and _18206_ (_09855_, _08493_, _07813_);
  not _18207_ (_09856_, _09855_);
  or _18208_ (_09857_, _09856_, word_in[8]);
  and _18209_ (_09858_, _08490_, _07992_);
  not _18210_ (_09859_, _09858_);
  not _18211_ (_09860_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _18212_ (_09861_, _08496_, _08008_);
  nor _18213_ (_09862_, _09861_, _09860_);
  and _18214_ (_09863_, _09861_, word_in[0]);
  or _18215_ (_09864_, _09863_, _09862_);
  or _18216_ (_09865_, _09864_, _09855_);
  and _18217_ (_09866_, _09865_, _09859_);
  and _18218_ (_09867_, _09866_, _09857_);
  and _18219_ (_09868_, _09764_, _07775_);
  and _18220_ (_09869_, _09858_, _08370_);
  or _18221_ (_09870_, _09869_, _09868_);
  or _18222_ (_09871_, _09870_, _09867_);
  not _18223_ (_09872_, _09868_);
  or _18224_ (_09873_, _09872_, word_in[24]);
  and _18225_ (_13437_, _09873_, _09871_);
  and _18226_ (_09874_, _09861_, word_in[1]);
  not _18227_ (_09875_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _18228_ (_09876_, _09861_, _09875_);
  nor _18229_ (_09878_, _09876_, _09874_);
  nor _18230_ (_09879_, _09878_, _09855_);
  and _18231_ (_09880_, _09855_, word_in[9]);
  or _18232_ (_09881_, _09880_, _09879_);
  and _18233_ (_09882_, _09881_, _09859_);
  and _18234_ (_09883_, _09858_, _08511_);
  or _18235_ (_09884_, _09883_, _09868_);
  or _18236_ (_09885_, _09884_, _09882_);
  or _18237_ (_09886_, _09872_, word_in[25]);
  and _18238_ (_13438_, _09886_, _09885_);
  not _18239_ (_09887_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _18240_ (_09888_, _09861_, _09887_);
  and _18241_ (_09889_, _09861_, word_in[2]);
  nor _18242_ (_09890_, _09889_, _09888_);
  nor _18243_ (_09891_, _09890_, _09855_);
  and _18244_ (_09892_, _09855_, word_in[10]);
  or _18245_ (_09893_, _09892_, _09891_);
  and _18246_ (_09894_, _09893_, _09859_);
  and _18247_ (_09895_, _09858_, _08525_);
  or _18248_ (_09896_, _09895_, _09868_);
  or _18249_ (_09898_, _09896_, _09894_);
  or _18250_ (_09899_, _09872_, word_in[26]);
  and _18251_ (_13439_, _09899_, _09898_);
  and _18252_ (_09901_, _09861_, word_in[3]);
  not _18253_ (_09903_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _18254_ (_09904_, _09861_, _09903_);
  nor _18255_ (_09906_, _09904_, _09901_);
  nor _18256_ (_09907_, _09906_, _09855_);
  and _18257_ (_09908_, _09855_, word_in[11]);
  or _18258_ (_09909_, _09908_, _09907_);
  and _18259_ (_09910_, _09909_, _09859_);
  and _18260_ (_09911_, _09858_, _08546_);
  or _18261_ (_09912_, _09911_, _09868_);
  or _18262_ (_09913_, _09912_, _09910_);
  or _18263_ (_09914_, _09872_, word_in[27]);
  and _18264_ (_08744_, _09914_, _09913_);
  or _18265_ (_09915_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand _18266_ (_09916_, _06205_, _07167_);
  and _18267_ (_09917_, _09916_, _05110_);
  and _18268_ (_08747_, _09917_, _09915_);
  not _18269_ (_09918_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _18270_ (_09919_, _09861_, _09918_);
  and _18271_ (_09920_, _09861_, word_in[4]);
  nor _18272_ (_09921_, _09920_, _09919_);
  nor _18273_ (_09922_, _09921_, _09855_);
  and _18274_ (_09923_, _09855_, word_in[12]);
  or _18275_ (_09924_, _09923_, _09922_);
  and _18276_ (_09925_, _09924_, _09859_);
  and _18277_ (_09926_, _09858_, _08564_);
  or _18278_ (_09927_, _09926_, _09868_);
  or _18279_ (_09928_, _09927_, _09925_);
  or _18280_ (_09929_, _09872_, word_in[28]);
  and _18281_ (_13440_, _09929_, _09928_);
  not _18282_ (_09930_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _18283_ (_09931_, _09861_, _09930_);
  and _18284_ (_09932_, _09861_, word_in[5]);
  or _18285_ (_09933_, _09932_, _09931_);
  or _18286_ (_09934_, _09933_, _09855_);
  or _18287_ (_09935_, _09856_, word_in[13]);
  and _18288_ (_09936_, _09935_, _09934_);
  or _18289_ (_09937_, _09936_, _09858_);
  or _18290_ (_09938_, _09859_, _08572_);
  and _18291_ (_09939_, _09938_, _09937_);
  or _18292_ (_09940_, _09939_, _09868_);
  or _18293_ (_09941_, _09872_, word_in[29]);
  and _18294_ (_13441_, _09941_, _09940_);
  not _18295_ (_09942_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _18296_ (_09943_, _09861_, _09942_);
  and _18297_ (_09944_, _09861_, word_in[6]);
  nor _18298_ (_09945_, _09944_, _09943_);
  nor _18299_ (_09946_, _09945_, _09855_);
  and _18300_ (_09947_, _09855_, word_in[14]);
  or _18301_ (_09948_, _09947_, _09946_);
  and _18302_ (_09949_, _09948_, _09859_);
  and _18303_ (_09950_, _09858_, _08593_);
  or _18304_ (_09951_, _09950_, _09868_);
  or _18305_ (_09952_, _09951_, _09949_);
  or _18306_ (_09953_, _09872_, word_in[30]);
  and _18307_ (_13442_, _09953_, _09952_);
  and _18308_ (_09954_, _09861_, word_in[7]);
  nor _18309_ (_09955_, _09861_, _07699_);
  nor _18310_ (_09956_, _09955_, _09954_);
  nor _18311_ (_09957_, _09956_, _09855_);
  and _18312_ (_09958_, _09855_, word_in[15]);
  or _18313_ (_09959_, _09958_, _09957_);
  and _18314_ (_09960_, _09959_, _09859_);
  and _18315_ (_09961_, _09858_, _08023_);
  or _18316_ (_09962_, _09961_, _09868_);
  or _18317_ (_09963_, _09962_, _09960_);
  or _18318_ (_09964_, _09872_, word_in[31]);
  and _18319_ (_13443_, _09964_, _09963_);
  and _18320_ (_09965_, _08642_, _07992_);
  not _18321_ (_09966_, _09965_);
  and _18322_ (_09967_, _08630_, _07813_);
  not _18323_ (_09968_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _18324_ (_09969_, _08633_, _07988_);
  nor _18325_ (_09970_, _09969_, _09968_);
  and _18326_ (_09971_, _09969_, _08495_);
  nor _18327_ (_09972_, _09971_, _09970_);
  nor _18328_ (_09973_, _09972_, _09967_);
  and _18329_ (_09974_, _09967_, word_in[8]);
  or _18330_ (_09975_, _09974_, _09973_);
  and _18331_ (_09976_, _09975_, _09966_);
  and _18332_ (_09977_, _09764_, _07746_);
  and _18333_ (_09978_, _09965_, _08370_);
  or _18334_ (_09979_, _09978_, _09977_);
  or _18335_ (_09980_, _09979_, _09976_);
  not _18336_ (_09981_, _09977_);
  or _18337_ (_09982_, _09981_, word_in[24]);
  and _18338_ (_08823_, _09982_, _09980_);
  not _18339_ (_09983_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _18340_ (_09984_, _09969_, _09983_);
  and _18341_ (_09985_, _09969_, _08513_);
  or _18342_ (_09986_, _09985_, _09984_);
  or _18343_ (_09987_, _09986_, _09967_);
  not _18344_ (_09988_, _09967_);
  or _18345_ (_09989_, _09988_, word_in[9]);
  and _18346_ (_09990_, _09989_, _09987_);
  or _18347_ (_09991_, _09990_, _09965_);
  or _18348_ (_09992_, _09966_, _08511_);
  and _18349_ (_09993_, _09992_, _09991_);
  or _18350_ (_09994_, _09993_, _09977_);
  or _18351_ (_09995_, _09981_, word_in[25]);
  and _18352_ (_08826_, _09995_, _09994_);
  not _18353_ (_09996_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor _18354_ (_09997_, _09969_, _09996_);
  and _18355_ (_09998_, _09969_, _08401_);
  nor _18356_ (_09999_, _09998_, _09997_);
  nor _18357_ (_10000_, _09999_, _09967_);
  and _18358_ (_10001_, _09967_, word_in[10]);
  or _18359_ (_10002_, _10001_, _10000_);
  and _18360_ (_10003_, _10002_, _09966_);
  and _18361_ (_10004_, _09965_, _08525_);
  or _18362_ (_10005_, _10004_, _09977_);
  or _18363_ (_10006_, _10005_, _10003_);
  or _18364_ (_10007_, _09981_, word_in[26]);
  and _18365_ (_08829_, _10007_, _10006_);
  not _18366_ (_10008_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor _18367_ (_10009_, _09969_, _10008_);
  and _18368_ (_10010_, _09969_, _08415_);
  nor _18369_ (_10011_, _10010_, _10009_);
  nor _18370_ (_10012_, _10011_, _09967_);
  and _18371_ (_10013_, _09967_, word_in[11]);
  or _18372_ (_10014_, _10013_, _10012_);
  and _18373_ (_10015_, _10014_, _09966_);
  and _18374_ (_10016_, _09965_, _08546_);
  or _18375_ (_10017_, _10016_, _09977_);
  or _18376_ (_10018_, _10017_, _10015_);
  or _18377_ (_10019_, _09981_, word_in[27]);
  and _18378_ (_08832_, _10019_, _10018_);
  or _18379_ (_10020_, _09966_, _08564_);
  not _18380_ (_10021_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _18381_ (_10022_, _09969_, _10021_);
  and _18382_ (_10023_, _09969_, _08429_);
  or _18383_ (_10024_, _10023_, _10022_);
  or _18384_ (_10025_, _10024_, _09967_);
  or _18385_ (_10026_, _09988_, word_in[12]);
  and _18386_ (_10027_, _10026_, _10025_);
  or _18387_ (_10028_, _10027_, _09965_);
  and _18388_ (_10029_, _10028_, _10020_);
  or _18389_ (_10030_, _10029_, _09977_);
  or _18390_ (_10031_, _09981_, word_in[28]);
  and _18391_ (_08835_, _10031_, _10030_);
  or _18392_ (_10032_, _09966_, _08572_);
  not _18393_ (_10033_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor _18394_ (_10034_, _09969_, _10033_);
  and _18395_ (_10035_, _09969_, _08443_);
  or _18396_ (_10036_, _10035_, _10034_);
  or _18397_ (_10037_, _10036_, _09967_);
  or _18398_ (_10038_, _09988_, word_in[13]);
  and _18399_ (_10039_, _10038_, _10037_);
  or _18400_ (_10040_, _10039_, _09965_);
  and _18401_ (_10041_, _10040_, _10032_);
  or _18402_ (_10042_, _10041_, _09977_);
  or _18403_ (_10043_, _09981_, word_in[29]);
  and _18404_ (_08839_, _10043_, _10042_);
  or _18405_ (_10044_, _09988_, word_in[14]);
  not _18406_ (_10045_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _18407_ (_10046_, _09969_, _10045_);
  and _18408_ (_10047_, _09969_, _08457_);
  or _18409_ (_10048_, _10047_, _10046_);
  or _18410_ (_10049_, _10048_, _09967_);
  and _18411_ (_10050_, _10049_, _09966_);
  and _18412_ (_10051_, _10050_, _10044_);
  and _18413_ (_10052_, _09965_, _08593_);
  or _18414_ (_10053_, _10052_, _09977_);
  or _18415_ (_10054_, _10053_, _10051_);
  or _18416_ (_10055_, _09981_, word_in[30]);
  and _18417_ (_08843_, _10055_, _10054_);
  nor _18418_ (_10056_, _09969_, _07814_);
  and _18419_ (_10057_, _09969_, _08011_);
  nor _18420_ (_10058_, _10057_, _10056_);
  nor _18421_ (_10059_, _10058_, _09967_);
  and _18422_ (_10060_, _09967_, word_in[15]);
  or _18423_ (_10061_, _10060_, _10059_);
  and _18424_ (_10062_, _10061_, _09966_);
  and _18425_ (_10063_, _09965_, _08023_);
  or _18426_ (_10064_, _10063_, _09977_);
  or _18427_ (_10065_, _10064_, _10062_);
  or _18428_ (_10066_, _09981_, word_in[31]);
  and _18429_ (_08846_, _10066_, _10065_);
  not _18430_ (_10067_, _08002_);
  or _18431_ (_10068_, _10067_, word_in[8]);
  not _18432_ (_10069_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _18433_ (_10070_, _08010_, _10069_);
  and _18434_ (_10071_, _08495_, _08010_);
  or _18435_ (_10072_, _10071_, _10070_);
  or _18436_ (_10073_, _10072_, _08002_);
  and _18437_ (_10074_, _10073_, _07998_);
  and _18438_ (_10075_, _10074_, _10068_);
  and _18439_ (_10076_, _08370_, _07996_);
  or _18440_ (_10077_, _10076_, _08022_);
  or _18441_ (_10078_, _10077_, _10075_);
  or _18442_ (_10079_, _08925_, _08027_);
  and _18443_ (_08906_, _10079_, _10078_);
  or _18444_ (_10080_, _10067_, word_in[9]);
  not _18445_ (_10081_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor _18446_ (_10082_, _08010_, _10081_);
  and _18447_ (_10083_, _08513_, _08010_);
  or _18448_ (_10084_, _10083_, _10082_);
  or _18449_ (_10085_, _10084_, _08002_);
  and _18450_ (_10086_, _10085_, _07998_);
  and _18451_ (_10087_, _10086_, _10080_);
  and _18452_ (_10088_, _08511_, _07996_);
  or _18453_ (_10089_, _10088_, _08022_);
  or _18454_ (_10090_, _10089_, _10087_);
  or _18455_ (_10091_, _08395_, _08027_);
  and _18456_ (_08909_, _10091_, _10090_);
  not _18457_ (_10092_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _18458_ (_10093_, _08010_, _10092_);
  and _18459_ (_10094_, _08401_, _08010_);
  or _18460_ (_10095_, _10094_, _10093_);
  or _18461_ (_10096_, _10095_, _08002_);
  or _18462_ (_10097_, _10067_, word_in[10]);
  and _18463_ (_10098_, _10097_, _10096_);
  or _18464_ (_10099_, _10098_, _07996_);
  or _18465_ (_10100_, _08525_, _07998_);
  and _18466_ (_10101_, _10100_, _10099_);
  or _18467_ (_10102_, _10101_, _08022_);
  or _18468_ (_10103_, _08411_, _08027_);
  and _18469_ (_08913_, _10103_, _10102_);
  not _18470_ (_10105_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _18471_ (_10106_, _08010_, _10105_);
  and _18472_ (_10107_, _08415_, _08010_);
  nor _18473_ (_10108_, _10107_, _10106_);
  nor _18474_ (_10109_, _10108_, _08002_);
  and _18475_ (_10110_, _08002_, word_in[11]);
  or _18476_ (_10111_, _10110_, _10109_);
  and _18477_ (_10112_, _10111_, _07998_);
  and _18478_ (_10113_, _08546_, _07996_);
  or _18479_ (_10114_, _10113_, _08022_);
  or _18480_ (_10115_, _10114_, _10112_);
  or _18481_ (_10116_, _08425_, _08027_);
  and _18482_ (_08916_, _10116_, _10115_);
  or _18483_ (_10117_, _10067_, word_in[12]);
  not _18484_ (_10118_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor _18485_ (_10119_, _08010_, _10118_);
  and _18486_ (_10120_, _08429_, _08010_);
  or _18487_ (_10121_, _10120_, _10119_);
  or _18488_ (_10122_, _10121_, _08002_);
  and _18489_ (_10123_, _10122_, _07998_);
  and _18490_ (_10124_, _10123_, _10117_);
  and _18491_ (_10125_, _08564_, _07996_);
  or _18492_ (_10126_, _10125_, _08022_);
  or _18493_ (_10127_, _10126_, _10124_);
  or _18494_ (_10128_, _08439_, _08027_);
  and _18495_ (_08920_, _10128_, _10127_);
  and _18496_ (_10129_, _08572_, _07996_);
  and _18497_ (_10130_, _08443_, _08010_);
  not _18498_ (_10131_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor _18499_ (_10132_, _08010_, _10131_);
  nor _18500_ (_10133_, _10132_, _10130_);
  nor _18501_ (_10134_, _10133_, _08002_);
  and _18502_ (_10135_, _08002_, word_in[13]);
  or _18503_ (_10136_, _10135_, _10134_);
  and _18504_ (_10137_, _10136_, _07998_);
  or _18505_ (_10138_, _10137_, _10129_);
  and _18506_ (_10139_, _10138_, _08027_);
  and _18507_ (_10140_, _08453_, _08022_);
  or _18508_ (_08923_, _10140_, _10139_);
  or _18509_ (_10141_, _10067_, word_in[14]);
  not _18510_ (_10142_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _18511_ (_10143_, _08010_, _10142_);
  and _18512_ (_10145_, _08457_, _08010_);
  or _18513_ (_10146_, _10145_, _10143_);
  or _18514_ (_10147_, _10146_, _08002_);
  and _18515_ (_10148_, _10147_, _07998_);
  and _18516_ (_10149_, _10148_, _10141_);
  and _18517_ (_10150_, _08593_, _07996_);
  or _18518_ (_10151_, _10150_, _08022_);
  or _18519_ (_10152_, _10151_, _10149_);
  or _18520_ (_10153_, _08469_, _08027_);
  and _18521_ (_08926_, _10153_, _10152_);
  nor _18522_ (_09231_, _05845_, rst);
  and _18523_ (_10154_, _06624_, _05419_);
  nor _18524_ (_10155_, _05447_, _06121_);
  and _18525_ (_10156_, _10155_, _05794_);
  and _18526_ (_10157_, _10156_, _10154_);
  and _18527_ (_10158_, _10157_, _08272_);
  or _18528_ (_10159_, _10158_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _18529_ (_10160_, _05806_, _05992_);
  and _18530_ (_10161_, _10160_, _06618_);
  and _18531_ (_10162_, _10161_, _05434_);
  not _18532_ (_10163_, _10162_);
  and _18533_ (_10164_, _10163_, _10159_);
  nand _18534_ (_10165_, _10158_, _05872_);
  and _18535_ (_10166_, _10165_, _10164_);
  nor _18536_ (_10167_, _10163_, _05938_);
  or _18537_ (_10168_, _10167_, _10166_);
  and _18538_ (_09234_, _10168_, _05110_);
  nor _18539_ (_10169_, _06173_, _05785_);
  not _18540_ (_10170_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _18541_ (_10171_, _05376_, _10170_);
  nor _18542_ (_10172_, _10171_, _10169_);
  or _18543_ (_10173_, _10172_, _06632_);
  and _18544_ (_10174_, _10173_, _10157_);
  and _18545_ (_10175_, _10160_, _05434_);
  and _18546_ (_10176_, _10175_, _06618_);
  and _18547_ (_10177_, _10176_, _06194_);
  nor _18548_ (_10178_, _05376_, _05485_);
  nand _18549_ (_10179_, _10178_, _10157_);
  nor _18550_ (_10180_, _10176_, _10170_);
  and _18551_ (_10181_, _10180_, _10179_);
  or _18552_ (_10182_, _10181_, _10177_);
  or _18553_ (_10183_, _10182_, _10174_);
  and _18554_ (_09629_, _10183_, _05110_);
  and _18555_ (_10184_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _18556_ (_10185_, _10184_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _18557_ (_10186_, _05711_, _05650_);
  and _18558_ (_10187_, _05575_, _05489_);
  nand _18559_ (_10188_, _05158_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _18560_ (_10189_, _10188_, _10184_);
  or _18561_ (_10190_, _10189_, _10187_);
  or _18562_ (_10191_, _10190_, _10186_);
  and _18563_ (_10192_, _10191_, _10185_);
  or _18564_ (_10193_, _10192_, _10157_);
  or _18565_ (_10194_, _05488_, _06646_);
  nand _18566_ (_10195_, _10194_, _10157_);
  or _18567_ (_10196_, _10195_, _05784_);
  and _18568_ (_10197_, _10196_, _10193_);
  or _18569_ (_10198_, _10197_, _10162_);
  nand _18570_ (_10199_, _10162_, _05841_);
  and _18571_ (_10200_, _10199_, _05110_);
  and _18572_ (_09633_, _10200_, _10198_);
  and _18573_ (_10201_, _10157_, _08133_);
  or _18574_ (_10202_, _10201_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _18575_ (_10203_, _10202_, _10163_);
  nand _18576_ (_10204_, _10201_, _05872_);
  and _18577_ (_10205_, _10204_, _10203_);
  nor _18578_ (_10206_, _10163_, _06054_);
  or _18579_ (_10207_, _10206_, _10205_);
  and _18580_ (_09636_, _10207_, _05110_);
  and _18581_ (_10208_, _05376_, _05485_);
  and _18582_ (_10209_, _10208_, _05782_);
  and _18583_ (_10210_, _10209_, _10157_);
  not _18584_ (_10211_, _10157_);
  nor _18585_ (_10212_, _10178_, _10208_);
  or _18586_ (_10213_, _10212_, _10211_);
  and _18587_ (_10214_, _10213_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  not _18588_ (_10215_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _18589_ (_10216_, _10179_, _10215_);
  or _18590_ (_10217_, _10216_, _10214_);
  or _18591_ (_10218_, _10217_, _10210_);
  and _18592_ (_10219_, _10218_, _10163_);
  nor _18593_ (_10220_, _10163_, _05334_);
  or _18594_ (_10221_, _10220_, _10219_);
  and _18595_ (_09639_, _10221_, _05110_);
  or _18596_ (_10222_, _06384_, _07153_);
  or _18597_ (_10223_, _05473_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _18598_ (_10224_, _10223_, _05110_);
  and _18599_ (_09737_, _10224_, _10222_);
  and _18600_ (_10225_, _07742_, word_in[0]);
  nand _18601_ (_10226_, _07603_, _09436_);
  or _18602_ (_10227_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _18603_ (_10228_, _10227_, _10226_);
  and _18604_ (_10229_, _10228_, _07624_);
  nand _18605_ (_10230_, _07603_, _09649_);
  or _18606_ (_10231_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _18607_ (_10232_, _10231_, _10230_);
  and _18608_ (_10233_, _10232_, _07636_);
  nand _18609_ (_10234_, _07603_, _09860_);
  or _18610_ (_10235_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _18611_ (_10236_, _10235_, _10234_);
  and _18612_ (_10237_, _10236_, _07633_);
  or _18613_ (_10238_, _10237_, _10233_);
  or _18614_ (_10239_, _10238_, _10229_);
  nand _18615_ (_10240_, _07603_, _10069_);
  or _18616_ (_10241_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _18617_ (_10242_, _10241_, _10240_);
  and _18618_ (_10243_, _10242_, _07644_);
  or _18619_ (_10244_, _10243_, _07659_);
  or _18620_ (_10245_, _10244_, _10239_);
  nand _18621_ (_10246_, _07603_, _08499_);
  or _18622_ (_10247_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _18623_ (_10248_, _10247_, _10246_);
  and _18624_ (_10249_, _10248_, _07624_);
  nand _18625_ (_10250_, _07603_, _08765_);
  or _18626_ (_10251_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _18627_ (_10252_, _10251_, _10250_);
  and _18628_ (_10253_, _10252_, _07636_);
  nand _18629_ (_10254_, _07603_, _09021_);
  or _18630_ (_10255_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _18631_ (_10257_, _10255_, _10254_);
  and _18632_ (_10258_, _10257_, _07633_);
  or _18633_ (_10259_, _10258_, _10253_);
  or _18634_ (_10260_, _10259_, _10249_);
  nand _18635_ (_10261_, _07603_, _09222_);
  or _18636_ (_10262_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _18637_ (_10263_, _10262_, _10261_);
  and _18638_ (_10264_, _10263_, _07644_);
  or _18639_ (_10265_, _10264_, _07612_);
  or _18640_ (_10266_, _10265_, _10260_);
  and _18641_ (_10267_, _10266_, _10245_);
  and _18642_ (_10268_, _10267_, _07683_);
  or _18643_ (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _10268_, _10225_);
  nor _18644_ (_10269_, _07683_, _08379_);
  nand _18645_ (_10270_, _07603_, _09456_);
  or _18646_ (_10271_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _18647_ (_10272_, _10271_, _10270_);
  and _18648_ (_10273_, _10272_, _07624_);
  nand _18649_ (_10274_, _07603_, _09875_);
  or _18650_ (_10275_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _18651_ (_10276_, _10275_, _10274_);
  and _18652_ (_10277_, _10276_, _07633_);
  nand _18653_ (_10278_, _07603_, _09667_);
  or _18654_ (_10279_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _18655_ (_10280_, _10279_, _10278_);
  and _18656_ (_10281_, _10280_, _07636_);
  or _18657_ (_10282_, _10281_, _10277_);
  or _18658_ (_10283_, _10282_, _10273_);
  nand _18659_ (_10284_, _07603_, _10081_);
  or _18660_ (_10285_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _18661_ (_10286_, _10285_, _10284_);
  and _18662_ (_10287_, _10286_, _07644_);
  or _18663_ (_10288_, _10287_, _07659_);
  or _18664_ (_10289_, _10288_, _10283_);
  nand _18665_ (_10290_, _07603_, _08515_);
  or _18666_ (_10291_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _18667_ (_10292_, _10291_, _10290_);
  and _18668_ (_10293_, _10292_, _07624_);
  nand _18669_ (_10294_, _07603_, _08779_);
  or _18670_ (_10295_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _18671_ (_10296_, _10295_, _10294_);
  and _18672_ (_10297_, _10296_, _07636_);
  nand _18673_ (_10298_, _07603_, _09035_);
  or _18674_ (_10299_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _18675_ (_10300_, _10299_, _10298_);
  and _18676_ (_10301_, _10300_, _07633_);
  or _18677_ (_10302_, _10301_, _10297_);
  or _18678_ (_10303_, _10302_, _10293_);
  nand _18679_ (_10304_, _07603_, _09239_);
  or _18680_ (_10305_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _18681_ (_10307_, _10305_, _10304_);
  and _18682_ (_10308_, _10307_, _07644_);
  or _18683_ (_10309_, _10308_, _07612_);
  or _18684_ (_10310_, _10309_, _10303_);
  and _18685_ (_10311_, _10310_, _10289_);
  and _18686_ (_10312_, _10311_, _07683_);
  or _18687_ (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _10312_, _10269_);
  and _18688_ (_10313_, _07742_, word_in[2]);
  nand _18689_ (_10314_, _07603_, _09471_);
  or _18690_ (_10315_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _18691_ (_10316_, _10315_, _10314_);
  and _18692_ (_10317_, _10316_, _07624_);
  nand _18693_ (_10318_, _07603_, _09680_);
  or _18694_ (_10319_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _18695_ (_10320_, _10319_, _10318_);
  and _18696_ (_10321_, _10320_, _07636_);
  nand _18697_ (_10322_, _07603_, _09887_);
  or _18698_ (_10323_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _18699_ (_10324_, _10323_, _10322_);
  and _18700_ (_10325_, _10324_, _07633_);
  or _18701_ (_10326_, _10325_, _10321_);
  or _18702_ (_10327_, _10326_, _10317_);
  nand _18703_ (_10328_, _07603_, _10092_);
  or _18704_ (_10329_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _18705_ (_10330_, _10329_, _10328_);
  and _18706_ (_10331_, _10330_, _07644_);
  or _18707_ (_10332_, _10331_, _07659_);
  or _18708_ (_10333_, _10332_, _10327_);
  nand _18709_ (_10334_, _07603_, _08528_);
  or _18710_ (_10335_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _18711_ (_10336_, _10335_, _10334_);
  and _18712_ (_10337_, _10336_, _07624_);
  nand _18713_ (_10338_, _07603_, _08791_);
  or _18714_ (_10339_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _18715_ (_10340_, _10339_, _10338_);
  and _18716_ (_10341_, _10340_, _07636_);
  nand _18717_ (_10342_, _07603_, _09048_);
  or _18718_ (_10343_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _18719_ (_10344_, _10343_, _10342_);
  and _18720_ (_10345_, _10344_, _07633_);
  or _18721_ (_10346_, _10345_, _10341_);
  or _18722_ (_10347_, _10346_, _10337_);
  nand _18723_ (_10348_, _07603_, _09252_);
  or _18724_ (_10349_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _18725_ (_10350_, _10349_, _10348_);
  and _18726_ (_10351_, _10350_, _07644_);
  or _18727_ (_10352_, _10351_, _07612_);
  or _18728_ (_10353_, _10352_, _10347_);
  and _18729_ (_10354_, _10353_, _10333_);
  and _18730_ (_10355_, _10354_, _07683_);
  or _18731_ (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _10355_, _10313_);
  and _18732_ (_10356_, _07742_, word_in[3]);
  nand _18733_ (_10357_, _07603_, _09482_);
  or _18734_ (_10358_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _18735_ (_10359_, _10358_, _10357_);
  and _18736_ (_10360_, _10359_, _07624_);
  nand _18737_ (_10361_, _07603_, _09692_);
  or _18738_ (_10362_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _18739_ (_10363_, _10362_, _10361_);
  and _18740_ (_10364_, _10363_, _07636_);
  nand _18741_ (_10365_, _07603_, _09903_);
  or _18742_ (_10366_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and _18743_ (_10367_, _10366_, _10365_);
  and _18744_ (_10368_, _10367_, _07633_);
  or _18745_ (_10369_, _10368_, _10364_);
  or _18746_ (_10370_, _10369_, _10360_);
  nand _18747_ (_10371_, _07603_, _10105_);
  or _18748_ (_10372_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _18749_ (_10373_, _10372_, _10371_);
  and _18750_ (_10374_, _10373_, _07644_);
  or _18751_ (_10375_, _10374_, _07659_);
  or _18752_ (_10376_, _10375_, _10370_);
  nand _18753_ (_10377_, _07603_, _08538_);
  or _18754_ (_10378_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _18755_ (_10379_, _10378_, _10377_);
  and _18756_ (_10380_, _10379_, _07624_);
  nand _18757_ (_10381_, _07603_, _08803_);
  or _18758_ (_10382_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _18759_ (_10383_, _10382_, _10381_);
  and _18760_ (_10384_, _10383_, _07636_);
  nand _18761_ (_10386_, _07603_, _09059_);
  or _18762_ (_10387_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _18763_ (_10388_, _10387_, _10386_);
  and _18764_ (_10389_, _10388_, _07633_);
  or _18765_ (_10390_, _10389_, _10384_);
  or _18766_ (_10391_, _10390_, _10380_);
  nand _18767_ (_10392_, _07603_, _09264_);
  or _18768_ (_10393_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _18769_ (_10394_, _10393_, _10392_);
  and _18770_ (_10395_, _10394_, _07644_);
  or _18771_ (_10396_, _10395_, _07612_);
  or _18772_ (_10397_, _10396_, _10391_);
  and _18773_ (_10398_, _10397_, _10376_);
  and _18774_ (_10399_, _10398_, _07683_);
  or _18775_ (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _10399_, _10356_);
  and _18776_ (_10401_, _07742_, word_in[4]);
  nand _18777_ (_10402_, _07603_, _09494_);
  or _18778_ (_10403_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _18779_ (_10404_, _10403_, _10402_);
  and _18780_ (_10405_, _10404_, _07624_);
  nand _18781_ (_10407_, _07603_, _09703_);
  or _18782_ (_10408_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _18783_ (_10409_, _10408_, _10407_);
  and _18784_ (_10410_, _10409_, _07636_);
  nand _18785_ (_10411_, _07603_, _09918_);
  or _18786_ (_10412_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and _18787_ (_10413_, _10412_, _10411_);
  and _18788_ (_10414_, _10413_, _07633_);
  or _18789_ (_10415_, _10414_, _10410_);
  or _18790_ (_10416_, _10415_, _10405_);
  nand _18791_ (_10417_, _07603_, _10118_);
  or _18792_ (_10418_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _18793_ (_10419_, _10418_, _10417_);
  and _18794_ (_10420_, _10419_, _07644_);
  or _18795_ (_10421_, _10420_, _07659_);
  or _18796_ (_10422_, _10421_, _10416_);
  nand _18797_ (_10423_, _07603_, _08553_);
  or _18798_ (_10424_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _18799_ (_10425_, _10424_, _10423_);
  and _18800_ (_10426_, _10425_, _07624_);
  nand _18801_ (_10428_, _07603_, _08815_);
  or _18802_ (_10429_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _18803_ (_10430_, _10429_, _10428_);
  and _18804_ (_10431_, _10430_, _07636_);
  nand _18805_ (_10432_, _07603_, _09071_);
  or _18806_ (_10433_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _18807_ (_10434_, _10433_, _10432_);
  and _18808_ (_10435_, _10434_, _07633_);
  or _18809_ (_10436_, _10435_, _10431_);
  or _18810_ (_10437_, _10436_, _10426_);
  nand _18811_ (_10438_, _07603_, _09276_);
  or _18812_ (_10439_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _18813_ (_10440_, _10439_, _10438_);
  and _18814_ (_10441_, _10440_, _07644_);
  or _18815_ (_10442_, _10441_, _07612_);
  or _18816_ (_10443_, _10442_, _10437_);
  and _18817_ (_10444_, _10443_, _10422_);
  and _18818_ (_10445_, _10444_, _07683_);
  or _18819_ (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _10445_, _10401_);
  and _18820_ (_10446_, _07742_, word_in[5]);
  nand _18821_ (_10447_, _07603_, _09506_);
  or _18822_ (_10448_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _18823_ (_10449_, _10448_, _10447_);
  and _18824_ (_10450_, _10449_, _07624_);
  nand _18825_ (_10451_, _07603_, _09930_);
  or _18826_ (_10452_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _18827_ (_10453_, _10452_, _10451_);
  and _18828_ (_10454_, _10453_, _07633_);
  nand _18829_ (_10455_, _07603_, _09716_);
  or _18830_ (_10456_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _18831_ (_10457_, _10456_, _10455_);
  and _18832_ (_10458_, _10457_, _07636_);
  or _18833_ (_10459_, _10458_, _10454_);
  or _18834_ (_10461_, _10459_, _10450_);
  nand _18835_ (_10462_, _07603_, _10131_);
  or _18836_ (_10463_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _18837_ (_10464_, _10463_, _10462_);
  and _18838_ (_10465_, _10464_, _07644_);
  or _18839_ (_10466_, _10465_, _07659_);
  or _18840_ (_10467_, _10466_, _10461_);
  nand _18841_ (_10468_, _07603_, _08575_);
  or _18842_ (_10469_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _18843_ (_10470_, _10469_, _10468_);
  and _18844_ (_10471_, _10470_, _07624_);
  nand _18845_ (_10473_, _07603_, _08830_);
  or _18846_ (_10474_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _18847_ (_10475_, _10474_, _10473_);
  and _18848_ (_10476_, _10475_, _07636_);
  nand _18849_ (_10477_, _07603_, _09082_);
  or _18850_ (_10478_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _18851_ (_10479_, _10478_, _10477_);
  and _18852_ (_10480_, _10479_, _07633_);
  or _18853_ (_10481_, _10480_, _10476_);
  or _18854_ (_10482_, _10481_, _10471_);
  nand _18855_ (_10483_, _07603_, _09288_);
  or _18856_ (_10484_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _18857_ (_10485_, _10484_, _10483_);
  and _18858_ (_10486_, _10485_, _07644_);
  or _18859_ (_10487_, _10486_, _07612_);
  or _18860_ (_10488_, _10487_, _10482_);
  and _18861_ (_10489_, _10488_, _10467_);
  and _18862_ (_10490_, _10489_, _07683_);
  or _18863_ (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _10490_, _10446_);
  and _18864_ (_10491_, _07742_, word_in[6]);
  nand _18865_ (_10492_, _07603_, _09518_);
  or _18866_ (_10493_, _07603_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _18867_ (_10494_, _10493_, _10492_);
  and _18868_ (_10495_, _10494_, _07624_);
  nand _18869_ (_10496_, _07603_, _09942_);
  or _18870_ (_10497_, _07603_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _18871_ (_10498_, _10497_, _10496_);
  and _18872_ (_10499_, _10498_, _07633_);
  nand _18873_ (_10500_, _07603_, _09728_);
  or _18874_ (_10501_, _07603_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _18875_ (_10502_, _10501_, _10500_);
  and _18876_ (_10503_, _10502_, _07636_);
  or _18877_ (_10504_, _10503_, _10499_);
  or _18878_ (_10505_, _10504_, _10495_);
  nand _18879_ (_10506_, _07603_, _10142_);
  or _18880_ (_10507_, _07603_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _18881_ (_10508_, _10507_, _10506_);
  and _18882_ (_10509_, _10508_, _07644_);
  or _18883_ (_10510_, _10509_, _07659_);
  or _18884_ (_10511_, _10510_, _10505_);
  nand _18885_ (_10512_, _07603_, _08585_);
  or _18886_ (_10513_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _18887_ (_10514_, _10513_, _10512_);
  and _18888_ (_10515_, _10514_, _07624_);
  nand _18889_ (_10516_, _07603_, _08847_);
  or _18890_ (_10518_, _07603_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _18891_ (_10519_, _10518_, _10516_);
  and _18892_ (_10520_, _10519_, _07636_);
  nand _18893_ (_10521_, _07603_, _09095_);
  or _18894_ (_10522_, _07603_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _18895_ (_10523_, _10522_, _10521_);
  and _18896_ (_10525_, _10523_, _07633_);
  or _18897_ (_10526_, _10525_, _10520_);
  or _18898_ (_10527_, _10526_, _10515_);
  nand _18899_ (_10528_, _07603_, _09300_);
  or _18900_ (_10529_, _07603_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _18901_ (_10530_, _10529_, _10528_);
  and _18902_ (_10531_, _10530_, _07644_);
  or _18903_ (_10532_, _10531_, _07612_);
  or _18904_ (_10533_, _10532_, _10527_);
  and _18905_ (_10534_, _10533_, _10511_);
  and _18906_ (_10535_, _10534_, _07683_);
  or _18907_ (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _10535_, _10491_);
  and _18908_ (_10536_, _07793_, word_in[8]);
  nand _18909_ (_10537_, _07603_, _09543_);
  or _18910_ (_10538_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _18911_ (_10540_, _10538_, _10537_);
  and _18912_ (_10541_, _10540_, _07796_);
  nand _18913_ (_10542_, _07603_, _09335_);
  or _18914_ (_10543_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _18915_ (_10544_, _10543_, _10542_);
  and _18916_ (_10545_, _10544_, _07794_);
  or _18917_ (_10546_, _10545_, _10541_);
  and _18918_ (_10547_, _10546_, _07757_);
  nand _18919_ (_10548_, _07603_, _08637_);
  or _18920_ (_10549_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _18921_ (_10550_, _10549_, _10548_);
  and _18922_ (_10551_, _10550_, _07796_);
  nand _18923_ (_10552_, _07603_, _08350_);
  or _18924_ (_10553_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _18925_ (_10554_, _10553_, _10552_);
  and _18926_ (_10555_, _10554_, _07794_);
  or _18927_ (_10556_, _10555_, _10551_);
  and _18928_ (_10557_, _10556_, _07760_);
  nand _18929_ (_10559_, _07603_, _09118_);
  or _18930_ (_10560_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _18931_ (_10561_, _10560_, _10559_);
  and _18932_ (_10563_, _10561_, _07796_);
  nand _18933_ (_10564_, _07603_, _08907_);
  or _18934_ (_10565_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _18935_ (_10566_, _10565_, _10564_);
  and _18936_ (_10568_, _10566_, _07794_);
  or _18937_ (_10569_, _10568_, _10563_);
  and _18938_ (_10570_, _10569_, _07841_);
  or _18939_ (_10571_, _10570_, _10557_);
  nand _18940_ (_10572_, _07603_, _09968_);
  or _18941_ (_10573_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _18942_ (_10574_, _10573_, _10572_);
  and _18943_ (_10575_, _10574_, _07796_);
  nand _18944_ (_10576_, _07603_, _09754_);
  or _18945_ (_10577_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _18946_ (_10578_, _10577_, _10576_);
  and _18947_ (_10579_, _10578_, _07794_);
  or _18948_ (_10580_, _10579_, _10575_);
  and _18949_ (_10581_, _10580_, _07813_);
  or _18950_ (_10583_, _10581_, _10571_);
  nor _18951_ (_10584_, _10583_, _10547_);
  nor _18952_ (_10586_, _10584_, _07793_);
  or _18953_ (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _10586_, _10536_);
  and _18954_ (_10588_, _07793_, word_in[9]);
  nand _18955_ (_10589_, _07603_, _09559_);
  or _18956_ (_10590_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _18957_ (_10591_, _10590_, _10589_);
  and _18958_ (_10592_, _10591_, _07796_);
  nand _18959_ (_10593_, _07603_, _09351_);
  or _18960_ (_10594_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _18961_ (_10595_, _10594_, _10593_);
  and _18962_ (_10596_, _10595_, _07794_);
  or _18963_ (_10598_, _10596_, _10592_);
  and _18964_ (_10599_, _10598_, _07757_);
  nand _18965_ (_10601_, _07603_, _08659_);
  or _18966_ (_10602_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _18967_ (_10603_, _10602_, _10601_);
  and _18968_ (_10604_, _10603_, _07796_);
  and _18969_ (_10605_, _07603_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _18970_ (_10606_, _07603_, _08515_);
  or _18971_ (_10607_, _10606_, _10605_);
  and _18972_ (_10608_, _10607_, _07794_);
  or _18973_ (_10609_, _10608_, _10604_);
  and _18974_ (_10610_, _10609_, _07760_);
  nand _18975_ (_10611_, _07603_, _09136_);
  or _18976_ (_10612_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _18977_ (_10613_, _10612_, _10611_);
  and _18978_ (_10614_, _10613_, _07796_);
  nand _18979_ (_10615_, _07603_, _08929_);
  or _18980_ (_10616_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _18981_ (_10617_, _10616_, _10615_);
  and _18982_ (_10618_, _10617_, _07794_);
  or _18983_ (_10619_, _10618_, _10614_);
  and _18984_ (_10621_, _10619_, _07841_);
  or _18985_ (_10622_, _10621_, _10610_);
  nand _18986_ (_10623_, _07603_, _09983_);
  or _18987_ (_10624_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _18988_ (_10625_, _10624_, _10623_);
  and _18989_ (_10626_, _10625_, _07796_);
  nand _18990_ (_10627_, _07603_, _09771_);
  or _18991_ (_10628_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _18992_ (_10629_, _10628_, _10627_);
  and _18993_ (_10630_, _10629_, _07794_);
  or _18994_ (_10631_, _10630_, _10626_);
  and _18995_ (_10632_, _10631_, _07813_);
  or _18996_ (_10633_, _10632_, _10622_);
  nor _18997_ (_10634_, _10633_, _10599_);
  nor _18998_ (_10635_, _10634_, _07793_);
  or _18999_ (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _10635_, _10588_);
  and _19000_ (_10636_, _07793_, word_in[10]);
  nand _19001_ (_10637_, _07603_, _09572_);
  or _19002_ (_10638_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _19003_ (_10639_, _10638_, _10637_);
  and _19004_ (_10640_, _10639_, _07796_);
  nand _19005_ (_10642_, _07603_, _09363_);
  or _19006_ (_10643_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _19007_ (_10644_, _10643_, _10642_);
  and _19008_ (_10646_, _10644_, _07794_);
  or _19009_ (_10647_, _10646_, _10640_);
  and _19010_ (_10648_, _10647_, _07757_);
  nand _19011_ (_10650_, _07603_, _08671_);
  or _19012_ (_10651_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _19013_ (_10652_, _10651_, _10650_);
  and _19014_ (_10653_, _10652_, _07796_);
  nand _19015_ (_10655_, _07603_, _08398_);
  or _19016_ (_10656_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _19017_ (_10657_, _10656_, _10655_);
  and _19018_ (_10658_, _10657_, _07794_);
  or _19019_ (_10659_, _10658_, _10653_);
  and _19020_ (_10661_, _10659_, _07760_);
  nand _19021_ (_10662_, _07603_, _09148_);
  or _19022_ (_10664_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _19023_ (_10665_, _10664_, _10662_);
  and _19024_ (_10666_, _10665_, _07796_);
  nand _19025_ (_10667_, _07603_, _08941_);
  or _19026_ (_10668_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _19027_ (_10669_, _10668_, _10667_);
  and _19028_ (_10670_, _10669_, _07794_);
  or _19029_ (_10671_, _10670_, _10666_);
  and _19030_ (_10672_, _10671_, _07841_);
  or _19031_ (_10673_, _10672_, _10661_);
  nand _19032_ (_10674_, _07603_, _09996_);
  or _19033_ (_10675_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _19034_ (_10676_, _10675_, _10674_);
  and _19035_ (_10677_, _10676_, _07796_);
  nand _19036_ (_10678_, _07603_, _09783_);
  or _19037_ (_10680_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and _19038_ (_10681_, _10680_, _10678_);
  and _19039_ (_10682_, _10681_, _07794_);
  or _19040_ (_10683_, _10682_, _10677_);
  and _19041_ (_10685_, _10683_, _07813_);
  or _19042_ (_10686_, _10685_, _10673_);
  nor _19043_ (_10687_, _10686_, _10648_);
  nor _19044_ (_10688_, _10687_, _07793_);
  or _19045_ (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _10688_, _10636_);
  and _19046_ (_10689_, _07793_, word_in[11]);
  nand _19047_ (_10690_, _07603_, _09585_);
  or _19048_ (_10691_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _19049_ (_10692_, _10691_, _10690_);
  and _19050_ (_10693_, _10692_, _07796_);
  nand _19051_ (_10694_, _07603_, _09375_);
  or _19052_ (_10695_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _19053_ (_10696_, _10695_, _10694_);
  and _19054_ (_10698_, _10696_, _07794_);
  or _19055_ (_10699_, _10698_, _10693_);
  and _19056_ (_10700_, _10699_, _07757_);
  nand _19057_ (_10701_, _07603_, _10008_);
  or _19058_ (_10702_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _19059_ (_10703_, _10702_, _10701_);
  and _19060_ (_10704_, _10703_, _07796_);
  nand _19061_ (_10706_, _07603_, _09795_);
  or _19062_ (_10707_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _19063_ (_10708_, _10707_, _10706_);
  and _19064_ (_10710_, _10708_, _07794_);
  or _19065_ (_10711_, _10710_, _10704_);
  and _19066_ (_10713_, _10711_, _07813_);
  nand _19067_ (_10715_, _07603_, _09160_);
  or _19068_ (_10716_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _19069_ (_10718_, _10716_, _10715_);
  and _19070_ (_10719_, _10718_, _07796_);
  nand _19071_ (_10721_, _07603_, _08953_);
  or _19072_ (_10722_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and _19073_ (_10723_, _10722_, _10721_);
  and _19074_ (_10725_, _10723_, _07794_);
  or _19075_ (_10726_, _10725_, _10719_);
  and _19076_ (_10727_, _10726_, _07841_);
  nand _19077_ (_10728_, _07603_, _08683_);
  or _19078_ (_10729_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _19079_ (_10731_, _10729_, _10728_);
  and _19080_ (_10732_, _10731_, _07796_);
  nand _19081_ (_10733_, _07603_, _08413_);
  or _19082_ (_10734_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _19083_ (_10735_, _10734_, _10733_);
  and _19084_ (_10737_, _10735_, _07794_);
  or _19085_ (_10738_, _10737_, _10732_);
  and _19086_ (_10740_, _10738_, _07760_);
  or _19087_ (_10741_, _10740_, _10727_);
  or _19088_ (_10742_, _10741_, _10713_);
  nor _19089_ (_10743_, _10742_, _10700_);
  nor _19090_ (_10744_, _10743_, _07793_);
  or _19091_ (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _10744_, _10689_);
  and _19092_ (_10745_, _07793_, word_in[12]);
  nand _19093_ (_10747_, _07603_, _09598_);
  or _19094_ (_10748_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _19095_ (_10749_, _10748_, _10747_);
  and _19096_ (_10750_, _10749_, _07796_);
  nand _19097_ (_10751_, _07603_, _09387_);
  or _19098_ (_10752_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _19099_ (_10753_, _10752_, _10751_);
  and _19100_ (_10754_, _10753_, _07794_);
  or _19101_ (_10756_, _10754_, _10750_);
  and _19102_ (_10757_, _10756_, _07757_);
  nand _19103_ (_10758_, _07603_, _08696_);
  or _19104_ (_10759_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _19105_ (_10760_, _10759_, _10758_);
  and _19106_ (_10761_, _10760_, _07796_);
  nand _19107_ (_10762_, _07603_, _08427_);
  or _19108_ (_10763_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _19109_ (_10764_, _10763_, _10762_);
  and _19110_ (_10765_, _10764_, _07794_);
  or _19111_ (_10766_, _10765_, _10761_);
  and _19112_ (_10767_, _10766_, _07760_);
  nand _19113_ (_10768_, _07603_, _09172_);
  or _19114_ (_10769_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _19115_ (_10770_, _10769_, _10768_);
  and _19116_ (_10771_, _10770_, _07796_);
  nand _19117_ (_10772_, _07603_, _08965_);
  or _19118_ (_10773_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _19119_ (_10774_, _10773_, _10772_);
  and _19120_ (_10775_, _10774_, _07794_);
  or _19121_ (_10776_, _10775_, _10771_);
  and _19122_ (_10777_, _10776_, _07841_);
  or _19123_ (_10778_, _10777_, _10767_);
  nand _19124_ (_10779_, _07603_, _10021_);
  or _19125_ (_10780_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _19126_ (_10781_, _10780_, _10779_);
  and _19127_ (_10782_, _10781_, _07796_);
  nand _19128_ (_10783_, _07603_, _09807_);
  or _19129_ (_10785_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _19130_ (_10786_, _10785_, _10783_);
  and _19131_ (_10787_, _10786_, _07794_);
  or _19132_ (_10788_, _10787_, _10782_);
  and _19133_ (_10790_, _10788_, _07813_);
  or _19134_ (_10791_, _10790_, _10778_);
  nor _19135_ (_10792_, _10791_, _10757_);
  nor _19136_ (_10793_, _10792_, _07793_);
  or _19137_ (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _10793_, _10745_);
  and _19138_ (_10794_, _07793_, word_in[13]);
  nand _19139_ (_10795_, _07603_, _09608_);
  or _19140_ (_10796_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _19141_ (_10797_, _10796_, _10795_);
  and _19142_ (_10798_, _10797_, _07796_);
  nand _19143_ (_10799_, _07603_, _09399_);
  or _19144_ (_10800_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _19145_ (_10801_, _10800_, _10799_);
  and _19146_ (_10802_, _10801_, _07794_);
  or _19147_ (_10804_, _10802_, _10798_);
  and _19148_ (_10805_, _10804_, _07757_);
  nand _19149_ (_10806_, _07603_, _08708_);
  or _19150_ (_10807_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _19151_ (_10808_, _10807_, _10806_);
  and _19152_ (_10809_, _10808_, _07796_);
  nand _19153_ (_10810_, _07603_, _08441_);
  or _19154_ (_10811_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _19155_ (_10812_, _10811_, _10810_);
  and _19156_ (_10814_, _10812_, _07794_);
  or _19157_ (_10815_, _10814_, _10809_);
  and _19158_ (_10816_, _10815_, _07760_);
  nand _19159_ (_10817_, _07603_, _09184_);
  or _19160_ (_10818_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _19161_ (_10819_, _10818_, _10817_);
  and _19162_ (_10820_, _10819_, _07796_);
  nand _19163_ (_10821_, _07603_, _08977_);
  or _19164_ (_10822_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _19165_ (_10823_, _10822_, _10821_);
  and _19166_ (_10824_, _10823_, _07794_);
  or _19167_ (_10825_, _10824_, _10820_);
  and _19168_ (_10826_, _10825_, _07841_);
  or _19169_ (_10827_, _10826_, _10816_);
  nand _19170_ (_10828_, _07603_, _10033_);
  or _19171_ (_10829_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _19172_ (_10830_, _10829_, _10828_);
  and _19173_ (_10831_, _10830_, _07796_);
  nand _19174_ (_10832_, _07603_, _09819_);
  or _19175_ (_10833_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _19176_ (_10834_, _10833_, _10832_);
  and _19177_ (_10835_, _10834_, _07794_);
  or _19178_ (_10836_, _10835_, _10831_);
  and _19179_ (_10837_, _10836_, _07813_);
  or _19180_ (_10838_, _10837_, _10827_);
  nor _19181_ (_10839_, _10838_, _10805_);
  nor _19182_ (_10840_, _10839_, _07793_);
  or _19183_ (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _10840_, _10794_);
  and _19184_ (_10841_, _07793_, word_in[14]);
  nand _19185_ (_10842_, _07603_, _09621_);
  or _19186_ (_10843_, _07603_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _19187_ (_10844_, _10843_, _10842_);
  and _19188_ (_10845_, _10844_, _07796_);
  nand _19189_ (_10846_, _07603_, _09411_);
  or _19190_ (_10847_, _07603_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _19191_ (_10848_, _10847_, _10846_);
  and _19192_ (_10849_, _10848_, _07794_);
  or _19193_ (_10850_, _10849_, _10845_);
  and _19194_ (_10851_, _10850_, _07757_);
  nand _19195_ (_10852_, _07603_, _10045_);
  or _19196_ (_10853_, _07603_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _19197_ (_10854_, _10853_, _10852_);
  and _19198_ (_10855_, _10854_, _07796_);
  nand _19199_ (_10856_, _07603_, _09831_);
  or _19200_ (_10857_, _07603_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _19201_ (_10858_, _10857_, _10856_);
  and _19202_ (_10859_, _10858_, _07794_);
  or _19203_ (_10860_, _10859_, _10855_);
  and _19204_ (_10861_, _10860_, _07813_);
  nand _19205_ (_10863_, _07603_, _09197_);
  or _19206_ (_10864_, _07603_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _19207_ (_10865_, _10864_, _10863_);
  and _19208_ (_10866_, _10865_, _07796_);
  nand _19209_ (_10867_, _07603_, _08990_);
  or _19210_ (_10868_, _07603_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _19211_ (_10869_, _10868_, _10867_);
  and _19212_ (_10870_, _10869_, _07794_);
  or _19213_ (_10871_, _10870_, _10866_);
  and _19214_ (_10872_, _10871_, _07841_);
  nand _19215_ (_10873_, _07603_, _08718_);
  or _19216_ (_10874_, _07603_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _19217_ (_10875_, _10874_, _10873_);
  and _19218_ (_10876_, _10875_, _07796_);
  nand _19219_ (_10877_, _07603_, _08455_);
  or _19220_ (_10878_, _07603_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _19221_ (_10879_, _10878_, _10877_);
  and _19222_ (_10881_, _10879_, _07794_);
  or _19223_ (_10882_, _10881_, _10876_);
  and _19224_ (_10884_, _10882_, _07760_);
  or _19225_ (_10885_, _10884_, _10872_);
  or _19226_ (_10886_, _10885_, _10861_);
  nor _19227_ (_10887_, _10886_, _10851_);
  nor _19228_ (_10888_, _10887_, _07793_);
  or _19229_ (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _10888_, _10841_);
  and _19230_ (_10889_, _07896_, word_in[16]);
  and _19231_ (_10890_, _10232_, _07624_);
  and _19232_ (_10891_, _10236_, _07636_);
  or _19233_ (_10892_, _10891_, _10890_);
  and _19234_ (_10893_, _10242_, _07633_);
  and _19235_ (_10894_, _10228_, _07644_);
  or _19236_ (_10895_, _10894_, _10893_);
  or _19237_ (_10896_, _10895_, _10892_);
  or _19238_ (_10897_, _10896_, _07907_);
  and _19239_ (_10898_, _10257_, _07636_);
  and _19240_ (_10899_, _10248_, _07644_);
  or _19241_ (_10900_, _10899_, _10898_);
  and _19242_ (_10901_, _10263_, _07633_);
  and _19243_ (_10902_, _10252_, _07624_);
  or _19244_ (_10903_, _10902_, _10901_);
  or _19245_ (_10904_, _10903_, _10900_);
  or _19246_ (_10905_, _10904_, _07863_);
  nand _19247_ (_10906_, _10905_, _10897_);
  nor _19248_ (_10907_, _10906_, _07896_);
  or _19249_ (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _10907_, _10889_);
  and _19250_ (_10908_, _07896_, word_in[17]);
  and _19251_ (_10909_, _10286_, _07633_);
  and _19252_ (_10910_, _10280_, _07624_);
  or _19253_ (_10911_, _10910_, _10909_);
  and _19254_ (_10912_, _10276_, _07636_);
  and _19255_ (_10913_, _10272_, _07644_);
  or _19256_ (_10914_, _10913_, _10912_);
  or _19257_ (_10915_, _10914_, _10911_);
  or _19258_ (_10916_, _10915_, _07907_);
  and _19259_ (_10917_, _10307_, _07633_);
  and _19260_ (_10918_, _10300_, _07636_);
  or _19261_ (_10919_, _10918_, _10917_);
  and _19262_ (_10920_, _10296_, _07624_);
  and _19263_ (_10921_, _10292_, _07644_);
  or _19264_ (_10922_, _10921_, _10920_);
  or _19265_ (_10923_, _10922_, _10919_);
  or _19266_ (_10924_, _10923_, _07863_);
  nand _19267_ (_10925_, _10924_, _10916_);
  nor _19268_ (_10926_, _10925_, _07896_);
  or _19269_ (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _10926_, _10908_);
  and _19270_ (_10927_, _07896_, word_in[18]);
  and _19271_ (_10928_, _10350_, _07633_);
  and _19272_ (_10929_, _10340_, _07624_);
  or _19273_ (_10930_, _10929_, _10928_);
  and _19274_ (_10931_, _10344_, _07636_);
  and _19275_ (_10932_, _10336_, _07644_);
  or _19276_ (_10933_, _10932_, _10931_);
  or _19277_ (_10934_, _10933_, _10930_);
  or _19278_ (_10936_, _10934_, _07863_);
  and _19279_ (_10937_, _10320_, _07624_);
  and _19280_ (_10938_, _10324_, _07636_);
  or _19281_ (_10939_, _10938_, _10937_);
  and _19282_ (_10940_, _10330_, _07633_);
  and _19283_ (_10941_, _10316_, _07644_);
  or _19284_ (_10943_, _10941_, _10940_);
  or _19285_ (_10944_, _10943_, _10939_);
  or _19286_ (_10945_, _10944_, _07907_);
  nand _19287_ (_10946_, _10945_, _10936_);
  nor _19288_ (_10947_, _10946_, _07896_);
  or _19289_ (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _10947_, _10927_);
  and _19290_ (_10948_, _07896_, word_in[19]);
  and _19291_ (_10949_, _10363_, _07624_);
  and _19292_ (_10950_, _10367_, _07636_);
  or _19293_ (_10951_, _10950_, _10949_);
  and _19294_ (_10952_, _10373_, _07633_);
  and _19295_ (_10953_, _10359_, _07644_);
  or _19296_ (_10954_, _10953_, _10952_);
  or _19297_ (_10955_, _10954_, _10951_);
  or _19298_ (_10956_, _10955_, _07907_);
  and _19299_ (_10957_, _10388_, _07636_);
  and _19300_ (_10958_, _10379_, _07644_);
  or _19301_ (_10959_, _10958_, _10957_);
  and _19302_ (_10960_, _10394_, _07633_);
  and _19303_ (_10961_, _10383_, _07624_);
  or _19304_ (_10962_, _10961_, _10960_);
  or _19305_ (_10963_, _10962_, _10959_);
  or _19306_ (_10964_, _10963_, _07863_);
  nand _19307_ (_10965_, _10964_, _10956_);
  nor _19308_ (_10967_, _10965_, _07896_);
  or _19309_ (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _10967_, _10948_);
  and _19310_ (_10968_, _07896_, word_in[20]);
  and _19311_ (_10969_, _10430_, _07624_);
  and _19312_ (_10970_, _10425_, _07644_);
  or _19313_ (_10971_, _10970_, _10969_);
  and _19314_ (_10972_, _10440_, _07633_);
  and _19315_ (_10973_, _10434_, _07636_);
  or _19316_ (_10975_, _10973_, _10972_);
  or _19317_ (_10976_, _10975_, _10971_);
  or _19318_ (_10977_, _10976_, _07863_);
  and _19319_ (_10978_, _10409_, _07624_);
  and _19320_ (_10980_, _10404_, _07644_);
  or _19321_ (_10981_, _10980_, _10978_);
  and _19322_ (_10982_, _10419_, _07633_);
  and _19323_ (_10983_, _10413_, _07636_);
  or _19324_ (_10984_, _10983_, _10982_);
  or _19325_ (_10986_, _10984_, _10981_);
  or _19326_ (_10987_, _10986_, _07907_);
  nand _19327_ (_10988_, _10987_, _10977_);
  nor _19328_ (_10989_, _10988_, _07896_);
  or _19329_ (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _10989_, _10968_);
  and _19330_ (_10990_, _07896_, word_in[21]);
  and _19331_ (_10991_, _10475_, _07624_);
  and _19332_ (_10992_, _10470_, _07644_);
  or _19333_ (_10993_, _10992_, _10991_);
  and _19334_ (_10994_, _10485_, _07633_);
  and _19335_ (_10995_, _10479_, _07636_);
  or _19336_ (_10996_, _10995_, _10994_);
  or _19337_ (_10997_, _10996_, _10993_);
  or _19338_ (_10998_, _10997_, _07863_);
  and _19339_ (_10999_, _10464_, _07633_);
  and _19340_ (_11000_, _10457_, _07624_);
  or _19341_ (_11001_, _11000_, _10999_);
  and _19342_ (_11002_, _10453_, _07636_);
  and _19343_ (_11003_, _10449_, _07644_);
  or _19344_ (_11005_, _11003_, _11002_);
  or _19345_ (_11007_, _11005_, _11001_);
  or _19346_ (_11008_, _11007_, _07907_);
  nand _19347_ (_11009_, _11008_, _10998_);
  nor _19348_ (_11010_, _11009_, _07896_);
  or _19349_ (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _11010_, _10990_);
  and _19350_ (_11011_, _07896_, word_in[22]);
  and _19351_ (_11012_, _10508_, _07633_);
  and _19352_ (_11013_, _10502_, _07624_);
  or _19353_ (_11014_, _11013_, _11012_);
  and _19354_ (_11015_, _10498_, _07636_);
  and _19355_ (_11016_, _10494_, _07644_);
  or _19356_ (_11017_, _11016_, _11015_);
  or _19357_ (_11018_, _11017_, _11014_);
  or _19358_ (_11019_, _11018_, _07907_);
  and _19359_ (_11020_, _10523_, _07636_);
  and _19360_ (_11021_, _10514_, _07644_);
  or _19361_ (_11022_, _11021_, _11020_);
  and _19362_ (_11023_, _10530_, _07633_);
  and _19363_ (_11024_, _10519_, _07624_);
  or _19364_ (_11025_, _11024_, _11023_);
  or _19365_ (_11026_, _11025_, _11022_);
  or _19366_ (_11027_, _11026_, _07863_);
  nand _19367_ (_11028_, _11027_, _11019_);
  nor _19368_ (_11029_, _11028_, _07896_);
  or _19369_ (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _11029_, _11011_);
  and _19370_ (_11030_, _07964_, word_in[24]);
  and _19371_ (_11031_, _10544_, _07796_);
  and _19372_ (_11032_, _10540_, _07794_);
  or _19373_ (_11033_, _11032_, _11031_);
  and _19374_ (_11034_, _11033_, _07938_);
  and _19375_ (_11035_, _10554_, _07796_);
  and _19376_ (_11036_, _10550_, _07794_);
  or _19377_ (_11037_, _11036_, _11035_);
  and _19378_ (_11038_, _11037_, _07944_);
  and _19379_ (_11039_, _10566_, _07796_);
  and _19380_ (_11040_, _10561_, _07794_);
  or _19381_ (_11041_, _11040_, _11039_);
  and _19382_ (_11042_, _11041_, _07973_);
  and _19383_ (_11043_, _10578_, _07796_);
  and _19384_ (_11044_, _10574_, _07794_);
  or _19385_ (_11045_, _11044_, _11043_);
  and _19386_ (_11046_, _11045_, _07981_);
  or _19387_ (_11047_, _11046_, _11042_);
  or _19388_ (_11048_, _11047_, _11038_);
  nor _19389_ (_11049_, _11048_, _11034_);
  nor _19390_ (_11050_, _11049_, _07964_);
  or _19391_ (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _11050_, _11030_);
  and _19392_ (_11051_, _07964_, word_in[25]);
  and _19393_ (_11052_, _10595_, _07796_);
  and _19394_ (_11053_, _10591_, _07794_);
  or _19395_ (_11054_, _11053_, _11052_);
  and _19396_ (_11055_, _11054_, _07938_);
  and _19397_ (_11056_, _10607_, _07796_);
  and _19398_ (_11057_, _10603_, _07794_);
  or _19399_ (_11059_, _11057_, _11056_);
  and _19400_ (_11060_, _11059_, _07944_);
  and _19401_ (_11061_, _10617_, _07796_);
  and _19402_ (_11062_, _10613_, _07794_);
  or _19403_ (_11063_, _11062_, _11061_);
  and _19404_ (_11064_, _11063_, _07973_);
  and _19405_ (_11065_, _10629_, _07796_);
  and _19406_ (_11066_, _10625_, _07794_);
  or _19407_ (_11067_, _11066_, _11065_);
  and _19408_ (_11068_, _11067_, _07981_);
  or _19409_ (_11069_, _11068_, _11064_);
  or _19410_ (_11070_, _11069_, _11060_);
  nor _19411_ (_11071_, _11070_, _11055_);
  nor _19412_ (_11072_, _11071_, _07964_);
  or _19413_ (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _11072_, _11051_);
  and _19414_ (_11074_, _07964_, word_in[26]);
  and _19415_ (_11075_, _10657_, _07796_);
  and _19416_ (_11076_, _10652_, _07794_);
  or _19417_ (_11077_, _11076_, _11075_);
  and _19418_ (_11078_, _11077_, _07944_);
  and _19419_ (_11079_, _10644_, _07796_);
  and _19420_ (_11080_, _10639_, _07794_);
  or _19421_ (_11081_, _11080_, _11079_);
  and _19422_ (_11082_, _11081_, _07938_);
  and _19423_ (_11083_, _10669_, _07796_);
  and _19424_ (_11084_, _10665_, _07794_);
  or _19425_ (_11085_, _11084_, _11083_);
  and _19426_ (_11086_, _11085_, _07973_);
  and _19427_ (_11087_, _10681_, _07796_);
  and _19428_ (_11088_, _10676_, _07794_);
  or _19429_ (_11089_, _11088_, _11087_);
  and _19430_ (_11090_, _11089_, _07981_);
  or _19431_ (_11091_, _11090_, _11086_);
  or _19432_ (_11092_, _11091_, _11082_);
  nor _19433_ (_11093_, _11092_, _11078_);
  nor _19434_ (_11094_, _11093_, _07964_);
  or _19435_ (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _11094_, _11074_);
  and _19436_ (_11096_, _07964_, word_in[27]);
  and _19437_ (_11097_, _10696_, _07796_);
  and _19438_ (_11098_, _10692_, _07794_);
  or _19439_ (_11099_, _11098_, _11097_);
  and _19440_ (_11100_, _11099_, _07938_);
  and _19441_ (_11101_, _10735_, _07796_);
  and _19442_ (_11102_, _10731_, _07794_);
  or _19443_ (_11103_, _11102_, _11101_);
  and _19444_ (_11104_, _11103_, _07944_);
  and _19445_ (_11105_, _10723_, _07796_);
  and _19446_ (_11106_, _10718_, _07794_);
  or _19447_ (_11107_, _11106_, _11105_);
  and _19448_ (_11108_, _11107_, _07973_);
  and _19449_ (_11109_, _10708_, _07796_);
  and _19450_ (_11110_, _10703_, _07794_);
  or _19451_ (_11111_, _11110_, _11109_);
  and _19452_ (_11113_, _11111_, _07981_);
  or _19453_ (_11114_, _11113_, _11108_);
  or _19454_ (_11116_, _11114_, _11104_);
  nor _19455_ (_11117_, _11116_, _11100_);
  nor _19456_ (_11118_, _11117_, _07964_);
  or _19457_ (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _11118_, _11096_);
  and _19458_ (_11119_, _07964_, word_in[28]);
  and _19459_ (_11120_, _10753_, _07796_);
  and _19460_ (_11122_, _10749_, _07794_);
  or _19461_ (_11123_, _11122_, _11120_);
  and _19462_ (_11124_, _11123_, _07938_);
  and _19463_ (_11125_, _10764_, _07796_);
  and _19464_ (_11127_, _10760_, _07794_);
  or _19465_ (_11128_, _11127_, _11125_);
  and _19466_ (_11129_, _11128_, _07944_);
  and _19467_ (_11130_, _10774_, _07796_);
  and _19468_ (_11131_, _10770_, _07794_);
  or _19469_ (_11132_, _11131_, _11130_);
  and _19470_ (_11133_, _11132_, _07973_);
  and _19471_ (_11134_, _10786_, _07796_);
  and _19472_ (_11135_, _10781_, _07794_);
  or _19473_ (_11136_, _11135_, _11134_);
  and _19474_ (_11137_, _11136_, _07981_);
  or _19475_ (_11139_, _11137_, _11133_);
  or _19476_ (_11140_, _11139_, _11129_);
  nor _19477_ (_11141_, _11140_, _11124_);
  nor _19478_ (_11142_, _11141_, _07964_);
  or _19479_ (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _11142_, _11119_);
  and _19480_ (_11143_, _07964_, word_in[29]);
  and _19481_ (_11144_, _10801_, _07796_);
  and _19482_ (_11145_, _10797_, _07794_);
  or _19483_ (_11146_, _11145_, _11144_);
  and _19484_ (_11147_, _11146_, _07938_);
  and _19485_ (_11149_, _10812_, _07796_);
  and _19486_ (_11151_, _10808_, _07794_);
  or _19487_ (_11152_, _11151_, _11149_);
  and _19488_ (_11153_, _11152_, _07944_);
  and _19489_ (_11155_, _10823_, _07796_);
  and _19490_ (_11156_, _10819_, _07794_);
  or _19491_ (_11157_, _11156_, _11155_);
  and _19492_ (_11158_, _11157_, _07973_);
  and _19493_ (_11159_, _10834_, _07796_);
  and _19494_ (_11160_, _10830_, _07794_);
  or _19495_ (_11162_, _11160_, _11159_);
  and _19496_ (_11163_, _11162_, _07981_);
  or _19497_ (_11165_, _11163_, _11158_);
  or _19498_ (_11166_, _11165_, _11153_);
  nor _19499_ (_11167_, _11166_, _11147_);
  nor _19500_ (_11168_, _11167_, _07964_);
  or _19501_ (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _11168_, _11143_);
  and _19502_ (_11169_, _07964_, word_in[30]);
  and _19503_ (_11170_, _10848_, _07796_);
  and _19504_ (_11171_, _10844_, _07794_);
  or _19505_ (_11172_, _11171_, _11170_);
  and _19506_ (_11173_, _11172_, _07938_);
  and _19507_ (_11174_, _10879_, _07796_);
  and _19508_ (_11175_, _10875_, _07794_);
  or _19509_ (_11176_, _11175_, _11174_);
  and _19510_ (_11177_, _11176_, _07944_);
  and _19511_ (_11178_, _10869_, _07796_);
  and _19512_ (_11179_, _10865_, _07794_);
  or _19513_ (_11180_, _11179_, _11178_);
  and _19514_ (_11181_, _11180_, _07973_);
  and _19515_ (_11182_, _10858_, _07796_);
  and _19516_ (_11183_, _10854_, _07794_);
  or _19517_ (_11184_, _11183_, _11182_);
  and _19518_ (_11185_, _11184_, _07981_);
  or _19519_ (_11186_, _11185_, _11181_);
  or _19520_ (_11187_, _11186_, _11177_);
  nor _19521_ (_11188_, _11187_, _11173_);
  nor _19522_ (_11189_, _11188_, _07964_);
  or _19523_ (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _11189_, _11169_);
  not _19524_ (_11190_, _06881_);
  not _19525_ (_11191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand _19526_ (_11192_, _06880_, _11191_);
  nor _19527_ (_11193_, _11192_, _11190_);
  not _19528_ (_11194_, _11193_);
  or _19529_ (_11196_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not _19530_ (_11197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _19531_ (_11199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _11197_);
  and _19532_ (_11200_, _11199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _19533_ (_11202_, _11200_, _11196_);
  and _19534_ (_11203_, _11202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _19535_ (_11204_, _11203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _19536_ (_11205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand _19537_ (_11206_, _11205_, _11202_);
  and _19538_ (_11207_, _11206_, _11204_);
  and _19539_ (_11208_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _19540_ (_11209_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _19541_ (_11211_, _11205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _19542_ (_11212_, _11211_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _19543_ (_11213_, _11212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _19544_ (_11214_, _11213_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _19545_ (_11215_, _11214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _19546_ (_11216_, _11215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _19547_ (_11217_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _19548_ (_11218_, _11217_, _11216_);
  and _19549_ (_11219_, _11218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _19550_ (_11220_, _11219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _19551_ (_11222_, _11220_, _11209_);
  and _19552_ (_11223_, _11222_, _11208_);
  not _19553_ (_11225_, _06882_);
  and _19554_ (_11226_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _19555_ (_11227_, _11226_, _11202_);
  and _19556_ (_11228_, _11227_, _11223_);
  or _19557_ (_11230_, _11228_, _11207_);
  and _19558_ (_11231_, _11230_, _11194_);
  and _19559_ (_11232_, _11193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _19560_ (_11233_, _05807_, _10208_);
  and _19561_ (_11234_, _11233_, _06888_);
  or _19562_ (_11235_, _11234_, _11232_);
  or _19563_ (_11236_, _11235_, _11231_);
  nand _19564_ (_11237_, _11234_, _05938_);
  and _19565_ (_11238_, _08133_, _05807_);
  and _19566_ (_11239_, _11238_, _06888_);
  not _19567_ (_11240_, _11239_);
  and _19568_ (_11241_, _11240_, _11237_);
  and _19569_ (_11242_, _11241_, _11236_);
  and _19570_ (_11243_, _11239_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _19571_ (_11245_, _11243_, _11242_);
  and _19572_ (_09843_, _11245_, _05110_);
  or _19573_ (_11246_, _06406_, _07153_);
  or _19574_ (_11247_, _05473_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _19575_ (_11248_, _11247_, _05110_);
  and _19576_ (_09877_, _11248_, _11246_);
  nand _19577_ (_11249_, _06338_, _05473_);
  or _19578_ (_11250_, _05473_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _19579_ (_11251_, _11250_, _05110_);
  and _19580_ (_09897_, _11251_, _11249_);
  nand _19581_ (_11252_, _06427_, _05473_);
  or _19582_ (_11253_, _05473_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _19583_ (_11254_, _11253_, _05110_);
  and _19584_ (_09900_, _11254_, _11252_);
  or _19585_ (_11255_, _06271_, _07153_);
  or _19586_ (_11256_, _05473_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _19587_ (_11257_, _11256_, _05110_);
  and _19588_ (_09902_, _11257_, _11255_);
  nand _19589_ (_11258_, _06315_, _05473_);
  or _19590_ (_11259_, _05473_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _19591_ (_11260_, _11259_, _05110_);
  and _19592_ (_09905_, _11260_, _11258_);
  and _19593_ (_11261_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _19594_ (_11262_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _19595_ (_11263_, _05846_, _11262_);
  not _19596_ (_11264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _19597_ (_11265_, _11264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _19598_ (_11266_, _11265_, _11263_);
  nor _19599_ (_11268_, _11266_, _11261_);
  or _19600_ (_11269_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _19601_ (_11271_, _11269_, _05110_);
  nor _19602_ (_10104_, _11271_, _11268_);
  not _19603_ (_11272_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor _19604_ (_11273_, _05464_, _11272_);
  nor _19605_ (_11274_, _06054_, _05465_);
  or _19606_ (_11275_, _11274_, _11273_);
  and _19607_ (_10144_, _11275_, _05110_);
  not _19608_ (_11276_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _19609_ (_11277_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , _11276_);
  and _19610_ (_10400_, _11277_, _05110_);
  nor _19611_ (_11279_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _19612_ (_11280_, _11279_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _19613_ (_10460_, _11280_, _05110_);
  and _19614_ (_11281_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _19615_ (_11282_, _11281_);
  and _19616_ (_11283_, _07070_, _06451_);
  and _19617_ (_11284_, _11283_, _06873_);
  and _19618_ (_11286_, _11284_, _06342_);
  or _19619_ (_11287_, _07137_, _06823_);
  nor _19620_ (_11288_, _11287_, _07074_);
  and _19621_ (_11289_, _06811_, _06451_);
  and _19622_ (_11290_, _07071_, _06276_);
  or _19623_ (_11292_, _11290_, _07038_);
  and _19624_ (_11293_, _11292_, _06460_);
  nor _19625_ (_11294_, _11293_, _11289_);
  and _19626_ (_11295_, _11294_, _11288_);
  or _19627_ (_11296_, _07087_, _06452_);
  and _19628_ (_11297_, _11296_, _06448_);
  nor _19629_ (_11298_, _11297_, _06449_);
  nor _19630_ (_11299_, _07041_, _06461_);
  nand _19631_ (_11300_, _06852_, _07063_);
  and _19632_ (_11301_, _07038_, _06864_);
  and _19633_ (_11302_, _06825_, _06460_);
  nor _19634_ (_11303_, _11302_, _11301_);
  and _19635_ (_11304_, _11303_, _11300_);
  and _19636_ (_11305_, _11304_, _11299_);
  and _19637_ (_11306_, _11305_, _11298_);
  nand _19638_ (_11307_, _11306_, _11295_);
  and _19639_ (_11308_, _06872_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _19640_ (_11309_, _11301_, _11308_);
  or _19641_ (_11310_, _11309_, _06870_);
  and _19642_ (_11311_, _11310_, _11307_);
  or _19643_ (_11312_, _11311_, _11286_);
  nand _19644_ (_11313_, _11312_, _05151_);
  and _19645_ (_11314_, _11313_, _11282_);
  and _19646_ (_11315_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2]);
  not _19647_ (_11316_, _11315_);
  nand _19648_ (_11317_, _11298_, _06440_);
  nand _19649_ (_11319_, _11317_, _06870_);
  nor _19650_ (_11320_, _11284_, _07056_);
  nand _19651_ (_11321_, _11320_, _11319_);
  nand _19652_ (_11322_, _11321_, _05151_);
  and _19653_ (_11323_, _11322_, _11316_);
  nand _19654_ (_11324_, _11323_, _05110_);
  nor _19655_ (_10472_, _11324_, _11314_);
  nor _19656_ (_11325_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _19657_ (_10517_, _11325_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _19658_ (_11326_, _10155_, _05797_);
  and _19659_ (_11327_, _11326_, _05805_);
  or _19660_ (_11328_, _11327_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _19661_ (_11329_, _06888_, _05808_);
  not _19662_ (_11330_, _11329_);
  and _19663_ (_11331_, _11330_, _11328_);
  nand _19664_ (_11332_, _11327_, _05872_);
  and _19665_ (_11333_, _11332_, _11331_);
  and _19666_ (_11334_, _11329_, _06799_);
  or _19667_ (_11335_, _11334_, _11333_);
  and _19668_ (_10524_, _11335_, _05110_);
  nor _19669_ (_11336_, _06205_, _06200_);
  and _19670_ (_11337_, _06920_, _06909_);
  not _19671_ (_11338_, _11337_);
  and _19672_ (_11339_, _06909_, _06271_);
  not _19673_ (_11340_, _06315_);
  and _19674_ (_11341_, _11340_, _06294_);
  and _19675_ (_11342_, _11341_, _11339_);
  and _19676_ (_11343_, _06338_, _06271_);
  nor _19677_ (_11344_, _06315_, _06294_);
  and _19678_ (_11345_, _11344_, _11343_);
  nor _19679_ (_11346_, _11345_, _11342_);
  and _19680_ (_11347_, _11346_, _11338_);
  nor _19681_ (_11348_, _11347_, _06427_);
  not _19682_ (_11349_, _11348_);
  not _19683_ (_11350_, _06922_);
  and _19684_ (_11351_, _11341_, _11343_);
  and _19685_ (_11353_, _06338_, _06928_);
  and _19686_ (_11354_, _11341_, _11353_);
  nor _19687_ (_11355_, _11354_, _11351_);
  nor _19688_ (_11356_, _11355_, _11350_);
  and _19689_ (_11357_, _06926_, _06362_);
  and _19690_ (_11358_, _06920_, _11339_);
  and _19691_ (_11359_, _11358_, _11357_);
  and _19692_ (_11360_, _11343_, _06920_);
  nor _19693_ (_11362_, _06924_, _06406_);
  nor _19694_ (_11363_, _06384_, _06362_);
  and _19695_ (_11365_, _11363_, _11362_);
  and _19696_ (_11366_, _11365_, _11360_);
  nor _19697_ (_11367_, _11366_, _11359_);
  not _19698_ (_11368_, _11367_);
  nor _19699_ (_11369_, _11368_, _11356_);
  and _19700_ (_11370_, _11369_, _11349_);
  nor _19701_ (_11371_, _06926_, _06916_);
  and _19702_ (_11372_, _11344_, _11339_);
  and _19703_ (_11373_, _11357_, _11372_);
  nor _19704_ (_11374_, _11373_, _11354_);
  nor _19705_ (_11376_, _11374_, _11371_);
  not _19706_ (_11377_, _06916_);
  nor _19707_ (_11378_, _11353_, _11339_);
  and _19708_ (_11379_, _11378_, _06920_);
  not _19709_ (_11380_, _11379_);
  and _19710_ (_11381_, _11380_, _11346_);
  nor _19711_ (_11382_, _11381_, _11377_);
  nor _19712_ (_11383_, _11382_, _11376_);
  and _19713_ (_11384_, _11383_, _11370_);
  not _19714_ (_11385_, _11365_);
  nor _19715_ (_11386_, _06338_, _06315_);
  and _19716_ (_11387_, _11386_, _06294_);
  nor _19717_ (_11388_, _11358_, _11387_);
  nor _19718_ (_11389_, _11388_, _11385_);
  not _19719_ (_11391_, _11389_);
  not _19720_ (_11393_, _06384_);
  and _19721_ (_11394_, _11393_, _06362_);
  and _19722_ (_11395_, _11394_, _11362_);
  and _19723_ (_11396_, _11353_, _06920_);
  and _19724_ (_11397_, _11396_, _06924_);
  nor _19725_ (_11398_, _11397_, _11395_);
  and _19726_ (_11399_, _11398_, _11391_);
  and _19727_ (_11400_, _11387_, _06928_);
  not _19728_ (_11401_, _11400_);
  nor _19729_ (_11402_, _06926_, _06915_);
  nor _19730_ (_11403_, _11402_, _11401_);
  not _19731_ (_11404_, _06927_);
  nor _19732_ (_11405_, _11360_, _06911_);
  nor _19733_ (_11406_, _11405_, _11404_);
  nor _19734_ (_11407_, _11406_, _11403_);
  and _19735_ (_11408_, _11407_, _11399_);
  not _19736_ (_11409_, _11351_);
  nor _19737_ (_11410_, _11371_, _11409_);
  not _19738_ (_11411_, _11357_);
  and _19739_ (_11412_, _11386_, _06918_);
  and _19740_ (_11414_, _11412_, _06928_);
  nor _19741_ (_11415_, _11414_, _06910_);
  nor _19742_ (_11416_, _11415_, _11411_);
  nor _19743_ (_11417_, _11416_, _11410_);
  and _19744_ (_11418_, _11417_, _11408_);
  nor _19745_ (_11419_, _11387_, _11337_);
  nor _19746_ (_11420_, _11419_, _06928_);
  nor _19747_ (_11421_, _11420_, _06929_);
  and _19748_ (_11422_, _06914_, _06406_);
  not _19749_ (_11423_, _11422_);
  nor _19750_ (_11424_, _11423_, _11421_);
  not _19751_ (_11425_, _11424_);
  nor _19752_ (_11426_, _11351_, _11396_);
  nor _19753_ (_11427_, _11426_, _11385_);
  not _19754_ (_11428_, _11427_);
  and _19755_ (_11429_, _11342_, _06927_);
  and _19756_ (_11430_, _11396_, _06916_);
  nor _19757_ (_11431_, _11430_, _11429_);
  and _19758_ (_11432_, _11431_, _11428_);
  and _19759_ (_11433_, _11432_, _11425_);
  and _19760_ (_11434_, _11433_, _11418_);
  and _19761_ (_11435_, _11378_, _06910_);
  nand _19762_ (_11436_, _11435_, _11365_);
  and _19763_ (_11437_, _11345_, _11357_);
  not _19764_ (_11438_, _11437_);
  and _19765_ (_11439_, _11438_, _11436_);
  and _19766_ (_11440_, _06910_, _06338_);
  and _19767_ (_11441_, _11440_, _06916_);
  not _19768_ (_11442_, _11441_);
  and _19769_ (_11443_, _11358_, _06927_);
  nor _19770_ (_11444_, _11342_, _11396_);
  nor _19771_ (_11445_, _11444_, _11411_);
  nor _19772_ (_11446_, _11445_, _11443_);
  and _19773_ (_11447_, _11446_, _11442_);
  and _19774_ (_11448_, _11447_, _11439_);
  and _19775_ (_11449_, _11344_, _11353_);
  nor _19776_ (_11450_, _11449_, _11360_);
  nor _19777_ (_11451_, _11450_, _11411_);
  nor _19778_ (_11452_, _11449_, _11358_);
  nor _19779_ (_11453_, _11452_, _11377_);
  nor _19780_ (_11454_, _11453_, _11451_);
  and _19781_ (_11455_, _11339_, _06910_);
  and _19782_ (_11456_, _11365_, _11455_);
  and _19783_ (_11457_, _11354_, _11365_);
  nor _19784_ (_11458_, _11457_, _11456_);
  not _19785_ (_11459_, _11458_);
  and _19786_ (_11460_, _11337_, _06928_);
  and _19787_ (_11461_, _06338_, _11340_);
  and _19788_ (_11462_, _11461_, _06918_);
  nor _19789_ (_11463_, _11462_, _11460_);
  nor _19790_ (_11464_, _11463_, _11385_);
  nor _19791_ (_11465_, _11464_, _11459_);
  and _19792_ (_11466_, _11465_, _11454_);
  and _19793_ (_11467_, _11466_, _11448_);
  and _19794_ (_11468_, _11467_, _11434_);
  and _19795_ (_11469_, _11468_, _11384_);
  nor _19796_ (_11470_, _11469_, _06255_);
  not _19797_ (_11471_, _11469_);
  and _19798_ (_11472_, _11400_, _06922_);
  not _19799_ (_11473_, _11472_);
  and _19800_ (_11474_, _06406_, _06384_);
  or _19801_ (_11475_, _11474_, _06924_);
  and _19802_ (_11476_, _11475_, _11358_);
  nor _19803_ (_11477_, _11476_, _11456_);
  and _19804_ (_11478_, _11477_, _11473_);
  and _19805_ (_11479_, _11478_, _11369_);
  and _19806_ (_11480_, _11479_, _11448_);
  nand _19807_ (_11481_, _11480_, _11471_);
  and _19808_ (_11482_, _11481_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _19809_ (_11483_, _11469_, _06255_);
  nor _19810_ (_11484_, _11483_, _11470_);
  and _19811_ (_11485_, _11484_, _11482_);
  nor _19812_ (_11486_, _11485_, _11470_);
  nor _19813_ (_11487_, _11486_, _06200_);
  and _19814_ (_11488_, _11487_, _06201_);
  nor _19815_ (_11489_, _11487_, _06201_);
  nor _19816_ (_11490_, _11489_, _11488_);
  nor _19817_ (_11491_, _11490_, _11336_);
  and _19818_ (_11492_, _06256_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _19819_ (_11493_, _11492_, _11336_);
  nor _19820_ (_11494_, _11493_, _11480_);
  or _19821_ (_11495_, _11494_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _19822_ (_11497_, _11495_, _11491_);
  and _19823_ (_10539_, _11497_, _05110_);
  not _19824_ (_11498_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  not _19825_ (_11499_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _19826_ (_11500_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _19827_ (_11501_, _11500_, _11499_);
  nor _19828_ (_11502_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor _19829_ (_11503_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _19830_ (_11504_, _11503_, _11502_);
  and _19831_ (_11505_, _11504_, _11501_);
  and _19832_ (_11506_, _11505_, _11498_);
  and _19833_ (_11507_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _19834_ (_11508_, _11507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _19835_ (_10558_, _11508_, _05110_);
  not _19836_ (_11510_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nand _19837_ (_11511_, _05474_, _11510_);
  nand _19838_ (_11512_, _11511_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _19839_ (_11513_, _11512_, _11506_);
  and _19840_ (_10562_, _11513_, _05110_);
  and _19841_ (_10567_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _05110_);
  not _19842_ (_11515_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _19843_ (_11516_, _06880_, _11515_);
  or _19844_ (_11517_, _11516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _19845_ (_11518_, _11517_, _11326_);
  not _19846_ (_11519_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _19847_ (_11520_, _05488_, _11519_);
  nand _19848_ (_11521_, _11520_, _11326_);
  or _19849_ (_11523_, _11521_, _05784_);
  and _19850_ (_11524_, _11523_, _11518_);
  or _19851_ (_11525_, _11524_, _11329_);
  nand _19852_ (_11526_, _11329_, _05841_);
  and _19853_ (_11527_, _11526_, _05110_);
  and _19854_ (_10582_, _11527_, _11525_);
  and _19855_ (_11528_, _11326_, _08133_);
  nand _19856_ (_11529_, _11528_, _05872_);
  or _19857_ (_11530_, _11528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _19858_ (_11532_, _11530_, _11330_);
  and _19859_ (_11533_, _11532_, _11529_);
  nor _19860_ (_11535_, _11330_, _06054_);
  or _19861_ (_11536_, _11535_, _11533_);
  and _19862_ (_10585_, _11536_, _05110_);
  and _19863_ (_11537_, _10178_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _19864_ (_11538_, _11537_, _10209_);
  and _19865_ (_11539_, _11538_, _11326_);
  not _19866_ (_11540_, _11326_);
  or _19867_ (_11541_, _11540_, _10212_);
  and _19868_ (_11542_, _11541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or _19869_ (_11543_, _11542_, _11329_);
  or _19870_ (_11544_, _11543_, _11539_);
  nand _19871_ (_11545_, _11329_, _05334_);
  and _19872_ (_11546_, _11545_, _05110_);
  and _19873_ (_10587_, _11546_, _11544_);
  and _19874_ (_11547_, _11326_, _06632_);
  not _19875_ (_11548_, _05866_);
  nand _19876_ (_11549_, _11326_, _05401_);
  or _19877_ (_11550_, _11549_, _11548_);
  and _19878_ (_11551_, _11550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _19879_ (_11552_, _11551_, _11329_);
  or _19880_ (_11553_, _11552_, _11547_);
  nand _19881_ (_11554_, _11329_, _06088_);
  and _19882_ (_11555_, _11554_, _05110_);
  and _19883_ (_10597_, _11555_, _11553_);
  and _19884_ (_11556_, _06173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _19885_ (_11557_, _11556_, _08245_);
  and _19886_ (_11558_, _11557_, _11326_);
  not _19887_ (_11559_, _10169_);
  nand _19888_ (_11560_, _11326_, _11559_);
  and _19889_ (_11561_, _11560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _19890_ (_11562_, _11561_, _11329_);
  or _19891_ (_11563_, _11562_, _11558_);
  nand _19892_ (_11564_, _11329_, _06229_);
  and _19893_ (_11565_, _11564_, _05110_);
  and _19894_ (_10600_, _11565_, _11563_);
  not _19895_ (_11566_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _19896_ (_11567_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor _19897_ (_11568_, _11567_, _11566_);
  and _19898_ (_11569_, _11567_, _11566_);
  nor _19899_ (_11570_, _11569_, _11568_);
  not _19900_ (_11571_, _11570_);
  and _19901_ (_11572_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _19902_ (_11573_, _11572_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _19903_ (_11574_, _11572_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _19904_ (_11575_, _11574_, _11573_);
  or _19905_ (_11576_, _11575_, _11567_);
  and _19906_ (_11577_, _11576_, _11571_);
  nor _19907_ (_11578_, _11568_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _19908_ (_11579_, _11568_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _19909_ (_11580_, _11579_, _11578_);
  or _19910_ (_11581_, _11573_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _19911_ (_03099_, _11581_, _05110_);
  and _19912_ (_11582_, _03099_, _11580_);
  and _19913_ (_10620_, _11582_, _11577_);
  and _19914_ (_10641_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _05110_);
  nor _19915_ (_11583_, _11240_, _06229_);
  nor _19916_ (_11584_, _11239_, _11234_);
  and _19917_ (_11585_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _19918_ (_11586_, _11585_, _11202_);
  and _19919_ (_11587_, _11586_, _11223_);
  nand _19920_ (_11588_, _11218_, _11202_);
  nor _19921_ (_11589_, _11588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _19922_ (_11590_, _11588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _19923_ (_11591_, _11590_, _11193_);
  or _19924_ (_11592_, _11591_, _11589_);
  or _19925_ (_11593_, _11592_, _11587_);
  or _19926_ (_11594_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _19927_ (_11595_, _11594_, _11593_);
  and _19928_ (_11596_, _11595_, _11584_);
  and _19929_ (_11597_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _19930_ (_11598_, _11597_, _11596_);
  or _19931_ (_11599_, _11598_, _11583_);
  and _19932_ (_10645_, _11599_, _05110_);
  not _19933_ (_11600_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _19934_ (_11601_, _11216_, _11202_);
  nor _19935_ (_11602_, _11601_, _11600_);
  or _19936_ (_11603_, _11602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _19937_ (_11604_, _11603_, _11588_);
  or _19938_ (_11605_, _11604_, _11193_);
  and _19939_ (_11606_, _11202_, _11225_);
  and _19940_ (_11607_, _11606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _19941_ (_11608_, _11607_, _11223_);
  or _19942_ (_11609_, _11608_, _11605_);
  or _19943_ (_11610_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _19944_ (_11611_, _11610_, _11609_);
  and _19945_ (_11612_, _11611_, _11584_);
  nor _19946_ (_11613_, _11240_, _05938_);
  and _19947_ (_11614_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _19948_ (_11615_, _11614_, _11613_);
  or _19949_ (_11616_, _11615_, _11612_);
  and _19950_ (_10649_, _11616_, _05110_);
  and _19951_ (_11617_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _07601_);
  and _19952_ (_11618_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _19953_ (_11619_, _11618_, _11617_);
  and _19954_ (_10654_, _11619_, _05110_);
  and _19955_ (_11620_, _11239_, _06799_);
  and _19956_ (_11621_, _11601_, _11600_);
  nor _19957_ (_11622_, _11621_, _11602_);
  or _19958_ (_11623_, _11622_, _11193_);
  and _19959_ (_11625_, _11606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _19960_ (_11626_, _11625_, _11223_);
  or _19961_ (_11627_, _11626_, _11623_);
  not _19962_ (_11628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand _19963_ (_11629_, _11193_, _11628_);
  and _19964_ (_11630_, _11629_, _11627_);
  and _19965_ (_11631_, _11630_, _11584_);
  and _19966_ (_11632_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _19967_ (_11633_, _11632_, _11631_);
  or _19968_ (_11634_, _11633_, _11620_);
  and _19969_ (_10660_, _11634_, _05110_);
  and _19970_ (_11635_, _06380_, _06311_);
  and _19971_ (_11636_, _11635_, _06423_);
  and _19972_ (_11637_, _11325_, _05475_);
  and _19973_ (_11638_, _11637_, _06266_);
  and _19974_ (_11639_, _06334_, _06289_);
  and _19975_ (_11640_, _11639_, _11638_);
  and _19976_ (_11641_, _06402_, _06357_);
  and _19977_ (_11642_, _11641_, _11640_);
  and _19978_ (_10663_, _11642_, _11636_);
  and _19979_ (_11644_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _19980_ (_11645_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _19981_ (_11646_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _19982_ (_11647_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _19983_ (_11648_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _19984_ (_11650_, _11648_, _11646_);
  and _19985_ (_11651_, _11650_, _11647_);
  nor _19986_ (_11652_, _11651_, _11646_);
  nor _19987_ (_11653_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _19988_ (_11654_, _11653_, _11645_);
  not _19989_ (_11655_, _11654_);
  nor _19990_ (_11656_, _11655_, _11652_);
  nor _19991_ (_11657_, _11656_, _11645_);
  not _19992_ (_11658_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _19993_ (_11660_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _19994_ (_11661_, _11660_, _11658_);
  and _19995_ (_11662_, _11661_, _11657_);
  and _19996_ (_11664_, _11657_, _11660_);
  nor _19997_ (_11665_, _11664_, _11658_);
  nor _19998_ (_11666_, _11665_, _11662_);
  not _19999_ (_11667_, _11666_);
  not _20000_ (_11669_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _20001_ (_11670_, _11657_, _11669_);
  nor _20002_ (_11671_, _11657_, _11669_);
  nor _20003_ (_11672_, _11671_, _11670_);
  not _20004_ (_11673_, _11672_);
  nor _20005_ (_11675_, _11650_, _11647_);
  nor _20006_ (_11676_, _11675_, _11651_);
  nand _20007_ (_11677_, _11676_, _11471_);
  not _20008_ (_11678_, _11677_);
  nor _20009_ (_11680_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _20010_ (_11681_, _11680_, _11647_);
  and _20011_ (_11682_, _11681_, _11481_);
  or _20012_ (_11683_, _11676_, _11471_);
  and _20013_ (_11684_, _11683_, _11677_);
  and _20014_ (_11685_, _11684_, _11682_);
  or _20015_ (_11686_, _11685_, _11678_);
  and _20016_ (_11687_, _11655_, _11652_);
  nor _20017_ (_11688_, _11687_, _11656_);
  and _20018_ (_11689_, _11688_, _11686_);
  and _20019_ (_11690_, _11689_, _11673_);
  not _20020_ (_11691_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _20021_ (_11692_, _11670_, _11691_);
  or _20022_ (_11693_, _11692_, _11664_);
  and _20023_ (_11695_, _11693_, _11690_);
  and _20024_ (_11696_, _11695_, _11667_);
  nor _20025_ (_11698_, _11695_, _11667_);
  nor _20026_ (_11699_, _11698_, _11696_);
  or _20027_ (_11700_, _11699_, _07437_);
  or _20028_ (_11701_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _20029_ (_11703_, _11701_, _11510_);
  and _20030_ (_11705_, _11703_, _11700_);
  or _20031_ (_11706_, _11705_, _11644_);
  and _20032_ (_10679_, _11706_, _05110_);
  and _20033_ (_11708_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _20034_ (_11709_, _11708_, _11202_);
  and _20035_ (_11710_, _11709_, _11223_);
  and _20036_ (_11711_, _11220_, _11202_);
  and _20037_ (_11712_, _11711_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _20038_ (_11713_, _11711_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _20039_ (_11714_, _11713_, _11712_);
  or _20040_ (_11715_, _11714_, _11193_);
  or _20041_ (_11716_, _11715_, _11710_);
  nor _20042_ (_11717_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor _20043_ (_11719_, _11717_, _11234_);
  and _20044_ (_11720_, _11719_, _11716_);
  and _20045_ (_11721_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _20046_ (_11722_, _11721_, _11239_);
  or _20047_ (_11723_, _11722_, _11720_);
  nand _20048_ (_11724_, _11239_, _05334_);
  and _20049_ (_11726_, _11724_, _05110_);
  and _20050_ (_10684_, _11726_, _11723_);
  and _20051_ (_11727_, _06824_, _06813_);
  and _20052_ (_11728_, _11727_, _06451_);
  and _20053_ (_11729_, _07038_, _06277_);
  and _20054_ (_11730_, _11729_, _06451_);
  nor _20055_ (_11731_, _11730_, _07147_);
  not _20056_ (_11732_, _11731_);
  nor _20057_ (_11734_, _11732_, _11728_);
  nor _20058_ (_11735_, _11734_, _06239_);
  not _20059_ (_11736_, _11314_);
  and _20060_ (_11737_, _07077_, _06277_);
  or _20061_ (_11738_, _11737_, _07088_);
  or _20062_ (_11740_, _11738_, _07122_);
  nand _20063_ (_11741_, _07115_, _06276_);
  and _20064_ (_11742_, _07077_, _06276_);
  nor _20065_ (_11743_, _11742_, _07081_);
  nand _20066_ (_11744_, _11743_, _11741_);
  or _20067_ (_11745_, _11744_, _07086_);
  nor _20068_ (_11746_, _11745_, _11740_);
  not _20069_ (_11747_, _07076_);
  nand _20070_ (_11748_, _06825_, _06810_);
  and _20071_ (_11749_, _06856_, _06810_);
  nor _20072_ (_11750_, _11749_, _11301_);
  and _20073_ (_11751_, _11750_, _11748_);
  and _20074_ (_11752_, _11751_, _11747_);
  and _20075_ (_11753_, _11752_, _11734_);
  and _20076_ (_11754_, _06864_, _06438_);
  or _20077_ (_11755_, _11754_, _07139_);
  and _20078_ (_11756_, _11292_, _06810_);
  nor _20079_ (_11757_, _11756_, _11755_);
  or _20080_ (_11758_, _07069_, _06463_);
  nand _20081_ (_11759_, _11758_, _06810_);
  not _20082_ (_11760_, _11759_);
  and _20083_ (_11761_, _06941_, _06277_);
  nor _20084_ (_11762_, _11761_, _11760_);
  and _20085_ (_11763_, _11762_, _11757_);
  nor _20086_ (_11764_, _07116_, _07051_);
  nor _20087_ (_11765_, _07132_, _07127_);
  and _20088_ (_11766_, _11765_, _11764_);
  nor _20089_ (_11767_, _06845_, _06817_);
  and _20090_ (_11768_, _11767_, _07110_);
  and _20091_ (_11769_, _11768_, _11766_);
  and _20092_ (_11770_, _11769_, _11763_);
  and _20093_ (_11771_, _11770_, _11753_);
  nand _20094_ (_11772_, _11771_, _11746_);
  nand _20095_ (_11773_, _11772_, _06870_);
  nor _20096_ (_11774_, _11309_, _11284_);
  nand _20097_ (_11775_, _11774_, _11773_);
  nand _20098_ (_11776_, _11775_, _05151_);
  and _20099_ (_11777_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _20100_ (_11778_, _11777_);
  and _20101_ (_11779_, _11778_, _11776_);
  and _20102_ (_11780_, _11779_, _11736_);
  and _20103_ (_11781_, _11780_, _11323_);
  nor _20104_ (_11782_, _10176_, _10215_);
  nor _20105_ (_11783_, _11782_, _10220_);
  or _20106_ (_11784_, _11783_, _05419_);
  nand _20107_ (_11785_, _11783_, _05419_);
  and _20108_ (_11786_, _11785_, _11784_);
  nor _20109_ (_11787_, _10180_, _10177_);
  nand _20110_ (_11788_, _11787_, _05390_);
  and _20111_ (_11789_, _05433_, _05337_);
  and _20112_ (_11790_, _11789_, _06173_);
  and _20113_ (_11791_, _11790_, _05461_);
  and _20114_ (_11792_, _11791_, _11788_);
  or _20115_ (_11793_, _11787_, _05390_);
  nor _20116_ (_11794_, _06366_, _05375_);
  and _20117_ (_11795_, _06366_, _05375_);
  nor _20118_ (_11796_, _11795_, _11794_);
  and _20119_ (_11797_, _11796_, _11793_);
  and _20120_ (_11798_, _11797_, _11792_);
  and _20121_ (_11799_, _11798_, _11786_);
  and _20122_ (_11800_, _11799_, _06088_);
  not _20123_ (_11801_, _11783_);
  not _20124_ (_11802_, _06366_);
  and _20125_ (_11803_, _11787_, _11802_);
  and _20126_ (_11804_, _11803_, _11801_);
  nand _20127_ (_11805_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor _20128_ (_11806_, _11787_, _06366_);
  and _20129_ (_11807_, _11806_, _11783_);
  nand _20130_ (_11808_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _20131_ (_11809_, _11808_, _11805_);
  nor _20132_ (_11810_, _11787_, _11802_);
  and _20133_ (_11811_, _11810_, _11801_);
  nand _20134_ (_11812_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and _20135_ (_11813_, _11787_, _06366_);
  and _20136_ (_11814_, _11813_, _11783_);
  nand _20137_ (_11815_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _20138_ (_11816_, _11815_, _11812_);
  and _20139_ (_11817_, _11816_, _11809_);
  not _20140_ (_11818_, _11799_);
  and _20141_ (_11819_, _11813_, _11801_);
  nand _20142_ (_11820_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and _20143_ (_11821_, _11803_, _11783_);
  nand _20144_ (_11822_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _20145_ (_11823_, _11822_, _11820_);
  and _20146_ (_11824_, _11806_, _11801_);
  nand _20147_ (_11825_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _20148_ (_11826_, _11810_, _11783_);
  nand _20149_ (_11827_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _20150_ (_11828_, _11827_, _11825_);
  and _20151_ (_11829_, _11828_, _11823_);
  and _20152_ (_11830_, _11829_, _11818_);
  and _20153_ (_11831_, _11830_, _11817_);
  nor _20154_ (_11832_, _11831_, _11800_);
  nand _20155_ (_11833_, _11832_, _11781_);
  nand _20156_ (_11834_, _11778_, _11776_);
  and _20157_ (_11835_, _11323_, _11314_);
  nand _20158_ (_11836_, _11835_, _11834_);
  or _20159_ (_11837_, _11836_, _07470_);
  and _20160_ (_11838_, _11837_, _11833_);
  and _20161_ (_11839_, _11834_, _11736_);
  nand _20162_ (_11840_, _11839_, _11323_);
  nand _20163_ (_11841_, _07206_, _08272_);
  or _20164_ (_11842_, _11841_, _06088_);
  and _20165_ (_11843_, _07206_, _08272_);
  nand _20166_ (_11844_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _20167_ (_11845_, _11844_, _11842_);
  nand _20168_ (_11846_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  or _20169_ (_11847_, _11841_, _06229_);
  and _20170_ (_11848_, _11847_, _11846_);
  nand _20171_ (_11849_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  or _20172_ (_11850_, _11841_, _05938_);
  and _20173_ (_11851_, _11850_, _11849_);
  not _20174_ (_11852_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  or _20175_ (_11853_, _11843_, _05369_);
  or _20176_ (_11854_, _11841_, _06798_);
  nand _20177_ (_11855_, _11854_, _11853_);
  nor _20178_ (_11856_, _11855_, _11852_);
  and _20179_ (_11857_, _11856_, _11851_);
  and _20180_ (_11858_, _11857_, _11848_);
  and _20181_ (_11859_, _11858_, _11845_);
  or _20182_ (_11860_, _11858_, _11845_);
  not _20183_ (_11861_, _11860_);
  nor _20184_ (_11862_, _11861_, _11859_);
  or _20185_ (_11863_, _11862_, _05341_);
  and _20186_ (_11864_, _11863_, _05384_);
  or _20187_ (_11865_, _11864_, _11843_);
  and _20188_ (_11866_, _11865_, _11842_);
  or _20189_ (_11867_, _11866_, _11840_);
  nand _20190_ (_11868_, _11835_, _11779_);
  or _20191_ (_11869_, _11868_, _11787_);
  and _20192_ (_11870_, _11869_, _11867_);
  and _20193_ (_11871_, _11870_, _11838_);
  or _20194_ (_11872_, _11871_, _05390_);
  nand _20195_ (_11873_, _11870_, _11838_);
  or _20196_ (_11874_, _11873_, _05389_);
  and _20197_ (_11875_, _11874_, _11872_);
  and _20198_ (_11876_, _11839_, _11323_);
  nor _20199_ (_11877_, _11841_, _06054_);
  or _20200_ (_11878_, _11841_, _05334_);
  nand _20201_ (_11879_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _20202_ (_11880_, _11879_, _11878_);
  and _20203_ (_11881_, _11880_, _11859_);
  and _20204_ (_11882_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _20205_ (_11883_, _11882_, _11877_);
  and _20206_ (_11884_, _11883_, _11881_);
  nor _20207_ (_11885_, _11883_, _11881_);
  or _20208_ (_11886_, _11885_, _11884_);
  nand _20209_ (_11887_, _11886_, _05790_);
  nand _20210_ (_11888_, _11887_, _05423_);
  and _20211_ (_11889_, _11888_, _11841_);
  or _20212_ (_11890_, _11889_, _11877_);
  nand _20213_ (_11891_, _11890_, _11876_);
  nand _20214_ (_11892_, _11799_, _06054_);
  nand _20215_ (_11893_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nand _20216_ (_11894_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _20217_ (_11895_, _11894_, _11893_);
  nand _20218_ (_11896_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nand _20219_ (_11897_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _20220_ (_11898_, _11897_, _11896_);
  and _20221_ (_11899_, _11898_, _11895_);
  nand _20222_ (_11900_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nand _20223_ (_11901_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _20224_ (_11902_, _11901_, _11900_);
  nand _20225_ (_11903_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nand _20226_ (_11904_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and _20227_ (_11905_, _11904_, _11903_);
  and _20228_ (_11906_, _11905_, _11902_);
  and _20229_ (_11907_, _11906_, _11818_);
  nand _20230_ (_11908_, _11907_, _11899_);
  and _20231_ (_11909_, _11908_, _11892_);
  nand _20232_ (_11910_, _11909_, _11781_);
  or _20233_ (_11911_, _11836_, _07507_);
  and _20234_ (_11912_, _11911_, _11910_);
  or _20235_ (_11914_, _11779_, _11736_);
  nor _20236_ (_11915_, _11780_, _11323_);
  nand _20237_ (_11916_, _11915_, _11914_);
  and _20238_ (_11917_, _11916_, _11912_);
  and _20239_ (_11918_, _11917_, _11891_);
  and _20240_ (_11919_, _11918_, _06121_);
  nand _20241_ (_11920_, _11917_, _11891_);
  and _20242_ (_11921_, _11920_, _05433_);
  nor _20243_ (_11922_, _11921_, _11919_);
  or _20244_ (_11923_, _11868_, _11783_);
  or _20245_ (_11924_, _11836_, _07490_);
  and _20246_ (_11925_, _11924_, _11923_);
  and _20247_ (_11926_, _11799_, _05334_);
  and _20248_ (_11927_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _20249_ (_11928_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _20250_ (_11929_, _11928_, _11927_);
  and _20251_ (_11930_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and _20252_ (_11931_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _20253_ (_11932_, _11931_, _11930_);
  and _20254_ (_11933_, _11932_, _11929_);
  nand _20255_ (_11934_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nand _20256_ (_11935_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _20257_ (_11936_, _11935_, _11934_);
  nand _20258_ (_11937_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nand _20259_ (_11938_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _20260_ (_11939_, _11938_, _11937_);
  and _20261_ (_11941_, _11939_, _11936_);
  and _20262_ (_11942_, _11941_, _11818_);
  and _20263_ (_11943_, _11942_, _11933_);
  nor _20264_ (_11944_, _11943_, _11926_);
  nand _20265_ (_11945_, _11944_, _11781_);
  not _20266_ (_11946_, _11323_);
  and _20267_ (_11948_, _11946_, _11314_);
  nor _20268_ (_11949_, _11880_, _11859_);
  or _20269_ (_11950_, _11949_, _11881_);
  nand _20270_ (_11951_, _11950_, _05790_);
  nand _20271_ (_11952_, _11951_, _05408_);
  nand _20272_ (_11953_, _11952_, _11841_);
  nand _20273_ (_11954_, _11953_, _11878_);
  and _20274_ (_11955_, _11954_, _11876_);
  nor _20275_ (_11956_, _11955_, _11948_);
  and _20276_ (_11957_, _11956_, _11945_);
  nand _20277_ (_11958_, _11957_, _11925_);
  or _20278_ (_11959_, _11958_, _05418_);
  and _20279_ (_11960_, _11957_, _11925_);
  or _20280_ (_11961_, _11960_, _05419_);
  and _20281_ (_11962_, _11961_, _11959_);
  and _20282_ (_11963_, _11843_, _05901_);
  nor _20283_ (_11964_, _11841_, _05841_);
  and _20284_ (_11965_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _20285_ (_11966_, _11965_, _11964_);
  nand _20286_ (_11967_, _11966_, _11884_);
  not _20287_ (_11968_, _11967_);
  and _20288_ (_11969_, _11841_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand _20289_ (_11970_, _11969_, _11968_);
  or _20290_ (_11971_, _11969_, _11968_);
  and _20291_ (_11972_, _11971_, _05790_);
  nand _20292_ (_11973_, _11972_, _11970_);
  and _20293_ (_11974_, _11841_, _05452_);
  and _20294_ (_11975_, _11974_, _11973_);
  nor _20295_ (_11976_, _11975_, _11963_);
  nand _20296_ (_11977_, _11976_, _11839_);
  nand _20297_ (_11978_, _11799_, _05901_);
  nand _20298_ (_11979_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand _20299_ (_11981_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _20300_ (_11982_, _11981_, _11979_);
  nand _20301_ (_11984_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nand _20302_ (_11985_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _20303_ (_11986_, _11985_, _11984_);
  and _20304_ (_11987_, _11986_, _11982_);
  nand _20305_ (_11988_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand _20306_ (_11989_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _20307_ (_11990_, _11989_, _11988_);
  nand _20308_ (_11992_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nand _20309_ (_11993_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _20310_ (_11994_, _11993_, _11992_);
  and _20311_ (_11995_, _11994_, _11990_);
  and _20312_ (_11996_, _11995_, _11818_);
  nand _20313_ (_11997_, _11996_, _11987_);
  and _20314_ (_11998_, _11997_, _11978_);
  nand _20315_ (_11999_, _11998_, _11781_);
  nor _20316_ (_12000_, _05474_, _05454_);
  and _20317_ (_12001_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  not _20318_ (_12002_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _20319_ (_12003_, _06251_, _12002_);
  nor _20320_ (_12004_, _12003_, _12001_);
  and _20321_ (_12005_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _20322_ (_12006_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _20323_ (_12007_, _12006_, _12005_);
  and _20324_ (_12008_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _20325_ (_12009_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _20326_ (_12010_, _12009_, _12008_);
  and _20327_ (_12011_, _12010_, _12007_);
  and _20328_ (_12012_, _12011_, _12004_);
  nor _20329_ (_12013_, _12012_, _07437_);
  nor _20330_ (_12014_, _12013_, _12000_);
  or _20331_ (_12016_, _12014_, _11914_);
  and _20332_ (_12017_, _12016_, _11323_);
  and _20333_ (_12018_, _12017_, _11999_);
  and _20334_ (_12020_, _12018_, _11977_);
  and _20335_ (_12021_, _12020_, _05460_);
  nor _20336_ (_12022_, _12020_, _05460_);
  nor _20337_ (_12023_, _12022_, _12021_);
  or _20338_ (_12024_, _11966_, _11884_);
  nand _20339_ (_12025_, _12024_, _11967_);
  nand _20340_ (_12026_, _12025_, _05790_);
  nand _20341_ (_12027_, _12026_, _05439_);
  and _20342_ (_12028_, _12027_, _11841_);
  or _20343_ (_12029_, _12028_, _11964_);
  nand _20344_ (_12030_, _12029_, _11876_);
  nand _20345_ (_12031_, _11799_, _05841_);
  nand _20346_ (_12032_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nand _20347_ (_12033_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _20348_ (_12034_, _12033_, _12032_);
  nand _20349_ (_12035_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nand _20350_ (_12036_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _20351_ (_12037_, _12036_, _12035_);
  and _20352_ (_12038_, _12037_, _12034_);
  nand _20353_ (_12039_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nand _20354_ (_12040_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _20355_ (_12041_, _12040_, _12039_);
  nand _20356_ (_12042_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nand _20357_ (_12043_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _20358_ (_12044_, _12043_, _12042_);
  and _20359_ (_12045_, _12044_, _12041_);
  and _20360_ (_12046_, _12045_, _11818_);
  nand _20361_ (_12048_, _12046_, _12038_);
  and _20362_ (_12049_, _12048_, _12031_);
  nand _20363_ (_12050_, _12049_, _11781_);
  and _20364_ (_12051_, _12050_, _12030_);
  nor _20365_ (_12052_, _05474_, _05441_);
  and _20366_ (_12053_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  not _20367_ (_12054_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _20368_ (_12056_, _06251_, _12054_);
  nor _20369_ (_12057_, _12056_, _12053_);
  and _20370_ (_12058_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _20371_ (_12059_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _20372_ (_12060_, _12059_, _12058_);
  and _20373_ (_12061_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _20374_ (_12062_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _20375_ (_12063_, _12062_, _12061_);
  and _20376_ (_12064_, _12063_, _12060_);
  and _20377_ (_12065_, _12064_, _12057_);
  nor _20378_ (_12066_, _12065_, _07437_);
  nor _20379_ (_12067_, _12066_, _12052_);
  nor _20380_ (_12068_, _12067_, _11836_);
  nor _20381_ (_12070_, _11915_, _12068_);
  nand _20382_ (_12071_, _12070_, _12051_);
  or _20383_ (_12072_, _12071_, _05447_);
  and _20384_ (_12073_, _12070_, _12051_);
  or _20385_ (_12074_, _12073_, _05448_);
  and _20386_ (_12075_, _12074_, _12072_);
  and _20387_ (_12077_, _12075_, _12023_);
  and _20388_ (_12078_, _12077_, _11962_);
  and _20389_ (_12080_, _12078_, _11922_);
  and _20390_ (_12082_, _12080_, _11875_);
  not _20391_ (_12083_, _05867_);
  and _20392_ (_12084_, _12083_, _05806_);
  and _20393_ (_12086_, _12084_, _12082_);
  and _20394_ (_12087_, _12086_, _11735_);
  not _20395_ (_12088_, _12087_);
  not _20396_ (_12089_, _06870_);
  nor _20397_ (_12090_, _07105_, _06866_);
  nor _20398_ (_12091_, _12090_, _12089_);
  not _20399_ (_12092_, _06997_);
  not _20400_ (_12093_, _11284_);
  not _20401_ (_12094_, _06873_);
  or _20402_ (_12095_, _11728_, _07147_);
  nor _20403_ (_12096_, _12095_, _11730_);
  nor _20404_ (_12097_, _12096_, _12094_);
  nor _20405_ (_12098_, _12096_, _12089_);
  nor _20406_ (_12099_, _12098_, _12097_);
  and _20407_ (_12100_, _12099_, _12093_);
  and _20408_ (_12101_, _07396_, _05696_);
  and _20409_ (_12102_, _07309_, _06640_);
  nand _20410_ (_12103_, _12102_, _12101_);
  nor _20411_ (_12104_, _12103_, _07211_);
  and _20412_ (_12105_, _12104_, _06516_);
  and _20413_ (_12106_, _12105_, _12100_);
  and _20414_ (_12108_, _12106_, _06759_);
  and _20415_ (_12109_, _12108_, _12092_);
  nor _20416_ (_12111_, _11735_, _06436_);
  nor _20417_ (_12112_, _12111_, _12093_);
  and _20418_ (_12114_, _12112_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _20419_ (_12115_, _11735_, _05185_);
  nor _20420_ (_12117_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _20421_ (_12118_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _20422_ (_12119_, _12118_, _12117_);
  nor _20423_ (_12120_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _20424_ (_12121_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _20425_ (_12123_, _12121_, _12120_);
  and _20426_ (_12125_, _12123_, _12119_);
  and _20427_ (_12126_, _12125_, _11286_);
  or _20428_ (_12127_, _12126_, _12115_);
  or _20429_ (_12128_, _12127_, _12114_);
  nor _20430_ (_12130_, _12128_, _12109_);
  and _20431_ (_12131_, _06811_, _06431_);
  not _20432_ (_12132_, _12131_);
  and _20433_ (_12134_, _06825_, _06464_);
  nor _20434_ (_12135_, _12134_, _06812_);
  and _20435_ (_12137_, _12135_, _12132_);
  and _20436_ (_12138_, _07138_, _06451_);
  and _20437_ (_12140_, _07087_, _06451_);
  or _20438_ (_12141_, _12140_, _11728_);
  or _20439_ (_12142_, _12141_, _12138_);
  nor _20440_ (_12144_, _12142_, _06828_);
  and _20441_ (_12145_, _12144_, _12137_);
  not _20442_ (_12146_, _12145_);
  and _20443_ (_12147_, _12146_, _12130_);
  not _20444_ (_12148_, _12147_);
  not _20445_ (_12149_, _07073_);
  and _20446_ (_12150_, _12149_, _06451_);
  nor _20447_ (_12151_, _12150_, _11732_);
  nor _20448_ (_12153_, _12151_, _12130_);
  not _20449_ (_12154_, _11301_);
  and _20450_ (_12156_, _07087_, _06448_);
  and _20451_ (_12158_, _06451_, _06438_);
  nor _20452_ (_12159_, _12158_, _12156_);
  and _20453_ (_12160_, _12159_, _12154_);
  not _20454_ (_12162_, _12160_);
  nor _20455_ (_12163_, _12162_, _12153_);
  and _20456_ (_12165_, _12163_, _12148_);
  nor _20457_ (_12166_, _11309_, _06873_);
  nor _20458_ (_12168_, _12166_, _12165_);
  nor _20459_ (_12169_, _12168_, _12091_);
  nor _20460_ (_12171_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _20461_ (_12172_, _12171_);
  nor _20462_ (_12173_, _12172_, _10176_);
  and _20463_ (_12175_, _12173_, _10211_);
  not _20464_ (_12176_, _12175_);
  and _20465_ (_12177_, _12176_, _12112_);
  not _20466_ (_12178_, _06628_);
  and _20467_ (_12179_, _06638_, _12178_);
  not _20468_ (_12180_, _12179_);
  and _20469_ (_12181_, _12180_, _11286_);
  nor _20470_ (_12182_, _12181_, _12177_);
  not _20471_ (_12183_, _12182_);
  nor _20472_ (_12184_, _12183_, _12169_);
  and _20473_ (_12185_, _11780_, _11946_);
  nor _20474_ (_12186_, _11856_, _11851_);
  nor _20475_ (_12187_, _12186_, _11857_);
  nor _20476_ (_12188_, _12187_, _05341_);
  nor _20477_ (_12189_, _12188_, _05346_);
  nor _20478_ (_12190_, _12189_, _11843_);
  not _20479_ (_12192_, _12190_);
  and _20480_ (_12193_, _12192_, _11850_);
  not _20481_ (_12194_, _12193_);
  and _20482_ (_12195_, _12194_, _11876_);
  nor _20483_ (_12197_, _12195_, _12185_);
  or _20484_ (_12198_, _11836_, _07439_);
  nand _20485_ (_12200_, _11799_, _05938_);
  nand _20486_ (_12201_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nand _20487_ (_12203_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and _20488_ (_12204_, _12203_, _12201_);
  nand _20489_ (_12205_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nand _20490_ (_12207_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _20491_ (_12208_, _12207_, _12205_);
  and _20492_ (_12209_, _12208_, _12204_);
  nand _20493_ (_12210_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nand _20494_ (_12211_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _20495_ (_12212_, _12211_, _12210_);
  nand _20496_ (_12213_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nand _20497_ (_12214_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _20498_ (_12215_, _12214_, _12213_);
  and _20499_ (_12216_, _12215_, _12212_);
  and _20500_ (_12217_, _12216_, _11818_);
  nand _20501_ (_12219_, _12217_, _12209_);
  and _20502_ (_12220_, _12219_, _12200_);
  nand _20503_ (_12221_, _12220_, _11781_);
  or _20504_ (_12222_, _11868_, _06445_);
  and _20505_ (_12223_, _12222_, _12221_);
  and _20506_ (_12224_, _12223_, _12198_);
  and _20507_ (_12225_, _12224_, _12197_);
  or _20508_ (_12227_, _12225_, _05365_);
  nand _20509_ (_12228_, _12224_, _12197_);
  or _20510_ (_12229_, _12228_, _05486_);
  nand _20511_ (_12230_, _12229_, _12227_);
  nand _20512_ (_12231_, _11799_, _06229_);
  nand _20513_ (_12232_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nand _20514_ (_12233_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _20515_ (_12234_, _12233_, _12232_);
  nand _20516_ (_12235_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nand _20517_ (_12236_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _20518_ (_12237_, _12236_, _12235_);
  and _20519_ (_12239_, _12237_, _12234_);
  nand _20520_ (_12240_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nand _20521_ (_12241_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _20522_ (_12242_, _12241_, _12240_);
  nand _20523_ (_12243_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nand _20524_ (_12245_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _20525_ (_12246_, _12245_, _12243_);
  and _20526_ (_12248_, _12246_, _12242_);
  and _20527_ (_12249_, _12248_, _11818_);
  nand _20528_ (_12250_, _12249_, _12239_);
  and _20529_ (_12252_, _12250_, _12231_);
  nand _20530_ (_12253_, _12252_, _11781_);
  or _20531_ (_12254_, _11836_, _07454_);
  and _20532_ (_12255_, _12254_, _12253_);
  nor _20533_ (_12256_, _11857_, _11848_);
  or _20534_ (_12257_, _12256_, _11858_);
  and _20535_ (_12258_, _12257_, _05790_);
  or _20536_ (_12259_, _12258_, _05393_);
  nand _20537_ (_12260_, _12259_, _11841_);
  nand _20538_ (_12262_, _12260_, _11847_);
  nand _20539_ (_12263_, _12262_, _11876_);
  not _20540_ (_12264_, _06411_);
  or _20541_ (_12265_, _11868_, _12264_);
  and _20542_ (_12266_, _12265_, _12263_);
  and _20543_ (_12268_, _12266_, _12255_);
  or _20544_ (_12269_, _12268_, _05401_);
  nand _20545_ (_12270_, _12266_, _12255_);
  or _20546_ (_12272_, _12270_, _05485_);
  nand _20547_ (_12273_, _12272_, _12269_);
  and _20548_ (_12274_, _11799_, _06798_);
  nand _20549_ (_12275_, _11826_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nand _20550_ (_12276_, _11807_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _20551_ (_12277_, _12276_, _12275_);
  nand _20552_ (_12278_, _11819_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nand _20553_ (_12279_, _11814_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _20554_ (_12280_, _12279_, _12278_);
  and _20555_ (_12281_, _12280_, _12277_);
  nand _20556_ (_12282_, _11811_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nand _20557_ (_12283_, _11804_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _20558_ (_12284_, _12283_, _12282_);
  nand _20559_ (_12285_, _11824_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nand _20560_ (_12286_, _11821_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _20561_ (_12287_, _12286_, _12285_);
  and _20562_ (_12288_, _12287_, _12284_);
  and _20563_ (_12289_, _12288_, _11818_);
  and _20564_ (_12290_, _12289_, _12281_);
  nor _20565_ (_12291_, _12290_, _12274_);
  nand _20566_ (_12292_, _12291_, _11781_);
  nor _20567_ (_12294_, _05474_, _05234_);
  and _20568_ (_12295_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  not _20569_ (_12297_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _20570_ (_12298_, _06251_, _12297_);
  nor _20571_ (_12300_, _12298_, _12295_);
  and _20572_ (_12301_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _20573_ (_12303_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _20574_ (_12304_, _12303_, _12301_);
  and _20575_ (_12305_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _20576_ (_12307_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _20577_ (_12308_, _12307_, _12305_);
  and _20578_ (_12310_, _12308_, _12304_);
  and _20579_ (_12311_, _12310_, _12300_);
  nor _20580_ (_12312_, _12311_, _07437_);
  nor _20581_ (_12313_, _12312_, _12294_);
  or _20582_ (_12314_, _12313_, _11836_);
  and _20583_ (_12315_, _12314_, _12292_);
  and _20584_ (_12316_, _11855_, _11852_);
  nor _20585_ (_12318_, _12316_, _11856_);
  nor _20586_ (_12319_, _12318_, _05341_);
  nor _20587_ (_12321_, _12319_, _05370_);
  nor _20588_ (_12322_, _12321_, _11843_);
  not _20589_ (_12323_, _12322_);
  and _20590_ (_12324_, _12323_, _11854_);
  or _20591_ (_12325_, _12324_, _11840_);
  or _20592_ (_12326_, _11868_, _11802_);
  and _20593_ (_12327_, _12326_, _12325_);
  nand _20594_ (_12328_, _12327_, _12315_);
  and _20595_ (_12329_, _12328_, _05375_);
  and _20596_ (_12330_, _12327_, _12315_);
  and _20597_ (_12332_, _12330_, _05911_);
  nor _20598_ (_12333_, _12332_, _12329_);
  and _20599_ (_12334_, _12333_, _05793_);
  and _20600_ (_12336_, _12334_, _12273_);
  and _20601_ (_12337_, _12336_, _12230_);
  and _20602_ (_12338_, _12337_, _12082_);
  and _20603_ (_12339_, _05460_, _05335_);
  nand _20604_ (_12340_, _12339_, _12338_);
  and _20605_ (_12341_, _12340_, _12184_);
  and _20606_ (_12343_, _12341_, _12088_);
  and _20607_ (_12344_, _12156_, _06873_);
  and _20608_ (_12345_, _12344_, _06610_);
  not _20609_ (_12346_, _07470_);
  and _20610_ (_12347_, _07105_, _06870_);
  and _20611_ (_12349_, _12347_, _12346_);
  and _20612_ (_12350_, _06870_, _06451_);
  nand _20613_ (_12351_, _12350_, _07038_);
  nor _20614_ (_12352_, _12347_, _11309_);
  and _20615_ (_12353_, _12352_, _12351_);
  not _20616_ (_12354_, _06828_);
  nand _20617_ (_12355_, _12135_, _12354_);
  and _20618_ (_12356_, _12355_, _06873_);
  nor _20619_ (_12357_, _12356_, _12097_);
  and _20620_ (_12358_, _12357_, _12353_);
  nor _20621_ (_12360_, _11283_, _06828_);
  and _20622_ (_12361_, _12360_, _12159_);
  and _20623_ (_12362_, _12361_, _12096_);
  and _20624_ (_12363_, _12362_, _12137_);
  nor _20625_ (_12364_, _12363_, _12094_);
  nor _20626_ (_12365_, _12344_, _12091_);
  not _20627_ (_12367_, _12365_);
  nor _20628_ (_12368_, _12367_, _12364_);
  and _20629_ (_12369_, _12368_, _12358_);
  and _20630_ (_12370_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _20631_ (_12371_, _12364_);
  and _20632_ (_12373_, _12358_, _12367_);
  and _20633_ (_12374_, _12373_, _12371_);
  and _20634_ (_12376_, \oc8051_top_1.oc8051_memory_interface1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _20635_ (_12377_, _12376_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _20636_ (_12378_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _20637_ (_12379_, _12378_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _20638_ (_12380_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _20639_ (_12381_, \oc8051_top_1.oc8051_memory_interface1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _20640_ (_12382_, _12381_, _12380_);
  and _20641_ (_12384_, _12382_, _12379_);
  and _20642_ (_12385_, _12384_, _12377_);
  and _20643_ (_12386_, _12385_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _20644_ (_12387_, _12385_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _20645_ (_12389_, _12387_, _12386_);
  and _20646_ (_12390_, _12389_, _12374_);
  not _20647_ (_12392_, _11309_);
  nor _20648_ (_12393_, _12392_, _06668_);
  or _20649_ (_12394_, _12393_, _12390_);
  or _20650_ (_12395_, _12394_, _12370_);
  or _20651_ (_12396_, _12395_, _12349_);
  nor _20652_ (_12397_, _12396_, _12345_);
  nand _20653_ (_12399_, _12397_, _12343_);
  and _20654_ (_12400_, _12358_, _12014_);
  nand _20655_ (_12401_, _12357_, _12353_);
  and _20656_ (_12402_, _12401_, _07176_);
  nor _20657_ (_12403_, _12402_, _12400_);
  not _20658_ (_12404_, _12403_);
  and _20659_ (_12405_, _12403_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _20660_ (_12406_, _12358_, _12067_);
  and _20661_ (_12407_, _12401_, _07582_);
  nor _20662_ (_12408_, _12407_, _12406_);
  and _20663_ (_12409_, _12408_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _20664_ (_12410_, _12403_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _20665_ (_12411_, _12410_, _12405_);
  and _20666_ (_12412_, _12411_, _12409_);
  or _20667_ (_12413_, _12412_, _12405_);
  nor _20668_ (_12414_, _12408_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _20669_ (_12415_, _12414_, _12409_);
  and _20670_ (_12416_, _12415_, _12411_);
  not _20671_ (_12417_, _07507_);
  or _20672_ (_12418_, _12401_, _12417_);
  nor _20673_ (_12419_, _05474_, _05578_);
  and _20674_ (_12420_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20675_ (_12421_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _20676_ (_12422_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _20677_ (_12423_, _12422_, _12421_);
  and _20678_ (_12424_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _20679_ (_12425_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _20680_ (_12426_, _12425_, _12424_);
  and _20681_ (_12427_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor _20682_ (_12428_, _06251_, _06207_);
  nor _20683_ (_12429_, _12428_, _12427_);
  and _20684_ (_12430_, _12429_, _12426_);
  and _20685_ (_12431_, _12430_, _12423_);
  nor _20686_ (_12432_, _12431_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20687_ (_12433_, _12432_, _12420_);
  nor _20688_ (_12434_, _12433_, _06200_);
  nor _20689_ (_12435_, _12434_, _12419_);
  not _20690_ (_12436_, _12435_);
  or _20691_ (_12437_, _12436_, _12358_);
  nand _20692_ (_12438_, _12437_, _12418_);
  or _20693_ (_12439_, _12438_, _05583_);
  and _20694_ (_12440_, _12358_, _07490_);
  nor _20695_ (_12441_, _05474_, _05117_);
  and _20696_ (_12442_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20697_ (_12443_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _20698_ (_12444_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _20699_ (_12445_, _12444_, _12443_);
  and _20700_ (_12446_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _20701_ (_12447_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _20702_ (_12448_, _12447_, _12446_);
  and _20703_ (_12449_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  not _20704_ (_12450_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _20705_ (_12451_, _06251_, _12450_);
  nor _20706_ (_12452_, _12451_, _12449_);
  and _20707_ (_12453_, _12452_, _12448_);
  and _20708_ (_12454_, _12453_, _12445_);
  nor _20709_ (_12455_, _12454_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20710_ (_12456_, _12455_, _12442_);
  nor _20711_ (_12457_, _12456_, _06200_);
  nor _20712_ (_12458_, _12457_, _12441_);
  and _20713_ (_12459_, _12458_, _12401_);
  nor _20714_ (_12460_, _12459_, _12440_);
  and _20715_ (_12461_, _12460_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand _20716_ (_12462_, _12438_, _05583_);
  and _20717_ (_12463_, _12462_, _12439_);
  nand _20718_ (_12464_, _12463_, _12461_);
  nand _20719_ (_12465_, _12464_, _12439_);
  and _20720_ (_12466_, _12465_, _12416_);
  or _20721_ (_12467_, _12466_, _12413_);
  and _20722_ (_12468_, _12358_, _07470_);
  and _20723_ (_12469_, _12401_, _07561_);
  nor _20724_ (_12470_, _12469_, _12468_);
  nor _20725_ (_12471_, _12470_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _20726_ (_12472_, _12470_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _20727_ (_12473_, _07454_);
  or _20728_ (_12474_, _12401_, _12473_);
  not _20729_ (_12475_, _07543_);
  or _20730_ (_12476_, _12358_, _12475_);
  nand _20731_ (_12477_, _12476_, _12474_);
  or _20732_ (_12478_, _12477_, _05220_);
  not _20733_ (_12479_, _12478_);
  not _20734_ (_12480_, _07439_);
  or _20735_ (_12481_, _12401_, _12480_);
  not _20736_ (_12482_, _07525_);
  or _20737_ (_12483_, _12358_, _12482_);
  and _20738_ (_12484_, _12483_, _12481_);
  nand _20739_ (_12485_, _12484_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _20740_ (_12486_, _12313_);
  or _20741_ (_12487_, _12401_, _12486_);
  nor _20742_ (_12488_, _05474_, _05236_);
  and _20743_ (_12489_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _20744_ (_12490_, _06245_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _20745_ (_12491_, _06257_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _20746_ (_12492_, _12491_, _12490_);
  and _20747_ (_12493_, _06243_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  not _20748_ (_12494_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _20749_ (_12495_, _06251_, _12494_);
  nor _20750_ (_12496_, _12495_, _12493_);
  and _20751_ (_12497_, _12496_, _12492_);
  and _20752_ (_12498_, _06260_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _20753_ (_12499_, _06262_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _20754_ (_12500_, _12499_, _12498_);
  and _20755_ (_12501_, _12500_, _12497_);
  nor _20756_ (_12502_, _12501_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20757_ (_12503_, _12502_, _12489_);
  nor _20758_ (_12504_, _12503_, _06200_);
  nor _20759_ (_12505_, _12504_, _12488_);
  not _20760_ (_12507_, _12505_);
  or _20761_ (_12508_, _12507_, _12358_);
  and _20762_ (_12509_, _12508_, _12487_);
  and _20763_ (_12510_, _12509_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _20764_ (_12512_, _12484_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _20765_ (_12513_, _12512_, _12485_);
  and _20766_ (_12514_, _12513_, _12510_);
  not _20767_ (_12515_, _12514_);
  nand _20768_ (_12516_, _12515_, _12485_);
  nand _20769_ (_12517_, _12477_, _05220_);
  and _20770_ (_12518_, _12517_, _12478_);
  and _20771_ (_12519_, _12518_, _12516_);
  or _20772_ (_12520_, _12519_, _12479_);
  nor _20773_ (_12521_, _12520_, _12472_);
  nor _20774_ (_12522_, _12521_, _12471_);
  nor _20775_ (_12523_, _12460_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _20776_ (_12524_, _12523_, _12461_);
  and _20777_ (_12525_, _12463_, _12524_);
  and _20778_ (_12526_, _12525_, _12416_);
  and _20779_ (_12527_, _12526_, _12522_);
  or _20780_ (_12528_, _12527_, _12467_);
  or _20781_ (_12529_, _12528_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _20782_ (_12530_, _12529_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _20783_ (_12531_, _12530_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _20784_ (_12532_, _12531_, _12404_);
  and _20785_ (_12533_, _12528_, _12377_);
  nor _20786_ (_12534_, _12533_, _12403_);
  or _20787_ (_12535_, _12534_, _12532_);
  nand _20788_ (_12536_, _12535_, _05195_);
  or _20789_ (_12537_, _12535_, _05195_);
  and _20790_ (_12538_, _12537_, _12536_);
  and _20791_ (_12539_, _12351_, _12371_);
  nor _20792_ (_12540_, _12539_, _12373_);
  and _20793_ (_12541_, _12540_, _12538_);
  or _20794_ (_12542_, _12541_, _12399_);
  not _20795_ (_12543_, _06205_);
  and _20796_ (_12544_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _20797_ (_12545_, _12544_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _20798_ (_12546_, _12545_, _12543_);
  and _20799_ (_12547_, _12546_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _20800_ (_12548_, _12547_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _20801_ (_12549_, _12548_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _20802_ (_12550_, _12549_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _20803_ (_12551_, _12550_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _20804_ (_12552_, _12551_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _20805_ (_12553_, _12552_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand _20806_ (_12554_, _12552_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _20807_ (_12555_, _12554_, _12553_);
  or _20808_ (_12556_, _12555_, _12343_);
  and _20809_ (_12557_, _12556_, _05110_);
  and _20810_ (_10697_, _12557_, _12542_);
  nand _20811_ (_12558_, _11239_, _05841_);
  and _20812_ (_12559_, _11222_, _11202_);
  and _20813_ (_12560_, _12559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _20814_ (_12561_, _12559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _20815_ (_12562_, _12561_, _12560_);
  and _20816_ (_12563_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _20817_ (_12564_, _12563_, _11202_);
  and _20818_ (_12565_, _12564_, _11223_);
  or _20819_ (_12566_, _12565_, _11193_);
  or _20820_ (_12567_, _12566_, _12562_);
  nor _20821_ (_12568_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor _20822_ (_12569_, _12568_, _11234_);
  and _20823_ (_12570_, _12569_, _12567_);
  and _20824_ (_12571_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _20825_ (_12572_, _12571_, _11239_);
  or _20826_ (_12573_, _12572_, _12570_);
  and _20827_ (_12574_, _12573_, _05110_);
  and _20828_ (_10705_, _12574_, _12558_);
  nor _20829_ (_12575_, _11712_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor _20830_ (_12576_, _12575_, _12559_);
  and _20831_ (_12577_, _11606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _20832_ (_12578_, _12577_, _11223_);
  or _20833_ (_12579_, _12578_, _11193_);
  or _20834_ (_12580_, _12579_, _12576_);
  or _20835_ (_12581_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _20836_ (_12583_, _12581_, _11584_);
  and _20837_ (_12584_, _12583_, _12580_);
  and _20838_ (_12585_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _20839_ (_12586_, _12585_, _12584_);
  nor _20840_ (_12587_, _11240_, _06054_);
  or _20841_ (_12588_, _12587_, _12586_);
  and _20842_ (_10709_, _12588_, _05110_);
  and _20843_ (_10712_, _11998_, _05110_);
  nor _20844_ (_10714_, _11783_, rst);
  and _20845_ (_12589_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _20846_ (_12590_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  or _20847_ (_12591_, _12590_, _12589_);
  and _20848_ (_10717_, _12591_, _05110_);
  or _20849_ (_12592_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  not _20850_ (_12594_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand _20851_ (_12595_, _06205_, _12594_);
  and _20852_ (_12596_, _12595_, _05110_);
  and _20853_ (_10720_, _12596_, _12592_);
  or _20854_ (_12597_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand _20855_ (_12598_, _06205_, _12494_);
  and _20856_ (_12599_, _12598_, _05110_);
  and _20857_ (_10724_, _12599_, _12597_);
  and _20858_ (_12601_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _20859_ (_12602_, _12601_, _11202_);
  and _20860_ (_12603_, _12602_, _11223_);
  and _20861_ (_12604_, _11206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor _20862_ (_12605_, _11206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _20863_ (_12606_, _12605_, _11193_);
  or _20864_ (_12607_, _12606_, _12604_);
  or _20865_ (_12608_, _12607_, _12603_);
  nor _20866_ (_12609_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nor _20867_ (_12610_, _12609_, _11234_);
  and _20868_ (_12611_, _12610_, _12608_);
  not _20869_ (_12612_, _11234_);
  nor _20870_ (_12613_, _12612_, _06229_);
  or _20871_ (_12615_, _12613_, _11239_);
  or _20872_ (_12616_, _12615_, _12611_);
  or _20873_ (_12617_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _20874_ (_12618_, _12617_, _05110_);
  and _20875_ (_10730_, _12618_, _12616_);
  nor _20876_ (_12619_, _12612_, _05841_);
  and _20877_ (_12620_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _20878_ (_12621_, _12620_, _11202_);
  and _20879_ (_12622_, _12621_, _11223_);
  nand _20880_ (_12623_, _11214_, _11202_);
  nor _20881_ (_12624_, _12623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _20882_ (_12625_, _12623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _20883_ (_12626_, _12625_, _11193_);
  or _20884_ (_12627_, _12626_, _12624_);
  or _20885_ (_12628_, _12627_, _12622_);
  nor _20886_ (_12629_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor _20887_ (_12630_, _12629_, _11234_);
  and _20888_ (_12631_, _12630_, _12628_);
  or _20889_ (_12632_, _12631_, _11239_);
  or _20890_ (_12633_, _12632_, _12619_);
  or _20891_ (_12634_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _20892_ (_12635_, _12634_, _05110_);
  and _20893_ (_10736_, _12635_, _12633_);
  and _20894_ (_12636_, _06024_, _05376_);
  and _20895_ (_12637_, _12636_, _06888_);
  and _20896_ (_12638_, _12637_, _05806_);
  not _20897_ (_12639_, _12638_);
  or _20898_ (_12640_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _20899_ (_12641_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _20900_ (_12642_, _12641_, _11202_);
  and _20901_ (_12643_, _12642_, _11223_);
  and _20902_ (_12645_, _11213_, _11202_);
  or _20903_ (_12646_, _12645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _20904_ (_12647_, _12646_, _12623_);
  or _20905_ (_12648_, _12647_, _11193_);
  or _20906_ (_12649_, _12648_, _12643_);
  and _20907_ (_12650_, _12649_, _12640_);
  and _20908_ (_12651_, _12650_, _12639_);
  nor _20909_ (_12652_, _12612_, _06054_);
  or _20910_ (_12653_, _12652_, _12651_);
  or _20911_ (_12654_, _12653_, _11239_);
  or _20912_ (_12655_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _20913_ (_12656_, _12655_, _05110_);
  and _20914_ (_10739_, _12656_, _12654_);
  or _20915_ (_12657_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _20916_ (_12658_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _20917_ (_12659_, _12658_, _11202_);
  and _20918_ (_12660_, _12659_, _11223_);
  and _20919_ (_12661_, _11212_, _11202_);
  nor _20920_ (_12662_, _12661_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor _20921_ (_12663_, _12662_, _12645_);
  or _20922_ (_12664_, _12663_, _11193_);
  or _20923_ (_12665_, _12664_, _12660_);
  and _20924_ (_12666_, _12665_, _12657_);
  and _20925_ (_12667_, _12666_, _12639_);
  nor _20926_ (_12668_, _12639_, _05334_);
  or _20927_ (_12669_, _12668_, _12667_);
  or _20928_ (_12670_, _12669_, _11239_);
  or _20929_ (_12671_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _20930_ (_12672_, _12671_, _05110_);
  and _20931_ (_10746_, _12672_, _12670_);
  and _20932_ (_12673_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _20933_ (_12674_, _12673_, _11202_);
  and _20934_ (_12675_, _12674_, _11223_);
  and _20935_ (_12676_, _11211_, _11202_);
  nor _20936_ (_12677_, _12676_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _20937_ (_12678_, _12677_, _12661_);
  or _20938_ (_12679_, _12678_, _11193_);
  or _20939_ (_12680_, _12679_, _12675_);
  nor _20940_ (_12681_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nor _20941_ (_12682_, _12681_, _11234_);
  and _20942_ (_12683_, _12682_, _12680_);
  nor _20943_ (_12684_, _12612_, _06088_);
  or _20944_ (_12686_, _12684_, _11239_);
  or _20945_ (_12687_, _12686_, _12683_);
  or _20946_ (_12688_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _20947_ (_12689_, _12688_, _05110_);
  and _20948_ (_10755_, _12689_, _12687_);
  and _20949_ (_12690_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _05110_);
  and _20950_ (_12691_, _12690_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not _20951_ (_12692_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _20952_ (_12693_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _20953_ (_12694_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _20954_ (_12695_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not _20955_ (_12696_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _20956_ (_12697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _20957_ (_12698_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _20958_ (_12699_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _20959_ (_12700_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _20960_ (_12701_, _11661_, _12700_);
  and _20961_ (_12702_, _12701_, _12699_);
  and _20962_ (_12703_, _12702_, _12698_);
  and _20963_ (_12704_, _12703_, _11657_);
  and _20964_ (_12705_, _12704_, _12697_);
  and _20965_ (_12706_, _12705_, _12696_);
  and _20966_ (_12707_, _12706_, _12695_);
  and _20967_ (_12708_, _12707_, _12694_);
  and _20968_ (_12709_, _12708_, _12693_);
  nor _20969_ (_12710_, _12709_, _12692_);
  and _20970_ (_12711_, _12709_, _12692_);
  nor _20971_ (_12712_, _12711_, _12710_);
  not _20972_ (_12713_, _12712_);
  nor _20973_ (_12714_, _12708_, _12693_);
  nor _20974_ (_12715_, _12714_, _12709_);
  nor _20975_ (_12716_, _12707_, _12694_);
  or _20976_ (_12717_, _12716_, _12708_);
  nor _20977_ (_12718_, _12706_, _12695_);
  nor _20978_ (_12719_, _12718_, _12707_);
  nor _20979_ (_12720_, _12705_, _12696_);
  nor _20980_ (_12722_, _12720_, _12706_);
  not _20981_ (_12723_, _12722_);
  nor _20982_ (_12724_, _12704_, _12697_);
  nor _20983_ (_12725_, _12724_, _12705_);
  not _20984_ (_12726_, _12725_);
  not _20985_ (_12727_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _20986_ (_12728_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _20987_ (_12729_, _12702_, _11657_);
  and _20988_ (_12730_, _12729_, _12728_);
  nor _20989_ (_12731_, _12730_, _12727_);
  or _20990_ (_12732_, _12731_, _12704_);
  and _20991_ (_12733_, _12701_, _11657_);
  nor _20992_ (_12734_, _12733_, _12699_);
  nor _20993_ (_12735_, _12734_, _12729_);
  not _20994_ (_12736_, _12735_);
  nor _20995_ (_12737_, _11662_, _12700_);
  or _20996_ (_12738_, _12737_, _12733_);
  and _20997_ (_12739_, _12738_, _11696_);
  and _20998_ (_12740_, _12739_, _12736_);
  nor _20999_ (_12741_, _12729_, _12728_);
  or _21000_ (_12742_, _12741_, _12730_);
  and _21001_ (_12743_, _12742_, _12740_);
  and _21002_ (_12744_, _12743_, _12732_);
  and _21003_ (_12745_, _12744_, _12726_);
  and _21004_ (_12747_, _12745_, _12723_);
  not _21005_ (_12748_, _12747_);
  nor _21006_ (_12749_, _12748_, _12719_);
  nand _21007_ (_12750_, _12749_, _12717_);
  or _21008_ (_12751_, _12750_, _12715_);
  nor _21009_ (_12752_, _12751_, _12713_);
  and _21010_ (_12753_, _12751_, _12713_);
  or _21011_ (_12754_, _12753_, _12752_);
  or _21012_ (_12755_, _12754_, _07437_);
  or _21013_ (_12756_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _21014_ (_12757_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and _21015_ (_12758_, _12757_, _12756_);
  and _21016_ (_12759_, _12758_, _12755_);
  or _21017_ (_10784_, _12759_, _12691_);
  and _21018_ (_12760_, _12344_, _06984_);
  nor _21019_ (_12761_, _12392_, _07028_);
  not _21020_ (_12762_, _12014_);
  and _21021_ (_12763_, _12347_, _12762_);
  and _21022_ (_12764_, _12386_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _21023_ (_12765_, _12764_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _21024_ (_12766_, _12765_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _21025_ (_12767_, _12766_, _05496_);
  or _21026_ (_12768_, _12766_, _05496_);
  and _21027_ (_12769_, _12768_, _12767_);
  and _21028_ (_12770_, _12769_, _12374_);
  and _21029_ (_12771_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _21030_ (_12772_, _12771_, _12770_);
  or _21031_ (_12773_, _12772_, _12763_);
  or _21032_ (_12775_, _12773_, _12761_);
  nor _21033_ (_12776_, _12775_, _12760_);
  nand _21034_ (_12777_, _12776_, _12343_);
  and _21035_ (_12778_, _12531_, _05195_);
  nor _21036_ (_12779_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _21037_ (_12780_, _12779_, _12778_);
  nand _21038_ (_12782_, _12780_, _05613_);
  and _21039_ (_12783_, _12782_, _12403_);
  and _21040_ (_12784_, _12533_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _21041_ (_12785_, _12784_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand _21042_ (_12786_, _12785_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _21043_ (_12787_, _12786_, _05613_);
  and _21044_ (_12788_, _12787_, _12404_);
  or _21045_ (_12789_, _12788_, _12783_);
  nand _21046_ (_12790_, _12789_, _05496_);
  or _21047_ (_12791_, _12789_, _05496_);
  and _21048_ (_12792_, _12791_, _12790_);
  and _21049_ (_12793_, _12792_, _12540_);
  or _21050_ (_12794_, _12793_, _12777_);
  and _21051_ (_12795_, _12545_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _21052_ (_12796_, _12795_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _21053_ (_12797_, _12796_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _21054_ (_12798_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _21055_ (_12799_, _12798_, _12797_);
  nand _21056_ (_12800_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _21057_ (_12801_, _12800_, _06205_);
  and _21058_ (_12802_, _12801_, _12799_);
  and _21059_ (_12803_, _12802_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _21060_ (_12804_, _12803_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _21061_ (_12805_, _12804_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand _21062_ (_12806_, _12805_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _21063_ (_12807_, _12805_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _21064_ (_12808_, _12807_, _12806_);
  or _21065_ (_12809_, _12808_, _12343_);
  and _21066_ (_12810_, _12809_, _05110_);
  and _21067_ (_10789_, _12810_, _12794_);
  and _21068_ (_10803_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _05110_);
  nor _21069_ (_12811_, _11309_, rst);
  and _21070_ (_10813_, _12811_, _12343_);
  and _21071_ (_12812_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor _21072_ (_12813_, _06229_, _06000_);
  and _21073_ (_12814_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or _21074_ (_12815_, _12814_, _12813_);
  and _21075_ (_12816_, _12815_, _05337_);
  or _21076_ (_12817_, _12816_, _12812_);
  and _21077_ (_10862_, _12817_, _05110_);
  and _21078_ (_12818_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _21079_ (_12819_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or _21080_ (_12820_, _12819_, _12818_);
  and _21081_ (_10880_, _12820_, _05110_);
  or _21082_ (_12821_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand _21083_ (_12822_, _06205_, _07514_);
  and _21084_ (_12823_, _12822_, _05110_);
  and _21085_ (_10883_, _12823_, _12821_);
  and _21086_ (_12824_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _21087_ (_12825_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  or _21088_ (_12826_, _12825_, _12824_);
  and _21089_ (_10935_, _12826_, _05110_);
  and _21090_ (_12827_, _08287_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not _21091_ (_12828_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _21092_ (_12829_, _08280_, _12828_);
  nor _21093_ (_12830_, _12829_, _08287_);
  or _21094_ (_12831_, _12830_, _12827_);
  nor _21095_ (_12832_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor _21096_ (_12833_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _21097_ (_12834_, _12833_, _12832_);
  nor _21098_ (_12835_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor _21099_ (_12836_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _21100_ (_12837_, _12836_, _12835_);
  and _21101_ (_12838_, _12837_, _12834_);
  nor _21102_ (_12839_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _21103_ (_12841_, _12839_, _12838_);
  and _21104_ (_12843_, _12841_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _21105_ (_12844_, _12843_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _21106_ (_12845_, _12844_, _08280_);
  nor _21107_ (_12847_, _12845_, _12831_);
  nor _21108_ (_12848_, _12847_, _08274_);
  nor _21109_ (_12849_, _08236_, _06798_);
  and _21110_ (_12850_, _12849_, _08274_);
  or _21111_ (_12851_, _12850_, _12848_);
  and _21112_ (_10942_, _12851_, _05110_);
  and _21113_ (_12853_, _08297_, _06194_);
  and _21114_ (_12854_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and _21115_ (_12855_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _21116_ (_12856_, _12855_, _12854_);
  nor _21117_ (_12857_, _12856_, _08274_);
  and _21118_ (_12858_, _08276_, _06230_);
  or _21119_ (_12859_, _12858_, _12857_);
  or _21120_ (_12860_, _12859_, _12853_);
  and _21121_ (_10966_, _12860_, _05110_);
  and _21122_ (_12861_, _08297_, _06230_);
  and _21123_ (_12862_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _21124_ (_12863_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor _21125_ (_12864_, _12863_, _12862_);
  nor _21126_ (_12865_, _12864_, _08274_);
  and _21127_ (_12866_, _08276_, _06559_);
  or _21128_ (_12867_, _12866_, _12865_);
  or _21129_ (_12868_, _12867_, _12861_);
  and _21130_ (_10974_, _12868_, _05110_);
  nor _21131_ (_10979_, _12313_, rst);
  and _21132_ (_12869_, _08297_, _06183_);
  and _21133_ (_12870_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _21134_ (_12871_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor _21135_ (_12872_, _12871_, _12870_);
  nor _21136_ (_12873_, _12872_, _08274_);
  not _21137_ (_12874_, _05334_);
  and _21138_ (_12875_, _08276_, _12874_);
  or _21139_ (_12876_, _12875_, _12873_);
  or _21140_ (_12877_, _12876_, _12869_);
  and _21141_ (_10985_, _12877_, _05110_);
  and _21142_ (_12878_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not _21143_ (_12879_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _21144_ (_12880_, pc_log_change, _12879_);
  or _21145_ (_12881_, _12880_, _12878_);
  and _21146_ (_11004_, _12881_, _05110_);
  and _21147_ (_12882_, _08297_, _12874_);
  and _21148_ (_12883_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _21149_ (_12884_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _21150_ (_12885_, _12884_, _12883_);
  nor _21151_ (_12887_, _12885_, _08274_);
  and _21152_ (_12888_, _08276_, _06194_);
  or _21153_ (_12889_, _12888_, _12887_);
  or _21154_ (_12890_, _12889_, _12882_);
  and _21155_ (_11006_, _12890_, _05110_);
  nand _21156_ (_12891_, _11280_, _07418_);
  or _21157_ (_12892_, _11280_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _21158_ (_12893_, _12892_, _05110_);
  and _21159_ (_11058_, _12893_, _12891_);
  not _21160_ (_12894_, _05901_);
  and _21161_ (_12895_, _08297_, _12894_);
  and _21162_ (_12896_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _21163_ (_12897_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor _21164_ (_12898_, _12897_, _12896_);
  nor _21165_ (_12899_, _12898_, _08274_);
  and _21166_ (_12900_, _08276_, _08224_);
  or _21167_ (_12901_, _12900_, _12899_);
  or _21168_ (_12902_, _12901_, _12895_);
  and _21169_ (_11073_, _12902_, _05110_);
  and _21170_ (_12903_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not _21171_ (_12904_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _21172_ (_12905_, _06205_, _12904_);
  or _21173_ (_12906_, _12905_, _12903_);
  and _21174_ (_11095_, _12906_, _05110_);
  and _21175_ (_12907_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not _21176_ (_12908_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _21177_ (_12909_, _06205_, _12908_);
  or _21178_ (_12910_, _12909_, _12907_);
  and _21179_ (_11112_, _12910_, _05110_);
  and _21180_ (_12911_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor _21181_ (_12912_, _06205_, _07571_);
  or _21182_ (_12913_, _12912_, _12911_);
  and _21183_ (_11115_, _12913_, _05110_);
  and _21184_ (_12914_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor _21185_ (_12915_, _06205_, _07514_);
  or _21186_ (_12916_, _12915_, _12914_);
  and _21187_ (_11121_, _12916_, _05110_);
  and _21188_ (_11126_, _11576_, _05110_);
  not _21189_ (_12917_, _06895_);
  or _21190_ (_12918_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  not _21191_ (_12919_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand _21192_ (_12920_, _08884_, _12919_);
  and _21193_ (_12921_, _12920_, _12918_);
  and _21194_ (_12922_, _12921_, _12917_);
  nor _21195_ (_12923_, _12917_, _06088_);
  or _21196_ (_12924_, _12923_, _12922_);
  and _21197_ (_11138_, _12924_, _05110_);
  or _21198_ (_12925_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand _21199_ (_12926_, _06205_, _12297_);
  and _21200_ (_12927_, _12926_, _05110_);
  and _21201_ (_11148_, _12927_, _12925_);
  or _21202_ (_12928_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand _21203_ (_12929_, _06205_, _06330_);
  and _21204_ (_12930_, _12929_, _05110_);
  and _21205_ (_11150_, _12930_, _12928_);
  or _21206_ (_12931_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand _21207_ (_12932_, _06205_, _07474_);
  and _21208_ (_12933_, _12932_, _05110_);
  and _21209_ (_11154_, _12933_, _12931_);
  and _21210_ (_12934_, _08297_, _08224_);
  and _21211_ (_12935_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _21212_ (_12936_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor _21213_ (_12937_, _12936_, _12935_);
  nor _21214_ (_12938_, _12937_, _08274_);
  and _21215_ (_12939_, _08276_, _06183_);
  or _21216_ (_12940_, _12939_, _12938_);
  or _21217_ (_12942_, _12940_, _12934_);
  and _21218_ (_11161_, _12942_, _05110_);
  and _21219_ (_12943_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _21220_ (_12944_, _12738_, _11696_);
  nor _21221_ (_12946_, _12944_, _12739_);
  or _21222_ (_12947_, _12946_, _07437_);
  or _21223_ (_12948_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _21224_ (_12949_, _12948_, _11510_);
  and _21225_ (_12950_, _12949_, _12947_);
  or _21226_ (_12952_, _12950_, _12943_);
  and _21227_ (_11164_, _12952_, _05110_);
  and _21228_ (_12953_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _21229_ (_12954_, _12743_, _12732_);
  nor _21230_ (_12955_, _12954_, _12744_);
  or _21231_ (_12956_, _12955_, _07437_);
  or _21232_ (_12957_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _21233_ (_12958_, _12957_, _11510_);
  and _21234_ (_12959_, _12958_, _12956_);
  or _21235_ (_12960_, _12959_, _12953_);
  and _21236_ (_11195_, _12960_, _05110_);
  or _21237_ (_12961_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand _21238_ (_12962_, _06205_, _07532_);
  and _21239_ (_12963_, _12962_, _05110_);
  and _21240_ (_11198_, _12963_, _12961_);
  nor _21241_ (_12964_, _12742_, _12740_);
  nor _21242_ (_12965_, _12964_, _12743_);
  or _21243_ (_12966_, _12965_, _07437_);
  or _21244_ (_12967_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _21245_ (_12968_, _12967_, _11510_);
  and _21246_ (_12969_, _12968_, _12966_);
  and _21247_ (_12970_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _21248_ (_12971_, _12970_, _12969_);
  and _21249_ (_11201_, _12971_, _05110_);
  and _21250_ (_12972_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _21251_ (_12973_, _12739_, _12736_);
  nor _21252_ (_12974_, _12973_, _12740_);
  or _21253_ (_12975_, _12974_, _07437_);
  or _21254_ (_12976_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _21255_ (_12977_, _12976_, _11510_);
  and _21256_ (_12978_, _12977_, _12975_);
  or _21257_ (_12979_, _12978_, _12972_);
  and _21258_ (_11210_, _12979_, _05110_);
  or _21259_ (_12980_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand _21260_ (_12981_, _06205_, _06352_);
  and _21261_ (_12982_, _12981_, _05110_);
  and _21262_ (_11221_, _12982_, _12980_);
  and _21263_ (_12983_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  not _21264_ (_12984_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _21265_ (_12985_, _06205_, _12984_);
  or _21266_ (_12986_, _12985_, _12983_);
  and _21267_ (_11224_, _12986_, _05110_);
  and _21268_ (_12987_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor _21269_ (_12988_, _06205_, _07532_);
  or _21270_ (_12989_, _12988_, _12987_);
  and _21271_ (_11229_, _12989_, _05110_);
  or _21272_ (_12990_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand _21273_ (_12991_, _06205_, _07425_);
  and _21274_ (_12992_, _12991_, _05110_);
  and _21275_ (_11244_, _12992_, _12990_);
  or _21276_ (_12993_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand _21277_ (_12994_, _06205_, _06370_);
  and _21278_ (_12995_, _12994_, _05110_);
  and _21279_ (_11267_, _12995_, _12993_);
  and _21280_ (_12996_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor _21281_ (_12997_, _06205_, _07553_);
  or _21282_ (_12998_, _12997_, _12996_);
  and _21283_ (_11270_, _12998_, _05110_);
  or _21284_ (_12999_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand _21285_ (_13000_, _06205_, _07494_);
  and _21286_ (_13001_, _13000_, _05110_);
  and _21287_ (_11278_, _13001_, _12999_);
  nand _21288_ (_13002_, _11280_, _06512_);
  or _21289_ (_13003_, _11280_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _21290_ (_13004_, _13003_, _05110_);
  and _21291_ (_11285_, _13004_, _13002_);
  or _21292_ (_13005_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand _21293_ (_13006_, _06205_, _06397_);
  and _21294_ (_13007_, _13006_, _05110_);
  and _21295_ (_11291_, _13007_, _13005_);
  or _21296_ (_13008_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand _21297_ (_13009_, _06205_, _07457_);
  and _21298_ (_13010_, _13009_, _05110_);
  and _21299_ (_11318_, _13010_, _13008_);
  or _21300_ (_13011_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand _21301_ (_13012_, _06205_, _07442_);
  and _21302_ (_13013_, _13012_, _05110_);
  and _21303_ (_11352_, _13013_, _13011_);
  or _21304_ (_13014_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand _21305_ (_13015_, _06205_, _06248_);
  and _21306_ (_13016_, _13015_, _05110_);
  and _21307_ (_11361_, _13016_, _13014_);
  or _21308_ (_13017_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand _21309_ (_13018_, _06205_, _06413_);
  and _21310_ (_13019_, _13018_, _05110_);
  and _21311_ (_11364_, _13019_, _13017_);
  or _21312_ (_13020_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand _21313_ (_13021_, _06205_, _06285_);
  and _21314_ (_13023_, _13021_, _05110_);
  and _21315_ (_11375_, _13023_, _13020_);
  or _21316_ (_13024_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand _21317_ (_13025_, _06205_, _06307_);
  and _21318_ (_13026_, _13025_, _05110_);
  and _21319_ (_11390_, _13026_, _13024_);
  and _21320_ (_13028_, _06177_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _21321_ (_13029_, _06184_, _12894_);
  or _21322_ (_13030_, _13029_, _13028_);
  and _21323_ (_11392_, _13030_, _05110_);
  or _21324_ (_13031_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand _21325_ (_13032_, _06205_, _12054_);
  and _21326_ (_13033_, _13032_, _05110_);
  and _21327_ (_11413_, _13033_, _13031_);
  and _21328_ (_13034_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _07601_);
  and _21329_ (_13035_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21330_ (_13036_, _13035_, _13034_);
  and _21331_ (_11496_, _13036_, _05110_);
  nor _21332_ (_11509_, _11580_, rst);
  and _21333_ (_11514_, _11570_, _05110_);
  and _21334_ (_13037_, _07601_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and _21335_ (_13038_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _21336_ (_13039_, _13038_, _13037_);
  and _21337_ (_11522_, _13039_, _05110_);
  and _21338_ (_13040_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _07601_);
  and _21339_ (_13041_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21340_ (_13042_, _13041_, _13040_);
  and _21341_ (_11531_, _13042_, _05110_);
  and _21342_ (_13043_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _07601_);
  and _21343_ (_13044_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21344_ (_13045_, _13044_, _13043_);
  and _21345_ (_11534_, _13045_, _05110_);
  and _21346_ (_13046_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor _21347_ (_13047_, _06205_, _12494_);
  or _21348_ (_13048_, _13047_, _13046_);
  and _21349_ (_11624_, _13048_, _05110_);
  and _21350_ (_13049_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor _21351_ (_13050_, _06205_, _06207_);
  or _21352_ (_13051_, _13050_, _13049_);
  and _21353_ (_11643_, _13051_, _05110_);
  and _21354_ (_13052_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor _21355_ (_13053_, _06205_, _12450_);
  or _21356_ (_13054_, _13053_, _13052_);
  and _21357_ (_11649_, _13054_, _05110_);
  and _21358_ (_13055_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _21359_ (_13056_, _06205_, _09467_);
  or _21360_ (_13057_, _13056_, _13055_);
  and _21361_ (_11659_, _13057_, _05110_);
  and _21362_ (_13058_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor _21363_ (_13059_, _06205_, _07167_);
  or _21364_ (_13060_, _13059_, _13058_);
  and _21365_ (_11663_, _13060_, _05110_);
  and _21366_ (_13061_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not _21367_ (_13062_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _21368_ (_13063_, _06205_, _13062_);
  or _21369_ (_13064_, _13063_, _13061_);
  and _21370_ (_11668_, _13064_, _05110_);
  and _21371_ (_13065_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  not _21372_ (_13066_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _21373_ (_13067_, _06205_, _13066_);
  or _21374_ (_13068_, _13067_, _13065_);
  and _21375_ (_11674_, _13068_, _05110_);
  and _21376_ (_13069_, _06807_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or _21377_ (_13070_, _11728_, _07120_);
  or _21378_ (_13071_, _13070_, _11732_);
  and _21379_ (_13072_, _06463_, _06448_);
  and _21380_ (_13073_, _11283_, _06342_);
  or _21381_ (_13074_, _13073_, _13072_);
  or _21382_ (_13075_, _13074_, _13071_);
  and _21383_ (_13076_, _06849_, _06277_);
  or _21384_ (_13077_, _12158_, _12138_);
  and _21385_ (_13078_, _06856_, _06434_);
  and _21386_ (_13079_, _07080_, _06451_);
  or _21387_ (_13080_, _13079_, _13078_);
  or _21388_ (_13081_, _13080_, _13077_);
  or _21389_ (_13082_, _13081_, _13076_);
  or _21390_ (_13083_, _13082_, _06940_);
  or _21391_ (_13084_, _13083_, _13075_);
  and _21392_ (_13085_, _13084_, _06842_);
  or _21393_ (_11679_, _13085_, _13069_);
  and _21394_ (_13086_, _06852_, _06276_);
  or _21395_ (_13087_, _06451_, _06447_);
  nand _21396_ (_13088_, _13087_, _13086_);
  and _21397_ (_13089_, _13088_, _06858_);
  or _21398_ (_13090_, _06849_, _06954_);
  or _21399_ (_11694_, _13090_, _13089_);
  and _21400_ (_13091_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  not _21401_ (_13092_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _21402_ (_13093_, _06205_, _13092_);
  or _21403_ (_13094_, _13093_, _13091_);
  and _21404_ (_11697_, _13094_, _05110_);
  and _21405_ (_13095_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not _21406_ (_13096_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _21407_ (_13097_, pc_log_change, _13096_);
  or _21408_ (_13098_, _13097_, _13095_);
  and _21409_ (_11702_, _13098_, _05110_);
  and _21410_ (_11704_, _11321_, _05110_);
  and _21411_ (_13099_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _21412_ (_13100_, _06205_, _12594_);
  or _21413_ (_13101_, _13100_, _13099_);
  and _21414_ (_11707_, _13101_, _05110_);
  and _21415_ (_13102_, _11412_, _06915_);
  and _21416_ (_13103_, _11358_, _06926_);
  or _21417_ (_13104_, _13103_, _11395_);
  nor _21418_ (_13105_, _13104_, _13102_);
  nand _21419_ (_13106_, _13105_, _11439_);
  or _21420_ (_13107_, _13106_, _11459_);
  and _21421_ (_13109_, _11387_, _11365_);
  and _21422_ (_13110_, _11342_, _06922_);
  and _21423_ (_13111_, _11345_, _06924_);
  or _21424_ (_13112_, _13111_, _13110_);
  or _21425_ (_13113_, _13112_, _13109_);
  or _21426_ (_13114_, _11441_, _11427_);
  and _21427_ (_13115_, _11412_, _11365_);
  or _21428_ (_13116_, _13115_, _11476_);
  or _21429_ (_13117_, _13116_, _13114_);
  or _21430_ (_13118_, _13117_, _13113_);
  or _21431_ (_13119_, _13118_, _13107_);
  or _21432_ (_13120_, _13119_, _06933_);
  and _21433_ (_13121_, _13120_, _05475_);
  nor _21434_ (_13122_, _06908_, _06238_);
  or _21435_ (_13123_, _13122_, rst);
  or _21436_ (_11718_, _13123_, _13121_);
  and _21437_ (_11725_, _11312_, _05110_);
  nor _21438_ (_13124_, _11484_, _11482_);
  nor _21439_ (_13125_, _13124_, _11485_);
  or _21440_ (_13126_, _13125_, _06200_);
  or _21441_ (_13127_, _05474_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _21442_ (_13128_, _13127_, _12757_);
  and _21443_ (_11733_, _13128_, _13126_);
  and _21444_ (_13129_, _11481_, _05474_);
  nand _21445_ (_13130_, _13129_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _21446_ (_13131_, _13129_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _21447_ (_13132_, _13131_, _12757_);
  and _21448_ (_11739_, _13132_, _13130_);
  nand _21449_ (_13133_, _06673_, _06229_);
  or _21450_ (_13134_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _21451_ (_13135_, _13134_, _05110_);
  and _21452_ (_11913_, _13135_, _13133_);
  nand _21453_ (_13136_, _11280_, _06668_);
  or _21454_ (_13137_, _11280_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _21455_ (_13138_, _13137_, _05110_);
  and _21456_ (_11940_, _13138_, _13136_);
  nand _21457_ (_13139_, _11280_, _07337_);
  or _21458_ (_13140_, _11280_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _21459_ (_13141_, _13140_, _05110_);
  and _21460_ (_11947_, _13141_, _13139_);
  or _21461_ (_13142_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nand _21462_ (_13143_, _06205_, _13062_);
  and _21463_ (_13144_, _13143_, _05110_);
  and _21464_ (_11980_, _13144_, _13142_);
  and _21465_ (_13145_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _21466_ (_13146_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor _21467_ (_13147_, _13146_, _13145_);
  nor _21468_ (_13148_, _13147_, _08274_);
  or _21469_ (_13149_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _11264_);
  and _21470_ (_13150_, _13149_, _08236_);
  and _21471_ (_13151_, _13150_, _08274_);
  or _21472_ (_13152_, _13151_, _13148_);
  and _21473_ (_11983_, _13152_, _05110_);
  or _21474_ (_13153_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand _21475_ (_13154_, _06205_, _07571_);
  and _21476_ (_13156_, _13154_, _05110_);
  and _21477_ (_11991_, _13156_, _13153_);
  and _21478_ (_13157_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _21479_ (_13158_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or _21480_ (_13159_, _13158_, _13157_);
  and _21481_ (_12015_, _13159_, _05110_);
  and _21482_ (_13160_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _21483_ (_13161_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  or _21484_ (_13162_, _13161_, _13160_);
  and _21485_ (_12019_, _13162_, _05110_);
  and _21486_ (_12047_, _11944_, _05110_);
  nor _21487_ (_12055_, _12067_, rst);
  and _21488_ (_13163_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _21489_ (_13164_, _13163_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _21490_ (_12069_, _13164_, _05110_);
  and _21491_ (_13165_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _21492_ (_13166_, _13165_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _21493_ (_12076_, _13166_, _05110_);
  and _21494_ (_13167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _05110_);
  and _21495_ (_13168_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _05110_);
  and _21496_ (_13170_, _13168_, _11505_);
  or _21497_ (_12079_, _13170_, _13167_);
  nor _21498_ (_12081_, _12435_, rst);
  and _21499_ (_13171_, _08869_, _05804_);
  nand _21500_ (_13172_, _13171_, _05841_);
  not _21501_ (_13174_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _21502_ (_13175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _13174_);
  not _21503_ (_13176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _21504_ (_13177_, _13176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nor _21505_ (_13178_, _13177_, _13175_);
  and _21506_ (_13179_, _11238_, _05804_);
  nor _21507_ (_13180_, _13179_, _13178_);
  not _21508_ (_13181_, _13180_);
  and _21509_ (_13182_, _13181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  not _21510_ (_13183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _21511_ (_13184_, t1_i);
  and _21512_ (_13185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _13184_);
  nor _21513_ (_13186_, _13185_, _13183_);
  not _21514_ (_13187_, _13186_);
  not _21515_ (_13188_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _21516_ (_13189_, _13188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _21517_ (_13190_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _21518_ (_13191_, _13190_);
  and _21519_ (_13192_, _13191_, _13189_);
  and _21520_ (_13193_, _13192_, _13187_);
  and _21521_ (_13194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _21522_ (_13195_, _13194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _21523_ (_13196_, _13195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _21524_ (_13197_, _13196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _21525_ (_13198_, _13197_, _13193_);
  and _21526_ (_13199_, _13198_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _21527_ (_13200_, _13199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _21528_ (_13201_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _21529_ (_13202_, _13201_, _13198_);
  nor _21530_ (_13203_, _13202_, _13200_);
  and _21531_ (_13204_, _13180_, _13203_);
  and _21532_ (_13205_, _13199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _21533_ (_13206_, _13205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _21534_ (_13207_, _13206_, _13175_);
  nand _21535_ (_13208_, _13207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _21536_ (_13209_, _13208_, _13179_);
  or _21537_ (_13210_, _13209_, _13204_);
  or _21538_ (_13211_, _13210_, _13182_);
  or _21539_ (_13212_, _13171_, _13211_);
  and _21540_ (_13213_, _13212_, _05110_);
  and _21541_ (_12085_, _13213_, _13172_);
  and _21542_ (_13214_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _21543_ (_13215_, _13214_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _21544_ (_12107_, _13215_, _05110_);
  and _21545_ (_13216_, _13196_, _13193_);
  nor _21546_ (_13217_, _13216_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _21547_ (_13218_, _13217_, _13198_);
  and _21548_ (_13219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nor _21549_ (_13220_, _13219_, _13179_);
  and _21550_ (_13221_, _13220_, _13218_);
  not _21551_ (_13222_, _13220_);
  and _21552_ (_13223_, _13222_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand _21553_ (_13224_, _13207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _21554_ (_13225_, _13224_, _13179_);
  or _21555_ (_13226_, _13225_, _13223_);
  or _21556_ (_13227_, _13226_, _13221_);
  or _21557_ (_13228_, _13227_, _13171_);
  nand _21558_ (_13229_, _13171_, _05334_);
  and _21559_ (_13230_, _13229_, _05110_);
  and _21560_ (_12110_, _13230_, _13228_);
  and _21561_ (_13231_, _13195_, _13193_);
  nor _21562_ (_13232_, _13231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _21563_ (_13233_, _13232_, _13216_);
  and _21564_ (_13234_, _13233_, _13220_);
  and _21565_ (_13235_, _13222_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _21566_ (_13236_, _13235_, _13234_);
  nand _21567_ (_13237_, _13207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _21568_ (_13238_, _13237_, _13179_);
  or _21569_ (_13239_, _13238_, _13171_);
  or _21570_ (_13240_, _13239_, _13236_);
  nand _21571_ (_13241_, _13171_, _06088_);
  and _21572_ (_13242_, _13241_, _05110_);
  and _21573_ (_12113_, _13242_, _13240_);
  and _21574_ (_13243_, _13193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _21575_ (_13244_, _13243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _21576_ (_13245_, _13244_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _21577_ (_13246_, _13245_, _13231_);
  nand _21578_ (_13247_, _13246_, _13220_);
  or _21579_ (_13248_, _13220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _21580_ (_13249_, _13248_, _13247_);
  and _21581_ (_13250_, _06894_, _05804_);
  and _21582_ (_13251_, _13202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _21583_ (_13252_, _13251_, _13175_);
  nand _21584_ (_13253_, _13252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _21585_ (_13254_, _13253_, _13179_);
  or _21586_ (_13255_, _13254_, _13250_);
  or _21587_ (_13256_, _13255_, _13249_);
  nand _21588_ (_13257_, _13250_, _06229_);
  and _21589_ (_13258_, _13257_, _05110_);
  and _21590_ (_12116_, _13258_, _13256_);
  nand _21591_ (_13259_, _13171_, _06054_);
  nand _21592_ (_13260_, _13207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _21593_ (_13261_, _13260_, _13179_);
  nor _21594_ (_13262_, _13198_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _21595_ (_13263_, _13262_, _13199_);
  and _21596_ (_13264_, _13263_, _13180_);
  and _21597_ (_13265_, _13181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _21598_ (_13266_, _13265_, _13264_);
  or _21599_ (_13267_, _13266_, _13261_);
  or _21600_ (_13268_, _13267_, _13171_);
  and _21601_ (_13269_, _13268_, _05110_);
  and _21602_ (_12122_, _13269_, _13259_);
  or _21603_ (_13270_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand _21604_ (_13271_, _06205_, _12908_);
  and _21605_ (_13272_, _13271_, _05110_);
  and _21606_ (_12124_, _13272_, _13270_);
  and _21607_ (_13273_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _21608_ (_13274_, _13273_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _21609_ (_12129_, _13274_, _05110_);
  not _21610_ (_13275_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _21611_ (_13276_, _13220_, _13275_);
  or _21612_ (_13277_, _13193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor _21613_ (_13278_, _13219_, _13243_);
  and _21614_ (_13279_, _13175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _21615_ (_13280_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _21616_ (_13281_, _13280_, _13201_);
  and _21617_ (_13282_, _13281_, _13197_);
  and _21618_ (_13283_, _13282_, _13279_);
  or _21619_ (_13284_, _13283_, _13278_);
  nand _21620_ (_13285_, _13284_, _13277_);
  nor _21621_ (_13286_, _13285_, _13179_);
  or _21622_ (_13287_, _13286_, _13250_);
  or _21623_ (_13288_, _13287_, _13276_);
  nand _21624_ (_13289_, _13250_, _06798_);
  and _21625_ (_13290_, _13289_, _05110_);
  and _21626_ (_12133_, _13290_, _13288_);
  nor _21627_ (_13291_, _13243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _21628_ (_13292_, _13291_, _13244_);
  nand _21629_ (_13294_, _13292_, _13220_);
  or _21630_ (_13295_, _13220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _21631_ (_13296_, _13295_, _13294_);
  nand _21632_ (_13297_, _13252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _21633_ (_13298_, _13297_, _13179_);
  or _21634_ (_13299_, _13298_, _13250_);
  or _21635_ (_13300_, _13299_, _13296_);
  nand _21636_ (_13301_, _13250_, _05938_);
  and _21637_ (_13302_, _13301_, _05110_);
  and _21638_ (_12136_, _13302_, _13300_);
  and _21639_ (_13303_, _12528_, _12376_);
  or _21640_ (_13304_, _13303_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _21641_ (_13305_, _13304_, _12534_);
  and _21642_ (_13306_, _12530_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _21643_ (_13308_, _13306_, _12531_);
  and _21644_ (_13309_, _13308_, _12403_);
  or _21645_ (_13310_, _13309_, _13305_);
  and _21646_ (_13311_, _13310_, _12540_);
  and _21647_ (_13312_, _12344_, _07305_);
  and _21648_ (_13313_, _12374_, _06918_);
  and _21649_ (_13314_, _12347_, _12473_);
  and _21650_ (_13315_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _21651_ (_13316_, _12392_, _07337_);
  or _21652_ (_13317_, _13316_, _13315_);
  or _21653_ (_13318_, _13317_, _13314_);
  or _21654_ (_13319_, _13318_, _13313_);
  nor _21655_ (_13320_, _13319_, _13312_);
  nand _21656_ (_13321_, _13320_, _12343_);
  or _21657_ (_13322_, _13321_, _13311_);
  nor _21658_ (_13323_, _12551_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _21659_ (_13324_, _13323_, _12552_);
  or _21660_ (_13325_, _13324_, _12343_);
  and _21661_ (_13326_, _13325_, _05110_);
  and _21662_ (_12139_, _13326_, _13322_);
  and _21663_ (_13327_, _07038_, _06870_);
  and _21664_ (_13328_, _13327_, _06451_);
  nor _21665_ (_13329_, _13328_, _12364_);
  nor _21666_ (_13330_, _13329_, _12373_);
  not _21667_ (_13331_, _12461_);
  nand _21668_ (_13332_, _12524_, _12522_);
  nand _21669_ (_13333_, _13332_, _13331_);
  or _21670_ (_13334_, _12463_, _13333_);
  nand _21671_ (_13335_, _12463_, _13333_);
  and _21672_ (_13336_, _13335_, _13334_);
  and _21673_ (_13337_, _13336_, _13330_);
  and _21674_ (_13338_, _12436_, _12347_);
  not _21675_ (_13339_, _06548_);
  or _21676_ (_13340_, _12369_, _12344_);
  and _21677_ (_13341_, _13340_, _13339_);
  and _21678_ (_13342_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _21679_ (_13343_, _12374_, _12417_);
  or _21680_ (_13344_, _13343_, _13342_);
  or _21681_ (_13345_, _13344_, _13341_);
  or _21682_ (_13346_, _13345_, _13338_);
  or _21683_ (_13348_, _13346_, _13337_);
  and _21684_ (_13349_, _13348_, _12343_);
  nor _21685_ (_13350_, _12546_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _21686_ (_13351_, _13350_, _12547_);
  nor _21687_ (_13352_, _13351_, _12343_);
  or _21688_ (_13353_, _13352_, _13349_);
  and _21689_ (_12143_, _13353_, _05110_);
  nand _21690_ (_13354_, _13179_, _06798_);
  not _21691_ (_13355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _21692_ (_13356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _21693_ (_13358_, _13356_, _13198_);
  and _21694_ (_13359_, _13251_, _13177_);
  nor _21695_ (_13361_, _13359_, _13358_);
  nor _21696_ (_13362_, _13361_, _13355_);
  and _21697_ (_13363_, _13361_, _13355_);
  nor _21698_ (_13364_, _13363_, _13362_);
  or _21699_ (_13365_, _13364_, _13179_);
  and _21700_ (_13366_, _13365_, _13354_);
  or _21701_ (_13367_, _13366_, _13171_);
  nand _21702_ (_13368_, _13171_, _13355_);
  and _21703_ (_13369_, _13368_, _05110_);
  and _21704_ (_12152_, _13369_, _13367_);
  nand _21705_ (_13370_, _13179_, _05938_);
  not _21706_ (_13371_, _13171_);
  nor _21707_ (_13372_, _13362_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _21708_ (_13373_, _13362_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _21709_ (_13374_, _13373_, _13372_);
  or _21710_ (_13375_, _13374_, _13179_);
  and _21711_ (_13376_, _13375_, _13371_);
  and _21712_ (_13377_, _13376_, _13370_);
  and _21713_ (_13378_, _13250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _21714_ (_13379_, _13378_, _13377_);
  and _21715_ (_12155_, _13379_, _05110_);
  nor _21716_ (_13380_, _11693_, _11690_);
  nor _21717_ (_13381_, _13380_, _11695_);
  or _21718_ (_13382_, _13381_, _07437_);
  or _21719_ (_13383_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _21720_ (_13384_, _13383_, _11510_);
  and _21721_ (_13385_, _13384_, _13382_);
  and _21722_ (_13386_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _21723_ (_13387_, _13386_, _13385_);
  and _21724_ (_12157_, _13387_, _05110_);
  nand _21725_ (_13388_, _13179_, _06088_);
  and _21726_ (_13389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _21727_ (_13390_, _13389_, _13197_);
  and _21728_ (_13391_, _13390_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _21729_ (_13392_, _13391_, _13193_);
  and _21730_ (_13393_, _13392_, _13356_);
  and _21731_ (_13394_, _13282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _21732_ (_13395_, _13394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _21733_ (_13396_, _13395_, _13193_);
  and _21734_ (_13397_, _13396_, _13177_);
  nor _21735_ (_13398_, _13397_, _13393_);
  or _21736_ (_13399_, _13398_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _21737_ (_13400_, _13398_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _21738_ (_13401_, _13400_, _13399_);
  nor _21739_ (_13402_, _13401_, _13179_);
  nor _21740_ (_13403_, _13402_, _13171_);
  and _21741_ (_13404_, _13403_, _13388_);
  and _21742_ (_13405_, _06062_, _05806_);
  and _21743_ (_13406_, _13405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _21744_ (_13407_, _13406_, _13404_);
  and _21745_ (_12161_, _13407_, _05110_);
  nand _21746_ (_13408_, _13179_, _06054_);
  and _21747_ (_13409_, _13197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _21748_ (_13410_, _13409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _21749_ (_13411_, _13410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _21750_ (_13412_, _13411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _21751_ (_13413_, _13412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _21752_ (_13414_, _13413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _21753_ (_13415_, _13414_, _13193_);
  and _21754_ (_13416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _21755_ (_13417_, _13416_, _13415_);
  or _21756_ (_13418_, _13417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not _21757_ (_13419_, _13177_);
  and _21758_ (_13420_, _13416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _21759_ (_13421_, _13420_, _13396_);
  nor _21760_ (_13422_, _13421_, _13419_);
  and _21761_ (_13423_, _13422_, _13418_);
  and _21762_ (_13424_, _13416_, _13393_);
  or _21763_ (_13425_, _13424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _21764_ (_13426_, _13420_, _13176_);
  nand _21765_ (_13427_, _13426_, _13392_);
  and _21766_ (_13428_, _13427_, _13419_);
  and _21767_ (_13429_, _13428_, _13425_);
  or _21768_ (_13430_, _13429_, _13423_);
  nor _21769_ (_13431_, _13430_, _13179_);
  nor _21770_ (_13432_, _13431_, _13171_);
  and _21771_ (_00002_, _13432_, _13408_);
  and _21772_ (_00003_, _13405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _21773_ (_00005_, _00003_, _00002_);
  and _21774_ (_12164_, _00005_, _05110_);
  nand _21775_ (_00006_, _13179_, _05334_);
  and _21776_ (_00007_, _13415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _21777_ (_00008_, _00007_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _21778_ (_00009_, _00008_, _13177_);
  nor _21779_ (_00010_, _00009_, _13417_);
  and _21780_ (_00011_, _13392_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _21781_ (_00012_, _00011_, _13176_);
  not _21782_ (_00013_, _00012_);
  nor _21783_ (_00014_, _00013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _21784_ (_00015_, _00013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _21785_ (_00016_, _00015_, _00014_);
  and _21786_ (_00017_, _00016_, _13419_);
  or _21787_ (_00019_, _00017_, _00010_);
  or _21788_ (_00020_, _00019_, _13179_);
  and _21789_ (_00021_, _00020_, _13371_);
  and _21790_ (_00022_, _00021_, _00006_);
  and _21791_ (_00023_, _13405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _21792_ (_00024_, _00023_, _00022_);
  and _21793_ (_12167_, _00024_, _05110_);
  or _21794_ (_00025_, _13373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _21795_ (_00026_, _00025_, _13398_);
  or _21796_ (_00027_, _00026_, _13179_);
  nand _21797_ (_00029_, _13179_, _06229_);
  nand _21798_ (_00030_, _00029_, _00027_);
  or _21799_ (_00032_, _00030_, _13405_);
  nand _21800_ (_00033_, _13405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _21801_ (_00034_, _00033_, _00032_);
  nor _21802_ (_12170_, _00034_, rst);
  and _21803_ (_00036_, _06473_, _05807_);
  not _21804_ (_00037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _21805_ (_00039_, t0_i);
  and _21806_ (_00040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _00039_);
  nor _21807_ (_00041_, _00040_, _00037_);
  not _21808_ (_00042_, _00041_);
  not _21809_ (_00043_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _21810_ (_00044_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor _21811_ (_00045_, _00044_, _00043_);
  and _21812_ (_00046_, _00045_, _00042_);
  not _21813_ (_00047_, _00046_);
  and _21814_ (_00048_, _11233_, _05804_);
  nor _21815_ (_00049_, _00048_, _00047_);
  or _21816_ (_00050_, _00049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _21817_ (_00051_, _00046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _21818_ (_00052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _21819_ (_00053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _21820_ (_00054_, _00053_, _00052_);
  and _21821_ (_00055_, _00054_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _21822_ (_00056_, _00055_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _21823_ (_00057_, _00056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _21824_ (_00058_, _00057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _21825_ (_00059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _21826_ (_00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _00059_);
  and _21827_ (_00061_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _21828_ (_00062_, _00061_, _00058_);
  nand _21829_ (_00063_, _00062_, _00051_);
  or _21830_ (_00064_, _00063_, _00048_);
  and _21831_ (_00065_, _00064_, _00050_);
  or _21832_ (_00066_, _00065_, _00036_);
  nand _21833_ (_00067_, _00036_, _06798_);
  and _21834_ (_00068_, _00067_, _05110_);
  and _21835_ (_12174_, _00068_, _00066_);
  not _21836_ (_00069_, _00048_);
  or _21837_ (_00070_, _00069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _21838_ (_00071_, _00051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _21839_ (_00072_, _00051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _21840_ (_00073_, _00072_, _00071_);
  and _21841_ (_00074_, _00058_, _00046_);
  and _21842_ (_00075_, _00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _21843_ (_00076_, _00075_, _00074_);
  or _21844_ (_00077_, _00076_, _00073_);
  or _21845_ (_00078_, _00077_, _00048_);
  and _21846_ (_00079_, _00078_, _00070_);
  or _21847_ (_00080_, _00079_, _00036_);
  nand _21848_ (_00081_, _00036_, _05938_);
  and _21849_ (_00082_, _00081_, _05110_);
  and _21850_ (_12191_, _00082_, _00080_);
  nand _21851_ (_00083_, _00036_, _06088_);
  and _21852_ (_00084_, _00054_, _00046_);
  not _21853_ (_00085_, _00084_);
  or _21854_ (_00086_, _00085_, _00048_);
  and _21855_ (_00087_, _00086_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _21856_ (_00088_, _00074_, _00060_);
  nand _21857_ (_00089_, _00088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _21858_ (_00090_, _00072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nand _21859_ (_00091_, _00090_, _00085_);
  and _21860_ (_00092_, _00091_, _00089_);
  nor _21861_ (_00093_, _00092_, _00048_);
  or _21862_ (_00094_, _00093_, _00087_);
  or _21863_ (_00095_, _00094_, _00036_);
  and _21864_ (_00096_, _00095_, _05110_);
  and _21865_ (_12196_, _00096_, _00083_);
  not _21866_ (_00097_, _00036_);
  or _21867_ (_00098_, _00069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _21868_ (_00099_, _00088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _21869_ (_00100_, _00072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor _21870_ (_00101_, _00100_, _00090_);
  or _21871_ (_00102_, _00101_, _00099_);
  or _21872_ (_00103_, _00102_, _00048_);
  and _21873_ (_00104_, _00103_, _00098_);
  and _21874_ (_00105_, _00104_, _00097_);
  nor _21875_ (_00106_, _00097_, _06229_);
  or _21876_ (_00107_, _00106_, _00105_);
  and _21877_ (_12199_, _00107_, _05110_);
  nor _21878_ (_00108_, _12744_, _12726_);
  nor _21879_ (_00109_, _00108_, _12745_);
  or _21880_ (_00110_, _00109_, _07437_);
  or _21881_ (_00111_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _21882_ (_00112_, _00111_, _12757_);
  and _21883_ (_00113_, _00112_, _00110_);
  and _21884_ (_00114_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _05110_);
  and _21885_ (_00115_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _21886_ (_12202_, _00115_, _00113_);
  nand _21887_ (_00116_, _08870_, _05334_);
  and _21888_ (_00117_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _21889_ (_00118_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _21890_ (_00119_, _00118_, _00117_);
  or _21891_ (_00120_, _00119_, _08870_);
  and _21892_ (_00121_, _00120_, _05110_);
  and _21893_ (_12206_, _00121_, _00116_);
  nand _21894_ (_00122_, _08870_, _05841_);
  and _21895_ (_00123_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _21896_ (_00124_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _21897_ (_00125_, _00124_, _00123_);
  or _21898_ (_00126_, _00125_, _08870_);
  and _21899_ (_00127_, _00126_, _05110_);
  and _21900_ (_12218_, _00127_, _00122_);
  not _21901_ (_00129_, _11219_);
  nor _21902_ (_00130_, _11711_, _00129_);
  and _21903_ (_00131_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _21904_ (_00132_, _00131_, _11223_);
  or _21905_ (_00133_, _00132_, _00130_);
  and _21906_ (_00134_, _00133_, _11202_);
  nor _21907_ (_00135_, _11711_, _12919_);
  or _21908_ (_00136_, _00135_, _11193_);
  or _21909_ (_00137_, _00136_, _00134_);
  nor _21910_ (_00138_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor _21911_ (_00139_, _00138_, _11234_);
  and _21912_ (_00140_, _00139_, _00137_);
  and _21913_ (_00141_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _21914_ (_00142_, _00141_, _11239_);
  or _21915_ (_00143_, _00142_, _00140_);
  nand _21916_ (_00144_, _11239_, _06088_);
  and _21917_ (_00145_, _00144_, _05110_);
  and _21918_ (_12226_, _00145_, _00143_);
  nand _21919_ (_00146_, _13179_, _05841_);
  not _21920_ (_00147_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _21921_ (_00148_, _13428_, _00147_);
  not _21922_ (_00149_, _00148_);
  nor _21923_ (_00150_, _00149_, _13422_);
  nor _21924_ (_00151_, _00150_, _00147_);
  and _21925_ (_00152_, _13177_, _00147_);
  and _21926_ (_00153_, _00152_, _13421_);
  nand _21927_ (_00154_, _13420_, _13393_);
  nor _21928_ (_00155_, _00154_, _00148_);
  or _21929_ (_00156_, _00155_, _00153_);
  or _21930_ (_00157_, _00156_, _00151_);
  or _21931_ (_00158_, _00157_, _13179_);
  and _21932_ (_00159_, _00158_, _13371_);
  and _21933_ (_00160_, _00159_, _00146_);
  and _21934_ (_00161_, _13250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _21935_ (_00162_, _00161_, _00160_);
  and _21936_ (_12238_, _00162_, _05110_);
  nand _21937_ (_00163_, _00036_, _06054_);
  and _21938_ (_00164_, _00084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _21939_ (_00165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nor _21940_ (_00166_, _00165_, _00048_);
  and _21941_ (_00167_, _00166_, _00164_);
  nand _21942_ (_00168_, _00167_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _21943_ (_00169_, _00167_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _21944_ (_00170_, _00169_, _00168_);
  nand _21945_ (_00171_, _00088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _21946_ (_00172_, _00171_, _00048_);
  or _21947_ (_00173_, _00172_, _00036_);
  or _21948_ (_00174_, _00173_, _00170_);
  and _21949_ (_00175_, _00174_, _05110_);
  and _21950_ (_12244_, _00175_, _00163_);
  nand _21951_ (_00176_, _00036_, _05841_);
  and _21952_ (_00177_, _00164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _21953_ (_00178_, _00177_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _21954_ (_00179_, _00057_, _00046_);
  nor _21955_ (_00180_, _00179_, _00165_);
  and _21956_ (_00181_, _00180_, _00178_);
  and _21957_ (_00182_, _00088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _21958_ (_00183_, _00182_, _00181_);
  nor _21959_ (_00184_, _00183_, _00048_);
  not _21960_ (_00185_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor _21961_ (_00186_, _00166_, _00185_);
  or _21962_ (_00187_, _00186_, _00184_);
  or _21963_ (_00188_, _00187_, _00036_);
  and _21964_ (_00189_, _00188_, _05110_);
  and _21965_ (_12247_, _00189_, _00176_);
  nand _21966_ (_00190_, _00036_, _05334_);
  nor _21967_ (_00191_, _00084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _21968_ (_00192_, _00191_, _00164_);
  and _21969_ (_00193_, _00088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _21970_ (_00194_, _00193_, _00192_);
  nor _21971_ (_00195_, _00194_, _00048_);
  and _21972_ (_00196_, _00048_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _21973_ (_00197_, _00196_, _00195_);
  or _21974_ (_00198_, _00197_, _00036_);
  and _21975_ (_00199_, _00198_, _05110_);
  and _21976_ (_12251_, _00199_, _00190_);
  and _21977_ (_00200_, _11326_, _08272_);
  nand _21978_ (_00201_, _00200_, _05872_);
  or _21979_ (_00202_, _00200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _21980_ (_00203_, _00202_, _11330_);
  and _21981_ (_00204_, _00203_, _00201_);
  nor _21982_ (_00205_, _11330_, _05938_);
  or _21983_ (_00206_, _00205_, _00204_);
  and _21984_ (_12261_, _00206_, _05110_);
  or _21985_ (_00207_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _21986_ (_00208_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _21987_ (_00209_, _00208_, _00207_);
  or _21988_ (_00210_, _00209_, _06895_);
  nand _21989_ (_00211_, _06895_, _05938_);
  and _21990_ (_00212_, _00211_, _05110_);
  and _21991_ (_12267_, _00212_, _00210_);
  or _21992_ (_00213_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand _21993_ (_00214_, _08884_, _11600_);
  and _21994_ (_00215_, _00214_, _00213_);
  or _21995_ (_00216_, _00215_, _06895_);
  nand _21996_ (_00217_, _06895_, _06798_);
  and _21997_ (_00218_, _00217_, _05110_);
  and _21998_ (_12271_, _00218_, _00216_);
  nor _21999_ (_00219_, _00069_, _05841_);
  and _22000_ (_00220_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _22001_ (_00221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _22002_ (_00222_, _00221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22003_ (_00223_, _00222_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _22004_ (_00224_, _00223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _22005_ (_00225_, _00224_, _00220_);
  and _22006_ (_00226_, _00225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22007_ (_00227_, _00226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _22008_ (_00228_, _00227_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _22009_ (_00229_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22010_ (_00230_, _00226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _22011_ (_00231_, _00230_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _22012_ (_00232_, _00231_, _00229_);
  and _22013_ (_00233_, _00224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22014_ (_00234_, _00233_, _00055_);
  and _22015_ (_00235_, _00234_, _00046_);
  or _22016_ (_00236_, _00235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _22017_ (_00237_, _00165_);
  and _22018_ (_00238_, _00235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _22019_ (_00239_, _00238_, _00237_);
  and _22020_ (_00240_, _00239_, _00236_);
  and _22021_ (_00241_, _00233_, _00074_);
  or _22022_ (_00242_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _22023_ (_00243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22024_ (_00244_, _00243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _22025_ (_00245_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _22026_ (_00246_, _00245_);
  and _22027_ (_00247_, _00246_, _00244_);
  and _22028_ (_00248_, _00247_, _00242_);
  or _22029_ (_00249_, _00248_, _00240_);
  or _22030_ (_00250_, _00249_, _00232_);
  and _22031_ (_00251_, _00250_, _00069_);
  or _22032_ (_00252_, _00251_, _00036_);
  or _22033_ (_00254_, _00252_, _00219_);
  or _22034_ (_00255_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _22035_ (_00256_, _00255_, _05110_);
  and _22036_ (_12293_, _00256_, _00254_);
  nand _22037_ (_00257_, _00048_, _06054_);
  and _22038_ (_00258_, _00074_, _00243_);
  and _22039_ (_00259_, _00258_, _00224_);
  nand _22040_ (_00260_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _22041_ (_00261_, _00244_, _00060_);
  or _22042_ (_00262_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22043_ (_00264_, _00262_, _00261_);
  and _22044_ (_00265_, _00264_, _00260_);
  or _22045_ (_00266_, _00225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22046_ (_00267_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not _22047_ (_00268_, _00226_);
  and _22048_ (_00269_, _00268_, _00267_);
  and _22049_ (_00270_, _00269_, _00266_);
  and _22050_ (_00271_, _00224_, _00164_);
  or _22051_ (_00272_, _00271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22052_ (_00274_, _00233_, _00164_);
  nor _22053_ (_00275_, _00274_, _00237_);
  and _22054_ (_00276_, _00275_, _00272_);
  or _22055_ (_00277_, _00276_, _00270_);
  or _22056_ (_00278_, _00277_, _00265_);
  or _22057_ (_00279_, _00278_, _00048_);
  and _22058_ (_00280_, _00279_, _00257_);
  or _22059_ (_00281_, _00280_, _00036_);
  or _22060_ (_00282_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _22061_ (_00283_, _00282_, _05110_);
  and _22062_ (_12296_, _00283_, _00281_);
  nand _22063_ (_00284_, _06890_, _05334_);
  and _22064_ (_00285_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _22065_ (_00286_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _22066_ (_00287_, _00286_, _00285_);
  or _22067_ (_00288_, _00287_, _06890_);
  and _22068_ (_00289_, _00288_, _08871_);
  and _22069_ (_00290_, _00289_, _00284_);
  and _22070_ (_00291_, _08870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _22071_ (_00292_, _00291_, _00290_);
  and _22072_ (_12299_, _00292_, _05110_);
  nand _22073_ (_00293_, _06890_, _06088_);
  and _22074_ (_00294_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _22075_ (_00295_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _22076_ (_00296_, _00295_, _00294_);
  or _22077_ (_00297_, _00296_, _06890_);
  and _22078_ (_00298_, _00297_, _08871_);
  and _22079_ (_00299_, _00298_, _00293_);
  and _22080_ (_00300_, _08870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _22081_ (_00301_, _00300_, _00299_);
  and _22082_ (_12302_, _00301_, _05110_);
  nand _22083_ (_00303_, _06890_, _06229_);
  and _22084_ (_00304_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _22085_ (_00305_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _22086_ (_00307_, _00305_, _00304_);
  or _22087_ (_00308_, _00307_, _06890_);
  and _22088_ (_00309_, _00308_, _08871_);
  and _22089_ (_00310_, _00309_, _00303_);
  and _22090_ (_00311_, _08870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _22091_ (_00312_, _00311_, _00310_);
  and _22092_ (_12306_, _00312_, _05110_);
  nand _22093_ (_00313_, _06890_, _05938_);
  or _22094_ (_00314_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _22095_ (_00315_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _22096_ (_00316_, _00315_, _00314_);
  or _22097_ (_00317_, _00316_, _06890_);
  and _22098_ (_00318_, _00317_, _08871_);
  and _22099_ (_00319_, _00318_, _00313_);
  and _22100_ (_00320_, _08870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _22101_ (_00321_, _00320_, _00319_);
  and _22102_ (_12309_, _00321_, _05110_);
  not _22103_ (_00322_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _22104_ (_00323_, _00258_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _22105_ (_00324_, _00323_, _00322_);
  nand _22106_ (_00325_, _00258_, _00221_);
  and _22107_ (_00326_, _00325_, _00261_);
  and _22108_ (_00327_, _00326_, _00324_);
  and _22109_ (_00328_, _00220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _22110_ (_00329_, _00328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _22111_ (_00330_, _00221_, _00220_);
  not _22112_ (_00331_, _00330_);
  and _22113_ (_00332_, _00331_, _00267_);
  and _22114_ (_00333_, _00332_, _00329_);
  nand _22115_ (_00334_, _00164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _22116_ (_00335_, _00334_, _00322_);
  and _22117_ (_00336_, _00221_, _00164_);
  nor _22118_ (_00337_, _00336_, _00237_);
  and _22119_ (_00338_, _00337_, _00335_);
  or _22120_ (_00339_, _00338_, _00333_);
  or _22121_ (_00340_, _00339_, _00327_);
  or _22122_ (_00341_, _00340_, _00048_);
  nand _22123_ (_00342_, _00048_, _05938_);
  and _22124_ (_00343_, _00342_, _00341_);
  or _22125_ (_00344_, _00343_, _00036_);
  nand _22126_ (_00345_, _00036_, _00322_);
  and _22127_ (_00346_, _00345_, _05110_);
  and _22128_ (_12317_, _00346_, _00344_);
  nand _22129_ (_00347_, _00048_, _06229_);
  or _22130_ (_00348_, _00336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22131_ (_00349_, _00222_, _00164_);
  nor _22132_ (_00350_, _00349_, _00237_);
  and _22133_ (_00351_, _00350_, _00348_);
  and _22134_ (_00352_, _00221_, _00074_);
  or _22135_ (_00353_, _00352_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _22136_ (_00354_, _00222_, _00074_);
  and _22137_ (_00355_, _00354_, _00244_);
  and _22138_ (_00356_, _00355_, _00353_);
  and _22139_ (_00357_, _00222_, _00220_);
  nand _22140_ (_00358_, _00357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _22141_ (_00359_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _22142_ (_00360_, _00359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22143_ (_00361_, _00360_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22144_ (_00362_, _00361_, _00358_);
  or _22145_ (_00363_, _00362_, _00356_);
  or _22146_ (_00364_, _00363_, _00351_);
  or _22147_ (_00365_, _00364_, _00048_);
  and _22148_ (_00366_, _00365_, _00347_);
  or _22149_ (_00367_, _00366_, _00036_);
  or _22150_ (_00368_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _22151_ (_00369_, _00368_, _05110_);
  and _22152_ (_12320_, _00369_, _00367_);
  nand _22153_ (_00370_, _00048_, _06088_);
  and _22154_ (_00371_, _00258_, _00222_);
  or _22155_ (_00372_, _00371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _22156_ (_00373_, _00371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _22157_ (_00374_, _00373_);
  and _22158_ (_00375_, _00374_, _00261_);
  and _22159_ (_00376_, _00375_, _00372_);
  and _22160_ (_00378_, _00223_, _00220_);
  or _22161_ (_00379_, _00357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _22162_ (_00380_, _00379_, _00267_);
  nor _22163_ (_00381_, _00380_, _00378_);
  or _22164_ (_00382_, _00349_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _22165_ (_00384_, _00223_, _00164_);
  nor _22166_ (_00386_, _00384_, _00237_);
  and _22167_ (_00388_, _00386_, _00382_);
  or _22168_ (_00389_, _00388_, _00381_);
  or _22169_ (_00390_, _00389_, _00376_);
  or _22170_ (_00391_, _00390_, _00048_);
  and _22171_ (_00392_, _00391_, _00370_);
  or _22172_ (_00393_, _00392_, _00036_);
  or _22173_ (_00394_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _22174_ (_00396_, _00394_, _05110_);
  and _22175_ (_12331_, _00396_, _00393_);
  nand _22176_ (_00397_, _00048_, _05334_);
  or _22177_ (_00398_, _00373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not _22178_ (_00400_, _00259_);
  and _22179_ (_00401_, _00400_, _00261_);
  and _22180_ (_00402_, _00401_, _00398_);
  not _22181_ (_00403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _22182_ (_00404_, _00378_, _00403_);
  and _22183_ (_00405_, _00378_, _00403_);
  or _22184_ (_00406_, _00405_, _00404_);
  and _22185_ (_00407_, _00406_, _00267_);
  or _22186_ (_00408_, _00384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _22187_ (_00409_, _00271_, _00237_);
  and _22188_ (_00410_, _00409_, _00408_);
  or _22189_ (_00412_, _00410_, _00407_);
  or _22190_ (_00413_, _00412_, _00402_);
  or _22191_ (_00414_, _00413_, _00048_);
  and _22192_ (_00416_, _00414_, _00397_);
  or _22193_ (_00418_, _00416_, _00036_);
  nand _22194_ (_00420_, _00036_, _00403_);
  and _22195_ (_00421_, _00420_, _05110_);
  and _22196_ (_12335_, _00421_, _00418_);
  nand _22197_ (_00423_, _06890_, _05841_);
  and _22198_ (_00424_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _22199_ (_00425_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _22200_ (_00426_, _00425_, _00424_);
  or _22201_ (_00427_, _00426_, _06890_);
  and _22202_ (_00428_, _00427_, _08871_);
  and _22203_ (_00429_, _00428_, _00423_);
  and _22204_ (_00430_, _06895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _22205_ (_00431_, _00430_, _00429_);
  and _22206_ (_12342_, _00431_, _05110_);
  or _22207_ (_00432_, _00258_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _22208_ (_00433_, _00323_, _00261_);
  and _22209_ (_00434_, _00433_, _00432_);
  or _22210_ (_00435_, _00220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  not _22211_ (_00436_, _00328_);
  and _22212_ (_00437_, _00436_, _00267_);
  and _22213_ (_00438_, _00437_, _00435_);
  or _22214_ (_00439_, _00164_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _22215_ (_00440_, _00334_, _00165_);
  and _22216_ (_00441_, _00440_, _00439_);
  or _22217_ (_00442_, _00441_, _00438_);
  or _22218_ (_00443_, _00442_, _00434_);
  or _22219_ (_00444_, _00443_, _00048_);
  nand _22220_ (_00445_, _00048_, _06798_);
  and _22221_ (_00446_, _00445_, _00444_);
  or _22222_ (_00447_, _00446_, _00036_);
  not _22223_ (_00448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _22224_ (_00449_, _00036_, _00448_);
  and _22225_ (_00450_, _00449_, _05110_);
  and _22226_ (_12348_, _00450_, _00447_);
  and _22227_ (_00452_, _08273_, _05804_);
  nor _22228_ (_00453_, _00452_, _00059_);
  and _22229_ (_00454_, _00452_, _06799_);
  or _22230_ (_00455_, _00454_, _00453_);
  and _22231_ (_12359_, _00455_, _05110_);
  nand _22232_ (_00456_, _00452_, _06229_);
  or _22233_ (_00457_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _22234_ (_00458_, _00457_, _05110_);
  and _22235_ (_12366_, _00458_, _00456_);
  nand _22236_ (_00459_, _00452_, _06088_);
  or _22237_ (_00460_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _22238_ (_00461_, _00460_, _05110_);
  and _22239_ (_12372_, _00461_, _00459_);
  nand _22240_ (_00463_, _00452_, _05938_);
  or _22241_ (_00464_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _22242_ (_00465_, _00464_, _05110_);
  and _22243_ (_12375_, _00465_, _00463_);
  nand _22244_ (_00466_, _00452_, _06054_);
  or _22245_ (_00468_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _22246_ (_00469_, _00468_, _05110_);
  and _22247_ (_12383_, _00469_, _00466_);
  nand _22248_ (_00470_, _00452_, _05841_);
  or _22249_ (_00471_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _22250_ (_00473_, _00471_, _05110_);
  and _22251_ (_12388_, _00473_, _00470_);
  nand _22252_ (_00474_, _00452_, _05334_);
  or _22253_ (_00475_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _22254_ (_00476_, _00475_, _05110_);
  and _22255_ (_12391_, _00476_, _00474_);
  nand _22256_ (_00477_, _08276_, _05901_);
  or _22257_ (_00478_, _08290_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  or _22258_ (_00479_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  and _22259_ (_00480_, _00479_, _00478_);
  or _22260_ (_00481_, _00480_, _08274_);
  and _22261_ (_00482_, _00481_, _05110_);
  and _22262_ (_12398_, _00482_, _00477_);
  and _22263_ (_12506_, _11775_, _05110_);
  and _22264_ (_00484_, _06856_, _06451_);
  not _22265_ (_00485_, _00484_);
  and _22266_ (_00486_, _06852_, _06446_);
  and _22267_ (_00487_, _00486_, _07062_);
  nor _22268_ (_00488_, _00487_, _06849_);
  and _22269_ (_00489_, _00488_, _00485_);
  or _22270_ (_12511_, _00489_, _06954_);
  and _22271_ (_00490_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _07601_);
  and _22272_ (_00491_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _22273_ (_00492_, _00491_, _00490_);
  and _22274_ (_12582_, _00492_, _05110_);
  nor _22275_ (_12593_, _12458_, rst);
  and _22276_ (_00493_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _07601_);
  and _22277_ (_00494_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _22278_ (_00495_, _00494_, _00493_);
  and _22279_ (_12600_, _00495_, _05110_);
  and _22280_ (_00496_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _05110_);
  and _22281_ (_00497_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _05110_);
  and _22282_ (_00498_, _00497_, _11506_);
  or _22283_ (_12644_, _00498_, _00496_);
  and _22284_ (_00499_, _11506_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _22285_ (_00500_, _00499_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _22286_ (_12685_, _00500_, _05110_);
  and _22287_ (_00501_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _07601_);
  and _22288_ (_00502_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _22289_ (_00503_, _00502_, _00501_);
  and _22290_ (_12721_, _00503_, _05110_);
  nor _22291_ (_12746_, _12505_, rst);
  and _22292_ (_12774_, _12029_, _05110_);
  and _22293_ (_12781_, _11890_, _05110_);
  nor _22294_ (_12840_, _11866_, rst);
  or _22295_ (_12842_, _12262_, rst);
  nand _22296_ (_12846_, _12193_, _05110_);
  nand _22297_ (_12852_, _12324_, _05110_);
  and _22298_ (_00504_, _06186_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _22299_ (_00505_, _06184_, _06559_);
  nand _22300_ (_00506_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor _22301_ (_00507_, _00506_, _06171_);
  or _22302_ (_00508_, _00507_, _00505_);
  or _22303_ (_00509_, _00508_, _00504_);
  and _22304_ (_12941_, _00509_, _05110_);
  nand _22305_ (_00510_, _08257_, _05938_);
  or _22306_ (_00511_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _22307_ (_00512_, _00511_, _05110_);
  and _22308_ (_12951_, _00512_, _00510_);
  and _22309_ (_00513_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not _22310_ (_00514_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _22311_ (_00515_, pc_log_change, _00514_);
  or _22312_ (_00516_, _00515_, _00513_);
  and _22313_ (_13022_, _00516_, _05110_);
  or _22314_ (_00517_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _22315_ (_00518_, pc_log_change, _05496_);
  and _22316_ (_00519_, _00518_, _05110_);
  and _22317_ (_13027_, _00519_, _00517_);
  and _22318_ (_13155_, _10472_, _11834_);
  and _22319_ (_00520_, _08615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _22320_ (_00521_, _07034_, _06169_);
  or _22321_ (_00522_, _00521_, _00520_);
  and _22322_ (_13169_, _00522_, _05110_);
  and _22323_ (_00523_, _10154_, _06626_);
  and _22324_ (_00524_, _00523_, _05488_);
  nand _22325_ (_00525_, _00524_, _05872_);
  or _22326_ (_00526_, _00524_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _22327_ (_00527_, _00526_, _05794_);
  and _22328_ (_00528_, _00527_, _00525_);
  not _22329_ (_00529_, _05793_);
  and _22330_ (_00530_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _22331_ (_00531_, _00523_, _05805_);
  nand _22332_ (_00532_, _00531_, _06780_);
  or _22333_ (_00533_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _22334_ (_00534_, _00533_, _05806_);
  and _22335_ (_00535_, _00534_, _00532_);
  or _22336_ (_00536_, _00535_, _00530_);
  or _22337_ (_00537_, _00536_, _00528_);
  and _22338_ (_13293_, _00537_, _05110_);
  and _22339_ (_00538_, _00523_, _08133_);
  nand _22340_ (_00539_, _00538_, _05872_);
  or _22341_ (_00540_, _00538_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _22342_ (_00541_, _00540_, _05794_);
  and _22343_ (_00542_, _00541_, _00539_);
  and _22344_ (_00543_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _22345_ (_00544_, _00531_, _06548_);
  or _22346_ (_00545_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _22347_ (_00546_, _00545_, _05806_);
  and _22348_ (_00547_, _00546_, _00544_);
  or _22349_ (_00548_, _00547_, _00543_);
  or _22350_ (_00549_, _00548_, _00542_);
  and _22351_ (_13307_, _00549_, _05110_);
  not _22352_ (_00550_, _00531_);
  or _22353_ (_00551_, _00550_, _05782_);
  or _22354_ (_00552_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _22355_ (_00553_, _00552_, _05794_);
  and _22356_ (_00554_, _00553_, _00551_);
  and _22357_ (_00555_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _22358_ (_00556_, _00531_, _07418_);
  and _22359_ (_00557_, _00556_, _05806_);
  and _22360_ (_00558_, _00557_, _00552_);
  or _22361_ (_00559_, _00558_, _00555_);
  or _22362_ (_00560_, _00559_, _00554_);
  and _22363_ (_13347_, _00560_, _05110_);
  and _22364_ (_00561_, _00523_, _06632_);
  nand _22365_ (_00562_, _00523_, _05401_);
  or _22366_ (_00563_, _00562_, _11548_);
  and _22367_ (_00564_, _00563_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _22368_ (_00565_, _00564_, _00561_);
  and _22369_ (_00566_, _00565_, _05794_);
  and _22370_ (_00567_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _22371_ (_00568_, _00531_, _06668_);
  or _22372_ (_00569_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _22373_ (_00570_, _00569_, _05806_);
  and _22374_ (_00571_, _00570_, _00568_);
  or _22375_ (_00572_, _00571_, _00567_);
  or _22376_ (_00573_, _00572_, _00566_);
  and _22377_ (_13357_, _00573_, _05110_);
  nand _22378_ (_00574_, _00523_, _11559_);
  and _22379_ (_00575_, _00574_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _22380_ (_00576_, _06173_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _22381_ (_00577_, _00576_, _08245_);
  and _22382_ (_00578_, _00577_, _00523_);
  or _22383_ (_00579_, _00578_, _00575_);
  and _22384_ (_00580_, _00579_, _05794_);
  and _22385_ (_00581_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _22386_ (_00582_, _00550_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nor _22387_ (_00583_, _00550_, _07337_);
  or _22388_ (_00584_, _00583_, _00582_);
  and _22389_ (_00585_, _00584_, _05806_);
  or _22390_ (_00586_, _00585_, _00581_);
  or _22391_ (_00587_, _00586_, _00580_);
  and _22392_ (_13360_, _00587_, _05110_);
  or _22393_ (_00588_, _12745_, _12723_);
  nor _22394_ (_00589_, _12747_, _07437_);
  and _22395_ (_00591_, _00589_, _00588_);
  nor _22396_ (_00592_, _07436_, _05195_);
  or _22397_ (_00593_, _00592_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _22398_ (_00594_, _00593_, _00591_);
  or _22399_ (_00595_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _11510_);
  and _22400_ (_00596_, _00595_, _05110_);
  and _22401_ (_00004_, _00596_, _00594_);
  and _22402_ (_00597_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor _22403_ (_00598_, _06088_, _06000_);
  and _22404_ (_00599_, _06011_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or _22405_ (_00600_, _00599_, _00598_);
  and _22406_ (_00601_, _00600_, _05337_);
  or _22407_ (_00602_, _00601_, _00597_);
  and _22408_ (_00018_, _00602_, _05110_);
  nand _22409_ (_00603_, _12750_, _12715_);
  and _22410_ (_00604_, _00603_, _12751_);
  or _22411_ (_00605_, _00604_, _07437_);
  or _22412_ (_00606_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _22413_ (_00607_, _00606_, _12757_);
  and _22414_ (_00608_, _00607_, _00605_);
  and _22415_ (_00609_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _22416_ (_00028_, _00609_, _00608_);
  nand _22417_ (_00610_, _08257_, _06798_);
  or _22418_ (_00611_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _22419_ (_00612_, _00611_, _05110_);
  and _22420_ (_00031_, _00612_, _00610_);
  or _22421_ (_00613_, _12749_, _12717_);
  and _22422_ (_00614_, _00613_, _12750_);
  or _22423_ (_00615_, _00614_, _07437_);
  or _22424_ (_00616_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _22425_ (_00617_, _00616_, _12757_);
  and _22426_ (_00618_, _00617_, _00615_);
  and _22427_ (_00619_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _22428_ (_00035_, _00619_, _00618_);
  and _22429_ (_00620_, _12748_, _12719_);
  nor _22430_ (_00621_, _00620_, _12749_);
  or _22431_ (_00622_, _00621_, _07437_);
  or _22432_ (_00623_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _22433_ (_00624_, _00623_, _12757_);
  and _22434_ (_00625_, _00624_, _00622_);
  and _22435_ (_00626_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _22436_ (_00038_, _00626_, _00625_);
  or _22437_ (_00627_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _22438_ (_00628_, _00627_, _05110_);
  nand _22439_ (_00629_, _08257_, _06088_);
  and _22440_ (_00128_, _00629_, _00628_);
  nor _22441_ (_00630_, _11681_, _11481_);
  nor _22442_ (_00631_, _00630_, _11682_);
  or _22443_ (_00632_, _00631_, _07437_);
  or _22444_ (_00633_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _22445_ (_00634_, _00633_, _12757_);
  and _22446_ (_00635_, _00634_, _00632_);
  and _22447_ (_00636_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _22448_ (_00253_, _00636_, _00635_);
  nand _22449_ (_00637_, _08257_, _06229_);
  or _22450_ (_00638_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _22451_ (_00639_, _00638_, _05110_);
  and _22452_ (_00263_, _00639_, _00637_);
  nor _22453_ (_00640_, _11689_, _11673_);
  nor _22454_ (_00641_, _00640_, _11690_);
  or _22455_ (_00642_, _00641_, _07437_);
  or _22456_ (_00643_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _22457_ (_00644_, _00643_, _12757_);
  and _22458_ (_00645_, _00644_, _00642_);
  and _22459_ (_00646_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _22460_ (_00273_, _00646_, _00645_);
  or _22461_ (_00647_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _11510_);
  and _22462_ (_00649_, _00647_, _05110_);
  or _22463_ (_00650_, _11688_, _11686_);
  nor _22464_ (_00651_, _11689_, _07437_);
  and _22465_ (_00652_, _00651_, _00650_);
  nor _22466_ (_00653_, _07436_, _05220_);
  or _22467_ (_00654_, _00653_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _22468_ (_00655_, _00654_, _00652_);
  and _22469_ (_00302_, _00655_, _00649_);
  nor _22470_ (_00656_, _11684_, _11682_);
  nor _22471_ (_00657_, _00656_, _11685_);
  or _22472_ (_00658_, _00657_, _07437_);
  or _22473_ (_00659_, _07436_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _22474_ (_00660_, _00659_, _12757_);
  and _22475_ (_00661_, _00660_, _00658_);
  and _22476_ (_00662_, _00114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _22477_ (_00306_, _00662_, _00661_);
  and _22478_ (_00663_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _22479_ (_00664_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _22480_ (_00665_, pc_log_change, _00664_);
  or _22481_ (_00666_, _00665_, _00663_);
  and _22482_ (_00377_, _00666_, _05110_);
  and _22483_ (_00667_, _00047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and _22484_ (_00668_, _00245_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _22485_ (_00669_, _00668_, _00667_);
  and _22486_ (_00670_, _00669_, _00244_);
  and _22487_ (_00671_, _00238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _22488_ (_00672_, _00671_, _00667_);
  and _22489_ (_00673_, _00672_, _00165_);
  or _22490_ (_00674_, _00667_, _00074_);
  and _22491_ (_00675_, _00674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _22492_ (_00676_, _00675_, _00673_);
  or _22493_ (_00677_, _00676_, _00670_);
  nor _22494_ (_00678_, _00036_, rst);
  and _22495_ (_00679_, _00678_, _00069_);
  and _22496_ (_00383_, _00679_, _00677_);
  nand _22497_ (_00680_, _00048_, _05901_);
  and _22498_ (_00681_, _00245_, _00243_);
  or _22499_ (_00682_, _00681_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _22500_ (_00683_, _00681_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _22501_ (_00684_, _00683_, _00682_);
  and _22502_ (_00685_, _00684_, _00261_);
  nand _22503_ (_00686_, _00230_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _22504_ (_00687_, _00230_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _22505_ (_00688_, _00687_, _00686_);
  and _22506_ (_00689_, _00688_, _00267_);
  or _22507_ (_00690_, _00238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _22508_ (_00691_, _00671_, _00237_);
  and _22509_ (_00692_, _00691_, _00690_);
  or _22510_ (_00693_, _00692_, _00689_);
  or _22511_ (_00694_, _00693_, _00685_);
  or _22512_ (_00695_, _00694_, _00048_);
  and _22513_ (_00696_, _00695_, _00680_);
  or _22514_ (_00697_, _00696_, _00036_);
  or _22515_ (_00698_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _22516_ (_00699_, _00698_, _05110_);
  and _22517_ (_00385_, _00699_, _00697_);
  and _22518_ (_00700_, _00166_, _00179_);
  or _22519_ (_00701_, _00700_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _22520_ (_00702_, _00243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _22521_ (_00703_, _00702_, _00059_);
  nand _22522_ (_00704_, _00703_, _00074_);
  or _22523_ (_00705_, _00704_, _00048_);
  and _22524_ (_00706_, _00705_, _00678_);
  and _22525_ (_00707_, _00706_, _00701_);
  nand _22526_ (_00708_, _00036_, _05110_);
  nor _22527_ (_00709_, _00708_, _05901_);
  or _22528_ (_00387_, _00709_, _00707_);
  nand _22529_ (_00710_, _00452_, _05901_);
  or _22530_ (_00711_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _22531_ (_00712_, _00711_, _05110_);
  and _22532_ (_00395_, _00712_, _00710_);
  not _22533_ (_00713_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _22534_ (_00714_, _00220_, _00713_);
  and _22535_ (_00715_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _22536_ (_00716_, _00715_, _00226_);
  or _22537_ (_00717_, _00716_, _00714_);
  and _22538_ (_00718_, _00717_, _00267_);
  and _22539_ (_00399_, _00718_, _00679_);
  and _22540_ (_00411_, t0_i, _05110_);
  nand _22541_ (_00719_, _13171_, _05901_);
  nor _22542_ (_00720_, _13202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _22543_ (_00721_, _00720_, _13251_);
  and _22544_ (_00722_, _00721_, _13180_);
  and _22545_ (_00723_, _13181_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nand _22546_ (_00724_, _13252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _22547_ (_00725_, _00724_, _13179_);
  or _22548_ (_00726_, _00725_, _00723_);
  or _22549_ (_00727_, _00726_, _00722_);
  or _22550_ (_00728_, _00727_, _13171_);
  and _22551_ (_00729_, _00728_, _05110_);
  and _22552_ (_00415_, _00729_, _00719_);
  not _22553_ (_00730_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _22554_ (_00731_, _13193_, _00730_);
  and _22555_ (_00732_, _13193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _22556_ (_00733_, _00732_, _13420_);
  and _22557_ (_00734_, _00733_, _13414_);
  and _22558_ (_00735_, _00734_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _22559_ (_00736_, _00735_, _00731_);
  and _22560_ (_00737_, _00736_, _13177_);
  and _22561_ (_00738_, _13420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _22562_ (_00739_, _00738_, _13391_);
  and _22563_ (_00740_, _00739_, _00732_);
  or _22564_ (_00741_, _00740_, _00731_);
  and _22565_ (_00742_, _00741_, _13356_);
  nand _22566_ (_00743_, _13193_, _13174_);
  and _22567_ (_00744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _22568_ (_00745_, _00744_, _00743_);
  or _22569_ (_00746_, _00745_, _13252_);
  or _22570_ (_00747_, _00746_, _00742_);
  or _22571_ (_00748_, _00747_, _00737_);
  nor _22572_ (_00749_, _13171_, _13179_);
  and _22573_ (_00750_, _00749_, _05110_);
  and _22574_ (_00417_, _00750_, _00748_);
  nand _22575_ (_00751_, _13179_, _05901_);
  not _22576_ (_00752_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _22577_ (_00753_, _00150_, _00752_);
  and _22578_ (_00754_, _00150_, _00752_);
  or _22579_ (_00755_, _00754_, _00753_);
  or _22580_ (_00756_, _00755_, _13179_);
  and _22581_ (_00757_, _00756_, _13371_);
  and _22582_ (_00758_, _00757_, _00751_);
  and _22583_ (_00759_, _13250_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _22584_ (_00760_, _00759_, _00758_);
  and _22585_ (_00419_, _00760_, _05110_);
  and _22586_ (_00422_, t1_i, _05110_);
  or _22587_ (_00761_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _22588_ (_00762_, _00761_, _05110_);
  nand _22589_ (_00763_, _08257_, _05841_);
  and _22590_ (_00451_, _00763_, _00762_);
  and _22591_ (_00764_, _12344_, _06745_);
  nor _22592_ (_00765_, _12392_, _06780_);
  not _22593_ (_00766_, _12067_);
  and _22594_ (_00768_, _12347_, _00766_);
  or _22595_ (_00770_, _12765_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _22596_ (_00771_, _00770_, _12766_);
  and _22597_ (_00772_, _00771_, _12374_);
  and _22598_ (_00773_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _22599_ (_00774_, _00773_, _00772_);
  or _22600_ (_00775_, _00774_, _00768_);
  or _22601_ (_00776_, _00775_, _00765_);
  nor _22602_ (_00777_, _00776_, _00764_);
  nand _22603_ (_00778_, _00777_, _12343_);
  nand _22604_ (_00779_, _12786_, _12404_);
  or _22605_ (_00780_, _12780_, _12404_);
  and _22606_ (_00781_, _00780_, _00779_);
  nor _22607_ (_00782_, _00781_, _05613_);
  and _22608_ (_00783_, _00781_, _05613_);
  or _22609_ (_00784_, _00783_, _00782_);
  and _22610_ (_00786_, _00784_, _13330_);
  or _22611_ (_00787_, _00786_, _00778_);
  nor _22612_ (_00788_, _12804_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _22613_ (_00789_, _00788_, _12805_);
  or _22614_ (_00790_, _00789_, _12343_);
  and _22615_ (_00791_, _00790_, _05110_);
  and _22616_ (_00462_, _00791_, _00787_);
  nor _22617_ (_00793_, _12785_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _22618_ (_00794_, _00793_, _00779_);
  nand _22619_ (_00795_, _12778_, _05123_);
  and _22620_ (_00797_, _00795_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _22621_ (_00798_, _00797_, _12780_);
  and _22622_ (_00799_, _00798_, _12403_);
  or _22623_ (_00800_, _00799_, _00794_);
  and _22624_ (_00801_, _00800_, _13330_);
  and _22625_ (_00802_, _12344_, _07277_);
  and _22626_ (_00803_, _12347_, _12417_);
  nor _22627_ (_00804_, _12392_, _06548_);
  nor _22628_ (_00805_, _12764_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _22629_ (_00806_, _00805_, _12765_);
  and _22630_ (_00807_, _00806_, _12374_);
  and _22631_ (_00808_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _22632_ (_00809_, _00808_, _00807_);
  or _22633_ (_00810_, _00809_, _00804_);
  or _22634_ (_00811_, _00810_, _00803_);
  nor _22635_ (_00812_, _00811_, _00802_);
  nand _22636_ (_00813_, _00812_, _12343_);
  or _22637_ (_00814_, _00813_, _00801_);
  nor _22638_ (_00815_, _12803_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _22639_ (_00816_, _00815_, _12804_);
  or _22640_ (_00817_, _00816_, _12343_);
  and _22641_ (_00818_, _00817_, _05110_);
  and _22642_ (_00467_, _00818_, _00814_);
  or _22643_ (_00819_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _22644_ (_00820_, _00819_, _05110_);
  nand _22645_ (_00821_, _08257_, _06054_);
  and _22646_ (_00472_, _00821_, _00820_);
  and _22647_ (_00822_, _12344_, _07204_);
  not _22648_ (_00823_, _07490_);
  and _22649_ (_00825_, _12347_, _00823_);
  and _22650_ (_00826_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _22651_ (_00827_, _12386_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _22652_ (_00828_, _00827_, _12764_);
  and _22653_ (_00829_, _00828_, _12374_);
  nor _22654_ (_00830_, _12392_, _07235_);
  or _22655_ (_00831_, _00830_, _00829_);
  or _22656_ (_00832_, _00831_, _00826_);
  or _22657_ (_00833_, _00832_, _00825_);
  nor _22658_ (_00834_, _00833_, _00822_);
  nand _22659_ (_00835_, _00834_, _12343_);
  and _22660_ (_00836_, _12784_, _12404_);
  and _22661_ (_00837_, _12778_, _12403_);
  nor _22662_ (_00838_, _00837_, _00836_);
  nand _22663_ (_00839_, _00838_, _05123_);
  or _22664_ (_00840_, _00838_, _05123_);
  and _22665_ (_00841_, _00840_, _00839_);
  and _22666_ (_00842_, _00841_, _12540_);
  or _22667_ (_00843_, _00842_, _00835_);
  nor _22668_ (_00844_, _12802_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _22669_ (_00845_, _00844_, _12803_);
  or _22670_ (_00846_, _00845_, _12343_);
  and _22671_ (_00847_, _00846_, _05110_);
  and _22672_ (_00483_, _00847_, _00843_);
  nor _22673_ (_00590_, _11787_, rst);
  and _22674_ (_00848_, _08614_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _22675_ (_00849_, _08617_, _06230_);
  nand _22676_ (_00850_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor _22677_ (_00851_, _00850_, _06004_);
  or _22678_ (_00852_, _00851_, _00849_);
  or _22679_ (_00853_, _00852_, _00848_);
  and _22680_ (_00648_, _00853_, _05110_);
  or _22681_ (_00854_, _12524_, _12522_);
  and _22682_ (_00855_, _13330_, _13332_);
  and _22683_ (_00856_, _00855_, _00854_);
  not _22684_ (_00857_, _12458_);
  and _22685_ (_00858_, _00857_, _12347_);
  not _22686_ (_00859_, _07235_);
  and _22687_ (_00860_, _13340_, _00859_);
  and _22688_ (_00861_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _22689_ (_00862_, _12374_, _00823_);
  or _22690_ (_00863_, _00862_, _00861_);
  or _22691_ (_00864_, _00863_, _00860_);
  or _22692_ (_00865_, _00864_, _00858_);
  or _22693_ (_00866_, _00865_, _00856_);
  and _22694_ (_00867_, _00866_, _12343_);
  nor _22695_ (_00868_, _07607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _22696_ (_00869_, _00868_, _12546_);
  nor _22697_ (_00870_, _00869_, _12343_);
  or _22698_ (_00872_, _00870_, _00867_);
  and _22699_ (_00767_, _00872_, _05110_);
  not _22700_ (_00873_, _12343_);
  or _22701_ (_00874_, _12471_, _12472_);
  not _22702_ (_00875_, _00874_);
  nand _22703_ (_00876_, _00875_, _12520_);
  or _22704_ (_00877_, _00875_, _12520_);
  and _22705_ (_00878_, _00877_, _13330_);
  and _22706_ (_00879_, _00878_, _00876_);
  not _22707_ (_00880_, _06668_);
  and _22708_ (_00881_, _13340_, _00880_);
  not _22709_ (_00882_, _07561_);
  and _22710_ (_00883_, _12347_, _00882_);
  and _22711_ (_00885_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _22712_ (_00886_, _12374_, _12346_);
  or _22713_ (_00887_, _00886_, _00885_);
  or _22714_ (_00888_, _00887_, _00883_);
  or _22715_ (_00889_, _00888_, _00881_);
  or _22716_ (_00890_, _00889_, _00879_);
  or _22717_ (_00891_, _00890_, _00873_);
  or _22718_ (_00892_, _12343_, _07609_);
  and _22719_ (_00893_, _00892_, _05110_);
  and _22720_ (_00769_, _00893_, _00891_);
  nand _22721_ (_00894_, _12374_, _12473_);
  or _22722_ (_00895_, _12518_, _12516_);
  nand _22723_ (_00896_, _00895_, _12540_);
  or _22724_ (_00897_, _00896_, _12519_);
  and _22725_ (_00898_, _12347_, _12475_);
  not _22726_ (_00899_, _07337_);
  and _22727_ (_00900_, _13340_, _00899_);
  and _22728_ (_00901_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _22729_ (_00902_, _00901_, _00900_);
  nor _22730_ (_00903_, _00902_, _00898_);
  and _22731_ (_00904_, _00903_, _00897_);
  nand _22732_ (_00905_, _00904_, _00894_);
  and _22733_ (_00906_, _00905_, _12343_);
  and _22734_ (_00907_, _00873_, _07620_);
  or _22735_ (_00908_, _00907_, _00906_);
  and _22736_ (_00785_, _00908_, _05110_);
  and _22737_ (_00909_, _12347_, _12482_);
  and _22738_ (_00910_, _12374_, _12480_);
  or _22739_ (_00911_, _00910_, _00909_);
  not _22740_ (_00912_, _06512_);
  and _22741_ (_00913_, _13340_, _00912_);
  and _22742_ (_00914_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _22743_ (_00916_, _00914_, _00913_);
  nor _22744_ (_00917_, _12513_, _12510_);
  nor _22745_ (_00918_, _00917_, _12514_);
  and _22746_ (_00919_, _00918_, _12540_);
  or _22747_ (_00920_, _00919_, _00916_);
  or _22748_ (_00922_, _00920_, _00911_);
  or _22749_ (_00923_, _00922_, _00873_);
  or _22750_ (_00924_, _12343_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _22751_ (_00925_, _00924_, _05110_);
  and _22752_ (_00792_, _00925_, _00923_);
  not _22753_ (_00926_, _07418_);
  and _22754_ (_00927_, _13340_, _00926_);
  and _22755_ (_00928_, _12507_, _12347_);
  and _22756_ (_00930_, _12374_, _12486_);
  and _22757_ (_00932_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _22758_ (_00934_, _00932_, _00930_);
  or _22759_ (_00935_, _00934_, _00928_);
  or _22760_ (_00936_, _00935_, _00927_);
  nor _22761_ (_00937_, _12509_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _22762_ (_00938_, _00937_, _12510_);
  and _22763_ (_00939_, _00938_, _12540_);
  or _22764_ (_00940_, _00939_, _00936_);
  or _22765_ (_00941_, _00940_, _00873_);
  or _22766_ (_00942_, _12343_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _22767_ (_00943_, _00942_, _05110_);
  and _22768_ (_00796_, _00943_, _00941_);
  and _22769_ (_00824_, _06411_, _05110_);
  and _22770_ (_00944_, _12344_, _07364_);
  and _22771_ (_00945_, _12374_, _11340_);
  and _22772_ (_00946_, _12347_, _12480_);
  and _22773_ (_00947_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _22774_ (_00948_, _12392_, _06512_);
  or _22775_ (_00949_, _00948_, _00947_);
  or _22776_ (_00950_, _00949_, _00946_);
  or _22777_ (_00951_, _00950_, _00945_);
  or _22778_ (_00952_, _00951_, _00944_);
  and _22779_ (_00953_, _12528_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _22780_ (_00954_, _00953_, _12403_);
  and _22781_ (_00955_, _12529_, _12403_);
  nor _22782_ (_00956_, _00955_, _00954_);
  or _22783_ (_00957_, _00956_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _22784_ (_00958_, _00956_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _22785_ (_00959_, _00958_, _00957_);
  and _22786_ (_00960_, _00959_, _12540_);
  nor _22787_ (_00961_, _00960_, _00952_);
  nand _22788_ (_00962_, _00961_, _12343_);
  nor _22789_ (_00963_, _12550_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _22790_ (_00964_, _00963_, _12551_);
  or _22791_ (_00965_, _00964_, _12343_);
  and _22792_ (_00966_, _00965_, _05110_);
  and _22793_ (_00871_, _00966_, _00962_);
  and _22794_ (_00967_, _12344_, _07391_);
  and _22795_ (_00968_, _12374_, _06909_);
  and _22796_ (_00969_, _12347_, _12486_);
  and _22797_ (_00970_, _12369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _22798_ (_00971_, _11309_, _00926_);
  or _22799_ (_00972_, _00971_, _00970_);
  or _22800_ (_00973_, _00972_, _00969_);
  or _22801_ (_00974_, _00973_, _00968_);
  or _22802_ (_00975_, _00974_, _00967_);
  nand _22803_ (_00976_, _12528_, _05240_);
  or _22804_ (_00977_, _12528_, _05240_);
  and _22805_ (_00978_, _00977_, _00976_);
  and _22806_ (_00979_, _00978_, _12403_);
  and _22807_ (_00980_, _00954_, _12529_);
  or _22808_ (_00981_, _00980_, _00979_);
  and _22809_ (_00982_, _00981_, _13330_);
  or _22810_ (_00983_, _00982_, _00975_);
  and _22811_ (_00984_, _00983_, _12343_);
  nor _22812_ (_00985_, _12549_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or _22813_ (_00986_, _00985_, _12550_);
  nor _22814_ (_00987_, _00986_, _12343_);
  or _22815_ (_00988_, _00987_, _00984_);
  and _22816_ (_00884_, _00988_, _05110_);
  and _22817_ (_00989_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not _22818_ (_00990_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor _22819_ (_00991_, pc_log_change, _00990_);
  or _22820_ (_00992_, _00991_, _00989_);
  and _22821_ (_00915_, _00992_, _05110_);
  and _22822_ (_00993_, _06904_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _22823_ (_00994_, _06901_, _12874_);
  or _22824_ (_00995_, _00994_, _00993_);
  and _22825_ (_00921_, _00995_, _05110_);
  or _22826_ (_00996_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _22827_ (_00997_, _00996_, _08243_);
  and _22828_ (_00998_, _05782_, _08272_);
  not _22829_ (_00999_, _08272_);
  nand _22830_ (_01000_, _00999_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _22831_ (_01002_, _01000_, _08243_);
  or _22832_ (_01003_, _01002_, _00998_);
  and _22833_ (_01004_, _01003_, _00997_);
  or _22834_ (_01005_, _01004_, _08253_);
  nand _22835_ (_01006_, _08253_, _05938_);
  and _22836_ (_01007_, _01006_, _05110_);
  and _22837_ (_00929_, _01007_, _01005_);
  and _22838_ (_01008_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _22839_ (_01009_, _07028_);
  and _22840_ (_01010_, _13340_, _01009_);
  not _22841_ (_01011_, _07176_);
  and _22842_ (_01012_, _12347_, _01011_);
  and _22843_ (_01013_, _12374_, _12762_);
  or _22844_ (_01014_, _01013_, _01012_);
  or _22845_ (_01015_, _01014_, _01010_);
  and _22846_ (_01016_, _12525_, _12522_);
  or _22847_ (_01017_, _01016_, _12465_);
  and _22848_ (_01018_, _01017_, _12415_);
  nor _22849_ (_01019_, _01018_, _12409_);
  nor _22850_ (_01020_, _01019_, _12411_);
  and _22851_ (_01021_, _01019_, _12411_);
  or _22852_ (_01022_, _01021_, _01020_);
  and _22853_ (_01023_, _01022_, _12540_);
  or _22854_ (_01024_, _01023_, _01015_);
  nor _22855_ (_01025_, _01024_, _01008_);
  nand _22856_ (_01026_, _01025_, _12343_);
  nor _22857_ (_01027_, _12548_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _22858_ (_01028_, _01027_, _12549_);
  or _22859_ (_01029_, _01028_, _12343_);
  and _22860_ (_01030_, _01029_, _05110_);
  and _22861_ (_00931_, _01030_, _01026_);
  not _22862_ (_01031_, _07582_);
  and _22863_ (_01032_, _12347_, _01031_);
  and _22864_ (_01033_, _12374_, _00766_);
  or _22865_ (_01034_, _01033_, _01032_);
  not _22866_ (_01035_, _06780_);
  and _22867_ (_01036_, _13340_, _01035_);
  and _22868_ (_01037_, _11309_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _22869_ (_01038_, _01037_, _01036_);
  nor _22870_ (_01039_, _01017_, _12415_);
  nor _22871_ (_01040_, _01039_, _01018_);
  and _22872_ (_01041_, _01040_, _12540_);
  or _22873_ (_01042_, _01041_, _01038_);
  or _22874_ (_01044_, _01042_, _01034_);
  and _22875_ (_01045_, _01044_, _12343_);
  nor _22876_ (_01046_, _12547_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _22877_ (_01047_, _01046_, _12548_);
  nor _22878_ (_01048_, _01047_, _12343_);
  or _22879_ (_01049_, _01048_, _01045_);
  and _22880_ (_00933_, _01049_, _05110_);
  not _22881_ (_01050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand _22882_ (_01051_, _01050_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _22883_ (_01052_, _01051_, _08235_);
  and _22884_ (_01053_, _01052_, _08237_);
  or _22885_ (_01054_, _01053_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _22886_ (_01055_, _01054_, _08243_);
  and _22887_ (_01056_, _05782_, _05805_);
  not _22888_ (_01057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _22889_ (_01058_, _05805_, _01057_);
  nand _22890_ (_01059_, _01058_, _08243_);
  or _22891_ (_01060_, _01059_, _01056_);
  and _22892_ (_01061_, _01060_, _01055_);
  or _22893_ (_01062_, _01061_, _08253_);
  nand _22894_ (_01063_, _08253_, _06798_);
  and _22895_ (_01064_, _01063_, _05110_);
  and _22896_ (_01043_, _01064_, _01062_);
  and _22897_ (_01065_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _22898_ (_01066_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _22899_ (_01447_, _01066_, _01065_);
  not _22900_ (_01067_, _08243_);
  or _22901_ (_01068_, _10212_, _01067_);
  and _22902_ (_01069_, _01068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _22903_ (_01070_, _01069_, _08253_);
  and _22904_ (_01071_, _10178_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _22905_ (_01072_, _01071_, _10209_);
  and _22906_ (_01073_, _01072_, _08243_);
  or _22907_ (_01074_, _01073_, _01070_);
  nand _22908_ (_01075_, _08253_, _05334_);
  and _22909_ (_01076_, _01075_, _05110_);
  and _22910_ (_01453_, _01076_, _01074_);
  and _22911_ (_01077_, _05795_, _05419_);
  and _22912_ (_01078_, _01077_, _05460_);
  and _22913_ (_01079_, _01078_, _06122_);
  not _22914_ (_01080_, _01079_);
  or _22915_ (_01081_, _10212_, _01080_);
  and _22916_ (_01082_, _01081_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _22917_ (_01083_, _01082_, _06148_);
  and _22918_ (_01084_, _10178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _22919_ (_01085_, _01084_, _10209_);
  and _22920_ (_01086_, _01085_, _06153_);
  or _22921_ (_01087_, _01086_, _01083_);
  nand _22922_ (_01088_, _06148_, _05334_);
  and _22923_ (_01089_, _01088_, _05110_);
  and _22924_ (_01459_, _01089_, _01087_);
  and _22925_ (_01090_, _06153_, _08272_);
  or _22926_ (_01091_, _01090_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _22927_ (_01092_, _01091_, _06149_);
  nand _22928_ (_01093_, _01090_, _05872_);
  and _22929_ (_01094_, _01093_, _01092_);
  nor _22930_ (_01095_, _06149_, _05938_);
  or _22931_ (_01096_, _01095_, _01094_);
  and _22932_ (_01460_, _01096_, _05110_);
  and _22933_ (_01097_, _10178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _22934_ (_01098_, _01097_, _10209_);
  and _22935_ (_01099_, _01098_, _06123_);
  not _22936_ (_01100_, _06123_);
  or _22937_ (_01101_, _10212_, _01100_);
  and _22938_ (_01102_, _01101_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _22939_ (_01103_, _01102_, _06129_);
  or _22940_ (_01104_, _01103_, _01099_);
  nand _22941_ (_01105_, _06129_, _05334_);
  and _22942_ (_01106_, _01105_, _05110_);
  and _22943_ (_01463_, _01106_, _01104_);
  and _22944_ (_01107_, _06123_, _08272_);
  nand _22945_ (_01108_, _01107_, _05872_);
  or _22946_ (_01109_, _01107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _22947_ (_01110_, _01109_, _06130_);
  and _22948_ (_01111_, _01110_, _01108_);
  nor _22949_ (_01112_, _06130_, _05938_);
  or _22950_ (_01113_, _01112_, _01111_);
  and _22951_ (_01465_, _01113_, _05110_);
  nand _22952_ (_01114_, _08243_, _05401_);
  and _22953_ (_01115_, _01114_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _22954_ (_01116_, _01115_, _08253_);
  and _22955_ (_01117_, _11559_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _22956_ (_01118_, _01117_, _06632_);
  and _22957_ (_01119_, _01118_, _08243_);
  or _22958_ (_01120_, _01119_, _01116_);
  nand _22959_ (_01121_, _08253_, _06088_);
  and _22960_ (_01122_, _01121_, _05110_);
  and _22961_ (_01468_, _01122_, _01120_);
  nor _22962_ (_01123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _22963_ (_01124_, _01123_, _05976_);
  nor _22964_ (_01125_, _01124_, _06105_);
  nand _22965_ (_01126_, _05980_, _05860_);
  not _22966_ (_01127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nand _22967_ (_01128_, _05973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _22968_ (_01129_, _01128_, _01127_);
  nor _22969_ (_01130_, _05972_, _05850_);
  or _22970_ (_01131_, _01130_, _05980_);
  or _22971_ (_01132_, _01131_, _01129_);
  and _22972_ (_01133_, _01132_, _06104_);
  and _22973_ (_01134_, _01133_, _01126_);
  or _22974_ (_01135_, _01134_, _01125_);
  nand _22975_ (_01136_, _05976_, _05860_);
  and _22976_ (_01137_, _01136_, _01135_);
  nand _22977_ (_01138_, _01137_, _06099_);
  not _22978_ (_01139_, _05971_);
  nor _22979_ (_01140_, _06099_, _01139_);
  nand _22980_ (_01141_, _01140_, _01127_);
  nor _22981_ (_01142_, _01123_, _05967_);
  and _22982_ (_01143_, _05946_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _22983_ (_01144_, _01143_, _05955_);
  and _22984_ (_01145_, _05951_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _22985_ (_01146_, _01145_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _22986_ (_01147_, _01146_, _05967_);
  and _22987_ (_01148_, _01147_, _01144_);
  or _22988_ (_01149_, _01148_, _01142_);
  and _22989_ (_01150_, _01149_, _05960_);
  and _22990_ (_01151_, _05967_, _05955_);
  or _22991_ (_01152_, _01151_, _05959_);
  nand _22992_ (_01153_, _01152_, _05860_);
  nand _22993_ (_01154_, _01153_, _06100_);
  or _22994_ (_01155_, _01154_, _01150_);
  and _22995_ (_01156_, _01155_, _01141_);
  and _22996_ (_01157_, _01156_, _01138_);
  or _22997_ (_01158_, _01157_, _05986_);
  nand _22998_ (_01159_, _05986_, _01127_);
  and _22999_ (_01160_, _01159_, _05110_);
  and _23000_ (_01471_, _01160_, _01158_);
  nand _23001_ (_01161_, _01140_, _06092_);
  nor _23002_ (_01162_, _05986_, _06099_);
  or _23003_ (_01163_, _01162_, _05850_);
  and _23004_ (_01164_, _01163_, _05110_);
  and _23005_ (_01475_, _01164_, _01161_);
  nand _23006_ (_01165_, _05969_, _06110_);
  nor _23007_ (_01166_, _01165_, _06099_);
  and _23008_ (_01167_, _05986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  not _23009_ (_01168_, _05982_);
  or _23010_ (_01169_, _06098_, _01168_);
  nor _23011_ (_01170_, _01169_, _05975_);
  and _23012_ (_01171_, _01170_, _06137_);
  or _23013_ (_01172_, _01171_, _01167_);
  or _23014_ (_01173_, _01172_, _01166_);
  and _23015_ (_01478_, _01173_, _05110_);
  and _23016_ (_01479_, _13167_, _05986_);
  and _23017_ (_01174_, _06625_, _05789_);
  and _23018_ (_01175_, _01174_, _05867_);
  nand _23019_ (_01176_, _01175_, _05872_);
  or _23020_ (_01177_, _01175_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _23021_ (_01178_, _01177_, _05794_);
  and _23022_ (_01179_, _01178_, _01176_);
  and _23023_ (_01180_, _05804_, _05992_);
  nand _23024_ (_01181_, _01180_, _05901_);
  or _23025_ (_01182_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _23026_ (_01183_, _01182_, _05806_);
  and _23027_ (_01184_, _01183_, _01181_);
  and _23028_ (_01185_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _23029_ (_01186_, _01185_, rst);
  or _23030_ (_01187_, _01186_, _01184_);
  or _23031_ (_01488_, _01187_, _01179_);
  and _23032_ (_01188_, _06153_, _08133_);
  or _23033_ (_01189_, _01188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _23034_ (_01190_, _01189_, _06149_);
  nand _23035_ (_01191_, _01188_, _05872_);
  and _23036_ (_01192_, _01191_, _01190_);
  nor _23037_ (_01193_, _06149_, _06054_);
  or _23038_ (_01194_, _01193_, _01192_);
  and _23039_ (_01494_, _01194_, _05110_);
  and _23040_ (_01195_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _23041_ (_01196_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _23042_ (_01498_, _01196_, _01195_);
  and _23043_ (_01197_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and _23044_ (_01198_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or _23045_ (_01500_, _01198_, _01197_);
  and _23046_ (_01199_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _23047_ (_01200_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _23048_ (_01513_, _01200_, _01199_);
  and _23049_ (_01201_, _06123_, _08133_);
  nand _23050_ (_01202_, _01201_, _05872_);
  or _23051_ (_01203_, _01201_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _23052_ (_01204_, _01203_, _06130_);
  and _23053_ (_01205_, _01204_, _01202_);
  nor _23054_ (_01206_, _06130_, _06054_);
  or _23055_ (_01207_, _01206_, _01205_);
  and _23056_ (_01516_, _01207_, _05110_);
  and _23057_ (_01520_, _00496_, _05986_);
  and _23058_ (_01208_, _05798_, _05805_);
  or _23059_ (_01209_, _01208_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _23060_ (_01210_, _01209_, _05844_);
  nand _23061_ (_01211_, _01208_, _05872_);
  and _23062_ (_01212_, _01211_, _01210_);
  and _23063_ (_01213_, _06799_, _05809_);
  or _23064_ (_01214_, _01213_, _01212_);
  and _23065_ (_01522_, _01214_, _05110_);
  nor _23066_ (_01215_, _01140_, _05986_);
  not _23067_ (_01216_, _01215_);
  and _23068_ (_01217_, _01216_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _23069_ (_01218_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _23070_ (_01219_, _05973_, _05850_);
  or _23071_ (_01220_, _01219_, _01218_);
  nor _23072_ (_01221_, _05972_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23073_ (_01222_, _01221_, _05980_);
  nand _23074_ (_01223_, _01222_, _01220_);
  or _23075_ (_01224_, _06114_, _05849_);
  and _23076_ (_01225_, _01224_, _01223_);
  or _23077_ (_01226_, _01225_, _05979_);
  not _23078_ (_01227_, _05977_);
  not _23079_ (_01228_, _05979_);
  or _23080_ (_01229_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _05850_);
  or _23081_ (_01230_, _01229_, _01228_);
  and _23082_ (_01231_, _01230_, _01227_);
  and _23083_ (_01232_, _01231_, _01226_);
  and _23084_ (_01233_, _05977_, _05849_);
  or _23085_ (_01234_, _01233_, _05976_);
  or _23086_ (_01235_, _01234_, _01232_);
  or _23087_ (_01236_, _01229_, _06103_);
  and _23088_ (_01237_, _01236_, _06099_);
  and _23089_ (_01238_, _01237_, _01235_);
  and _23090_ (_01239_, _05951_, _05850_);
  or _23091_ (_01240_, _01239_, _01218_);
  and _23092_ (_01241_, _05946_, _05850_);
  nor _23093_ (_01242_, _01241_, _05955_);
  nand _23094_ (_01243_, _01242_, _01240_);
  or _23095_ (_01244_, _05956_, _05849_);
  and _23096_ (_01245_, _01244_, _01243_);
  or _23097_ (_01246_, _01245_, _05966_);
  not _23098_ (_01247_, _05963_);
  not _23099_ (_01248_, _05966_);
  or _23100_ (_01249_, _01229_, _01248_);
  and _23101_ (_01250_, _01249_, _01247_);
  and _23102_ (_01251_, _01250_, _01246_);
  and _23103_ (_01252_, _05963_, _05849_);
  or _23104_ (_01253_, _01252_, _05959_);
  or _23105_ (_01254_, _01253_, _01251_);
  and _23106_ (_01255_, _06100_, _05960_);
  and _23107_ (_01256_, _01229_, _06100_);
  or _23108_ (_01257_, _01256_, _01255_);
  and _23109_ (_01258_, _01257_, _01254_);
  or _23110_ (_01259_, _01258_, _01238_);
  and _23111_ (_01260_, _01259_, _06137_);
  or _23112_ (_01261_, _01260_, _01217_);
  and _23113_ (_01527_, _01261_, _05110_);
  and _23114_ (_01531_, _06388_, _05110_);
  nor _23115_ (_01262_, _05841_, _05465_);
  and _23116_ (_01263_, _05465_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or _23117_ (_01264_, _01263_, _01262_);
  and _23118_ (_01540_, _01264_, _05110_);
  and _23119_ (_01561_, _06366_, _05110_);
  and _23120_ (_01265_, _05798_, _10208_);
  or _23121_ (_01266_, _01265_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _23122_ (_01267_, _01266_, _05844_);
  nand _23123_ (_01268_, _01265_, _05872_);
  and _23124_ (_01269_, _01268_, _01267_);
  nor _23125_ (_01270_, _05844_, _05334_);
  or _23126_ (_01271_, _01270_, _01269_);
  and _23127_ (_01565_, _01271_, _05110_);
  and _23128_ (_01272_, _05798_, _06472_);
  nand _23129_ (_01273_, _01272_, _05872_);
  or _23130_ (_01274_, _01272_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _23131_ (_01275_, _01274_, _05844_);
  and _23132_ (_01276_, _01275_, _01273_);
  nor _23133_ (_01277_, _06229_, _05844_);
  or _23134_ (_01278_, _01277_, _01276_);
  and _23135_ (_01567_, _01278_, _05110_);
  and _23136_ (_01279_, _05986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _23137_ (_01280_, _01279_, _01215_);
  and _23138_ (_01571_, _01280_, _05110_);
  and _23139_ (_01281_, _05986_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _23140_ (_01282_, _01281_, _01215_);
  and _23141_ (_01574_, _01282_, _05110_);
  and _23142_ (_01283_, _08615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _23143_ (_01284_, _08617_, _12894_);
  or _23144_ (_01285_, _01284_, _01283_);
  and _23145_ (_01577_, _01285_, _05110_);
  or _23146_ (_01286_, _05966_, _05955_);
  and _23147_ (_01287_, _05952_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _23148_ (_01288_, _01287_, _01286_);
  and _23149_ (_01289_, _01288_, _01247_);
  and _23150_ (_01290_, _01289_, _01255_);
  nand _23151_ (_01291_, _05975_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nand _23152_ (_01292_, _01291_, _05981_);
  and _23153_ (_01293_, _01292_, _05978_);
  and _23154_ (_01294_, _01293_, _06099_);
  or _23155_ (_01295_, _01294_, _05986_);
  or _23156_ (_01296_, _01295_, _01290_);
  nand _23157_ (_01297_, _05986_, _11499_);
  and _23158_ (_01298_, _01297_, _05110_);
  and _23159_ (_01581_, _01298_, _01296_);
  nor _23160_ (_01299_, _05951_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _23161_ (_01300_, _01299_, _05946_);
  or _23162_ (_01301_, _01300_, _05955_);
  and _23163_ (_01302_, _01301_, _01248_);
  or _23164_ (_01303_, _01302_, _05963_);
  and _23165_ (_01304_, _01303_, _01255_);
  and _23166_ (_01305_, _06099_, _06103_);
  or _23167_ (_01306_, _05973_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _23168_ (_01307_, _01306_, _05972_);
  or _23169_ (_01308_, _01307_, _05980_);
  and _23170_ (_01309_, _01308_, _01228_);
  or _23171_ (_01310_, _01309_, _05977_);
  and _23172_ (_01311_, _01310_, _01305_);
  or _23173_ (_01312_, _01311_, _05986_);
  or _23174_ (_01313_, _01312_, _01304_);
  or _23175_ (_01314_, _06137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _23176_ (_01315_, _01314_, _05110_);
  and _23177_ (_01590_, _01315_, _01313_);
  nor _23178_ (_01316_, _11268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _23179_ (_01317_, _01316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _23180_ (_01318_, _01316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _23181_ (_01319_, _01318_, _05110_);
  and _23182_ (_01600_, _01319_, _01317_);
  not _23183_ (_01320_, _06560_);
  nor _23184_ (_01321_, _01320_, _05901_);
  and _23185_ (_01322_, _01320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or _23186_ (_01323_, _01322_, _01321_);
  and _23187_ (_01604_, _01323_, _05110_);
  and _23188_ (_01324_, _08750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not _23189_ (_01325_, _08745_);
  and _23190_ (_01326_, _08754_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor _23191_ (_01327_, _01326_, _01325_);
  or _23192_ (_01328_, _01327_, _01324_);
  and _23193_ (_01329_, _08754_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _23194_ (_01330_, _01329_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _23195_ (_01331_, _01330_, _05110_);
  and _23196_ (_01619_, _01331_, _01328_);
  or _23197_ (_01332_, _06984_, _07177_);
  nor _23198_ (_01333_, _07208_, _07028_);
  and _23199_ (_01334_, _07208_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _23200_ (_01335_, _01334_, _06471_);
  or _23201_ (_01336_, _01335_, _01333_);
  and _23202_ (_01337_, _01336_, _05110_);
  and _23203_ (_01636_, _01337_, _01332_);
  and _23204_ (_01338_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not _23205_ (_01339_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _23206_ (_01340_, pc_log_change, _01339_);
  or _23207_ (_01341_, _01340_, _01338_);
  and _23208_ (_01646_, _01341_, _05110_);
  nand _23209_ (_01342_, _07028_, _06477_);
  or _23210_ (_01343_, _06477_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _23211_ (_01344_, _01343_, _05110_);
  and _23212_ (_01669_, _01344_, _01342_);
  or _23213_ (_01345_, _05718_, _05716_);
  not _23214_ (_01346_, _05653_);
  nand _23215_ (_01347_, _05716_, _01346_);
  and _23216_ (_01348_, _01347_, _05650_);
  and _23217_ (_01349_, _01348_, _01345_);
  nand _23218_ (_01350_, _05646_, _05519_);
  and _23219_ (_01351_, _05647_, _05489_);
  and _23220_ (_01352_, _01351_, _01350_);
  and _23221_ (_01353_, _06485_, ABINPUT000000[0]);
  and _23222_ (_01354_, _06487_, ABINPUT000[0]);
  nor _23223_ (_01355_, _01354_, _01353_);
  nand _23224_ (_01356_, _01355_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _23225_ (_01357_, _01356_, _01352_);
  or _23226_ (_01358_, _01357_, _01349_);
  or _23227_ (_01359_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and _23228_ (_01360_, _01359_, _01358_);
  and _23229_ (_01361_, _01360_, _10211_);
  not _23230_ (_01362_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _23231_ (_01363_, _06472_, _01362_);
  or _23232_ (_01364_, _01363_, _08245_);
  and _23233_ (_01365_, _01364_, _10157_);
  nor _23234_ (_01366_, _01365_, _01361_);
  nand _23235_ (_01367_, _01366_, _10163_);
  nand _23236_ (_01368_, _10162_, _06229_);
  and _23237_ (_01369_, _01368_, _05110_);
  and _23238_ (_01741_, _01369_, _01367_);
  nor _23239_ (_01370_, _06054_, _06010_);
  and _23240_ (_01371_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _23241_ (_01372_, _01371_, _05995_);
  or _23242_ (_01373_, _01372_, _01370_);
  or _23243_ (_01374_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _23244_ (_01375_, _01374_, _05110_);
  and _23245_ (_01746_, _01375_, _01373_);
  or _23246_ (_01376_, _11202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor _23247_ (_01377_, _06882_, _06897_);
  nand _23248_ (_01378_, _01377_, _11223_);
  nand _23249_ (_01379_, _01378_, _11203_);
  and _23250_ (_01380_, _01379_, _01376_);
  or _23251_ (_01381_, _01380_, _11193_);
  and _23252_ (_01382_, _11193_, _06897_);
  nor _23253_ (_01383_, _01382_, _11234_);
  and _23254_ (_01384_, _01383_, _01381_);
  and _23255_ (_01385_, _11234_, _06799_);
  or _23256_ (_01386_, _01385_, _11239_);
  or _23257_ (_01387_, _01386_, _01384_);
  nand _23258_ (_01388_, _11239_, _06885_);
  and _23259_ (_01389_, _01388_, _05110_);
  and _23260_ (_01752_, _01389_, _01387_);
  or _23261_ (_01390_, _06137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23262_ (_01391_, _01390_, _05110_);
  or _23263_ (_01392_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _05850_);
  and _23264_ (_01393_, _01392_, _06103_);
  or _23265_ (_01394_, _01393_, _06105_);
  and _23266_ (_01395_, _05980_, _05859_);
  or _23267_ (_01396_, _01219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nand _23268_ (_01397_, _01396_, _01222_);
  nand _23269_ (_01398_, _01397_, _06104_);
  or _23270_ (_01399_, _01398_, _01395_);
  and _23271_ (_01400_, _01399_, _01394_);
  and _23272_ (_01401_, _05976_, _05859_);
  or _23273_ (_01402_, _01401_, _01400_);
  and _23274_ (_01403_, _01402_, _06099_);
  and _23275_ (_01404_, _05971_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23276_ (_01405_, _01152_, _05859_);
  or _23277_ (_01406_, _01239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _23278_ (_01407_, _01242_, _05967_);
  and _23279_ (_01408_, _01407_, _01406_);
  not _23280_ (_01409_, _05967_);
  and _23281_ (_01410_, _01392_, _01409_);
  or _23282_ (_01411_, _01410_, _01408_);
  and _23283_ (_01412_, _01411_, _05960_);
  or _23284_ (_01413_, _01412_, _01405_);
  and _23285_ (_01414_, _01413_, _01139_);
  nor _23286_ (_01415_, _01414_, _01404_);
  nor _23287_ (_01416_, _01415_, _06099_);
  or _23288_ (_01417_, _01416_, _01403_);
  or _23289_ (_01418_, _01417_, _05986_);
  and _23290_ (_01756_, _01418_, _01391_);
  and _23291_ (_01419_, _01216_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _23292_ (_01420_, _01128_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _23293_ (_01421_, _01420_, _01131_);
  or _23294_ (_01422_, _06114_, _05851_);
  and _23295_ (_01423_, _01422_, _01421_);
  or _23296_ (_01424_, _01423_, _05979_);
  or _23297_ (_01425_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _23298_ (_01426_, _01425_, _01228_);
  and _23299_ (_01427_, _01426_, _01227_);
  and _23300_ (_01428_, _01427_, _01424_);
  and _23301_ (_01429_, _05977_, _05851_);
  or _23302_ (_01430_, _01429_, _05976_);
  or _23303_ (_01431_, _01430_, _01428_);
  or _23304_ (_01432_, _01425_, _06103_);
  and _23305_ (_01433_, _01432_, _06099_);
  and _23306_ (_01434_, _01433_, _01431_);
  not _23307_ (_01435_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _23308_ (_01436_, _01145_, _01435_);
  nand _23309_ (_01437_, _01436_, _01144_);
  or _23310_ (_01438_, _05956_, _05851_);
  and _23311_ (_01439_, _01438_, _01437_);
  or _23312_ (_01440_, _01439_, _05966_);
  or _23313_ (_01441_, _01425_, _01248_);
  and _23314_ (_01442_, _01441_, _01247_);
  and _23315_ (_01443_, _01442_, _01440_);
  and _23316_ (_01444_, _05963_, _05851_);
  or _23317_ (_01445_, _01444_, _05959_);
  or _23318_ (_01446_, _01445_, _01443_);
  and _23319_ (_01448_, _01425_, _06100_);
  or _23320_ (_01449_, _01448_, _01255_);
  and _23321_ (_01450_, _01449_, _01446_);
  or _23322_ (_01451_, _01450_, _01434_);
  and _23323_ (_01452_, _01451_, _06137_);
  or _23324_ (_01454_, _01452_, _01419_);
  and _23325_ (_01759_, _01454_, _05110_);
  nand _23326_ (_01455_, _06100_, _06092_);
  and _23327_ (_01456_, _06092_, _06099_);
  or _23328_ (_01457_, _01456_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and _23329_ (_01458_, _01457_, _05110_);
  and _23330_ (_01763_, _01458_, _01455_);
  nor _23331_ (_01461_, _05986_, _05850_);
  and _23332_ (_01462_, _01461_, _06099_);
  or _23333_ (_01464_, _01462_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  nand _23334_ (_01466_, _01461_, _06100_);
  and _23335_ (_01467_, _01466_, _05110_);
  and _23336_ (_01767_, _01467_, _01464_);
  and _23337_ (_01469_, _06123_, _05805_);
  or _23338_ (_01470_, _01469_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _23339_ (_01472_, _01470_, _06130_);
  nand _23340_ (_01473_, _01469_, _05872_);
  and _23341_ (_01474_, _01473_, _01472_);
  and _23342_ (_01476_, _06799_, _06129_);
  or _23343_ (_01477_, _01476_, _01474_);
  and _23344_ (_01795_, _01477_, _05110_);
  and _23345_ (_01480_, _06632_, _06123_);
  nand _23346_ (_01481_, _06123_, _05401_);
  or _23347_ (_01482_, _01481_, _11548_);
  and _23348_ (_01483_, _01482_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _23349_ (_01484_, _01483_, _06129_);
  or _23350_ (_01485_, _01484_, _01480_);
  nand _23351_ (_01486_, _06129_, _06088_);
  and _23352_ (_01487_, _01486_, _05110_);
  and _23353_ (_01799_, _01487_, _01485_);
  and _23354_ (_01489_, _06173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _23355_ (_01490_, _01489_, _08245_);
  and _23356_ (_01491_, _01490_, _06123_);
  nand _23357_ (_01492_, _06123_, _11559_);
  and _23358_ (_01493_, _01492_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _23359_ (_01495_, _01493_, _06129_);
  or _23360_ (_01496_, _01495_, _01491_);
  nand _23361_ (_01497_, _06229_, _06129_);
  and _23362_ (_01499_, _01497_, _05110_);
  and _23363_ (_01801_, _01499_, _01496_);
  and _23364_ (_01501_, _06123_, _05488_);
  nand _23365_ (_01502_, _01501_, _05872_);
  or _23366_ (_01503_, _01501_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _23367_ (_01504_, _01503_, _06130_);
  and _23368_ (_01505_, _01504_, _01502_);
  nor _23369_ (_01506_, _06130_, _05841_);
  or _23370_ (_01507_, _01506_, _01505_);
  and _23371_ (_01804_, _01507_, _05110_);
  and _23372_ (_01508_, _06153_, _05805_);
  or _23373_ (_01509_, _01508_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _23374_ (_01510_, _01509_, _06149_);
  nand _23375_ (_01511_, _01508_, _05872_);
  and _23376_ (_01512_, _01511_, _01510_);
  and _23377_ (_01514_, _06799_, _06148_);
  or _23378_ (_01515_, _01514_, _01512_);
  and _23379_ (_01812_, _01515_, _05110_);
  and _23380_ (_01517_, _06632_, _01079_);
  nand _23381_ (_01518_, _01079_, _05401_);
  or _23382_ (_01519_, _01518_, _11548_);
  and _23383_ (_01521_, _01519_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _23384_ (_01523_, _01521_, _06148_);
  or _23385_ (_01524_, _01523_, _01517_);
  nand _23386_ (_01525_, _06148_, _06088_);
  and _23387_ (_01526_, _01525_, _05110_);
  and _23388_ (_01822_, _01526_, _01524_);
  or _23389_ (_01528_, _01518_, _05866_);
  and _23390_ (_01529_, _01528_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _23391_ (_01530_, _01529_, _06148_);
  and _23392_ (_01532_, _06173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _23393_ (_01533_, _01532_, _08245_);
  and _23394_ (_01534_, _01533_, _06153_);
  or _23395_ (_01535_, _01534_, _01530_);
  nand _23396_ (_01536_, _06229_, _06148_);
  and _23397_ (_01537_, _01536_, _05110_);
  and _23398_ (_01826_, _01537_, _01535_);
  and _23399_ (_01538_, _06153_, _05488_);
  or _23400_ (_01539_, _01538_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _23401_ (_01541_, _01539_, _06149_);
  nand _23402_ (_01542_, _01538_, _05872_);
  and _23403_ (_01543_, _01542_, _01541_);
  nor _23404_ (_01544_, _06149_, _05841_);
  or _23405_ (_01545_, _01544_, _01543_);
  and _23406_ (_01845_, _01545_, _05110_);
  or _23407_ (_01546_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _23408_ (_01547_, _01546_, _11326_);
  and _23409_ (_01548_, _05867_, _05782_);
  nand _23410_ (_01549_, _12083_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _23411_ (_01550_, _01549_, _11326_);
  or _23412_ (_01551_, _01550_, _01548_);
  and _23413_ (_01552_, _01551_, _01547_);
  or _23414_ (_01553_, _01552_, _11329_);
  nand _23415_ (_01554_, _11329_, _05901_);
  and _23416_ (_01555_, _01554_, _05110_);
  and _23417_ (_01851_, _01555_, _01553_);
  nand _23418_ (_01556_, _06890_, _05901_);
  and _23419_ (_01557_, _08872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _23420_ (_01558_, _06883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _23421_ (_01559_, _01558_, _01557_);
  or _23422_ (_01560_, _01559_, _06890_);
  and _23423_ (_01562_, _01560_, _08871_);
  and _23424_ (_01563_, _01562_, _01556_);
  and _23425_ (_01564_, _06895_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _23426_ (_01566_, _01564_, _01563_);
  and _23427_ (_01860_, _01566_, _05110_);
  and _23428_ (_01568_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _23429_ (_01569_, pc_log_change, _05478_);
  or _23430_ (_01570_, _01569_, _01568_);
  and _23431_ (_01869_, _01570_, _05110_);
  nor _23432_ (_01572_, _05841_, _06010_);
  and _23433_ (_01573_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _23434_ (_01575_, _01573_, _05995_);
  or _23435_ (_01576_, _01575_, _01572_);
  or _23436_ (_01578_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _23437_ (_01579_, _01578_, _05110_);
  and _23438_ (_01905_, _01579_, _01576_);
  nor _23439_ (_01580_, _11584_, _11515_);
  and _23440_ (_01582_, _11192_, _06881_);
  and _23441_ (_01583_, _01582_, _11202_);
  and _23442_ (_01584_, _01583_, _11223_);
  and _23443_ (_01585_, _01584_, _11584_);
  or _23444_ (_01586_, _01585_, _01580_);
  and _23445_ (_01908_, _01586_, _05110_);
  nand _23446_ (_01587_, _11239_, _05901_);
  or _23447_ (_01588_, _12560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _23448_ (_01589_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _23449_ (_01591_, _01589_, _11202_);
  nand _23450_ (_01592_, _01591_, _11223_);
  and _23451_ (_01594_, _01592_, _01588_);
  or _23452_ (_01595_, _01594_, _11193_);
  nor _23453_ (_01596_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor _23454_ (_01597_, _01596_, _11234_);
  and _23455_ (_01598_, _01597_, _01595_);
  and _23456_ (_01599_, _11234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _23457_ (_01601_, _01599_, _11239_);
  or _23458_ (_01602_, _01601_, _01598_);
  and _23459_ (_01603_, _01602_, _05110_);
  and _23460_ (_01911_, _01603_, _01587_);
  nor _23461_ (_01605_, _12612_, _05901_);
  and _23462_ (_01606_, _11601_, _11215_);
  and _23463_ (_01607_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _23464_ (_01608_, _01607_, _11223_);
  or _23465_ (_01609_, _01608_, _01606_);
  and _23466_ (_01610_, _01609_, _11202_);
  and _23467_ (_01611_, _11601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _23468_ (_01612_, _01611_, _11193_);
  or _23469_ (_01613_, _01612_, _01610_);
  nor _23470_ (_01614_, _11194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor _23471_ (_01616_, _01614_, _11234_);
  and _23472_ (_01617_, _01616_, _01613_);
  or _23473_ (_01618_, _01617_, _11239_);
  or _23474_ (_01620_, _01618_, _01605_);
  or _23475_ (_01621_, _11240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _23476_ (_01622_, _01621_, _05110_);
  and _23477_ (_01914_, _01622_, _01620_);
  and _23478_ (_01623_, _11202_, _11190_);
  and _23479_ (_01624_, _01623_, _11584_);
  or _23480_ (_01625_, _01624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _23481_ (_01626_, _11223_);
  nand _23482_ (_01627_, _01624_, _01626_);
  and _23483_ (_01628_, _01627_, _05110_);
  and _23484_ (_01917_, _01628_, _01625_);
  nand _23485_ (_01629_, _08870_, _05901_);
  and _23486_ (_01630_, _08886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _23487_ (_01631_, _08884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _23488_ (_01632_, _01631_, _01630_);
  or _23489_ (_01633_, _01632_, _08870_);
  and _23490_ (_01634_, _01633_, _05110_);
  and _23491_ (_01920_, _01634_, _01629_);
  and _23492_ (_01931_, t2ex_i, _05110_);
  nor _23493_ (_01635_, t2ex_i, rst);
  and _23494_ (_01934_, _01635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  nor _23495_ (_01637_, t2_i, rst);
  and _23496_ (_01937_, _01637_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  and _23497_ (_01940_, t2_i, _05110_);
  or _23498_ (_01638_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not _23499_ (_01639_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _23500_ (_01640_, pc_log_change, _01639_);
  and _23501_ (_01641_, _01640_, _05110_);
  and _23502_ (_02010_, _01641_, _01638_);
  or _23503_ (_01642_, _06860_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _23504_ (_01643_, _06861_, _05110_);
  and _23505_ (_01644_, _01643_, _01642_);
  and _23506_ (_01645_, _06811_, _06434_);
  or _23507_ (_01647_, _01645_, _06947_);
  or _23508_ (_01648_, _01647_, _06816_);
  and _23509_ (_01649_, _07079_, _07040_);
  or _23510_ (_01650_, _01649_, _07046_);
  or _23511_ (_01651_, _07081_, _06453_);
  or _23512_ (_01652_, _01651_, _07089_);
  or _23513_ (_01653_, _01652_, _01650_);
  or _23514_ (_01654_, _01653_, _01648_);
  or _23515_ (_01655_, _07093_, _07052_);
  or _23516_ (_01656_, _01655_, _07074_);
  and _23517_ (_01657_, _06457_, _07067_);
  and _23518_ (_01658_, _06852_, _06455_);
  or _23519_ (_01659_, _01658_, _01657_);
  or _23520_ (_01660_, _01659_, _07078_);
  or _23521_ (_01661_, _01660_, _06449_);
  or _23522_ (_01662_, _07048_, _07041_);
  or _23523_ (_01663_, _01662_, _01661_);
  and _23524_ (_01664_, _13086_, _06434_);
  and _23525_ (_01665_, _07138_, _06464_);
  or _23526_ (_01666_, _01665_, _01664_);
  and _23527_ (_01667_, _07079_, _06830_);
  or _23528_ (_01668_, _01667_, _07039_);
  and _23529_ (_01670_, _07087_, _06434_);
  or _23530_ (_01671_, _01670_, _01668_);
  or _23531_ (_01672_, _01671_, _01666_);
  or _23532_ (_01673_, _13078_, _11749_);
  not _23533_ (_01674_, _07095_);
  nand _23534_ (_01675_, _11300_, _01674_);
  or _23535_ (_01676_, _01675_, _01673_);
  or _23536_ (_01677_, _01676_, _01672_);
  or _23537_ (_01678_, _01677_, _01663_);
  or _23538_ (_01679_, _01678_, _01656_);
  or _23539_ (_01680_, _01679_, _01654_);
  and _23540_ (_01681_, _01680_, _06842_);
  or _23541_ (_02048_, _01681_, _01644_);
  nand _23542_ (_01682_, _06294_, _05473_);
  or _23543_ (_01683_, _05473_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _23544_ (_01684_, _01683_, _05110_);
  and _23545_ (_02086_, _01684_, _01682_);
  and _23546_ (_01685_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _23547_ (_01686_, _05938_, _06010_);
  or _23548_ (_01687_, _01686_, _01685_);
  or _23549_ (_01688_, _01687_, _05995_);
  or _23550_ (_01689_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _23551_ (_01690_, _01689_, _05110_);
  and _23552_ (_02207_, _01690_, _01688_);
  nand _23553_ (_01691_, _06673_, _05938_);
  or _23554_ (_01692_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _23555_ (_01693_, _01692_, _05110_);
  and _23556_ (_02218_, _01693_, _01691_);
  nor _23557_ (_01694_, _06088_, _06010_);
  and _23558_ (_01695_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _23559_ (_01696_, _01695_, _05995_);
  or _23560_ (_01697_, _01696_, _01694_);
  or _23561_ (_01698_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _23562_ (_01699_, _01698_, _05110_);
  and _23563_ (_02222_, _01699_, _01697_);
  or _23564_ (_01700_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand _23565_ (_01701_, _06205_, _12450_);
  and _23566_ (_01702_, _01701_, _05110_);
  and _23567_ (_02255_, _01702_, _01700_);
  and _23568_ (_01703_, _06807_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _23569_ (_01704_, _07075_, _13076_);
  or _23570_ (_01705_, _01704_, _01652_);
  or _23571_ (_01706_, _11760_, _07096_);
  and _23572_ (_01707_, _12149_, _06864_);
  and _23573_ (_01708_, _01665_, _11802_);
  or _23574_ (_01709_, _01708_, _01707_);
  or _23575_ (_01710_, _01709_, _01706_);
  or _23576_ (_01711_, _06838_, _06828_);
  and _23577_ (_01712_, _07069_, _06434_);
  and _23578_ (_01713_, _07038_, _06434_);
  or _23579_ (_01714_, _01713_, _13078_);
  or _23580_ (_01715_, _01714_, _01712_);
  or _23581_ (_01716_, _01715_, _01711_);
  or _23582_ (_01717_, _01716_, _01710_);
  or _23583_ (_01718_, _01717_, _01705_);
  and _23584_ (_01719_, _01718_, _06842_);
  or _23585_ (_02391_, _01719_, _01703_);
  not _23586_ (_01720_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _23587_ (_01721_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and _23588_ (_01722_, _01721_, _01720_);
  and _23589_ (_01723_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _05110_);
  and _23590_ (_02407_, _01723_, _01722_);
  and _23591_ (_01724_, _12330_, _12228_);
  nand _23592_ (_01725_, _12018_, _11977_);
  and _23593_ (_01726_, _12073_, _01725_);
  and _23594_ (_01727_, _01726_, _11918_);
  and _23595_ (_01728_, _01727_, _11960_);
  and _23596_ (_01729_, _12268_, _11871_);
  and _23597_ (_01730_, _01729_, _01728_);
  and _23598_ (_01731_, _01730_, _01724_);
  and _23599_ (_01732_, _01731_, _06471_);
  and _23600_ (_01733_, _12071_, _01725_);
  and _23601_ (_01734_, _01733_, _11918_);
  and _23602_ (_01735_, _01734_, _11960_);
  and _23603_ (_01736_, _12268_, _11873_);
  and _23604_ (_01737_, _12330_, _12225_);
  and _23605_ (_01738_, _01737_, _01736_);
  and _23606_ (_01739_, _01738_, _01735_);
  and _23607_ (_01740_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _23608_ (_01742_, _12270_, _11873_);
  and _23609_ (_01743_, _01737_, _01742_);
  and _23610_ (_01744_, _01743_, _01735_);
  and _23611_ (_01745_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _23612_ (_01747_, _01745_, _01740_);
  and _23613_ (_01748_, _12328_, _12225_);
  and _23614_ (_01749_, _01748_, _01742_);
  and _23615_ (_01750_, _01749_, _01735_);
  and _23616_ (_01751_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _23617_ (_01753_, _01724_, _01736_);
  and _23618_ (_01754_, _01753_, _01735_);
  and _23619_ (_01755_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _23620_ (_01757_, _01755_, _01751_);
  or _23621_ (_01758_, _01757_, _01747_);
  and _23622_ (_01760_, _01738_, _01728_);
  and _23623_ (_01761_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _23624_ (_01762_, _12328_, _12228_);
  and _23625_ (_01764_, _01762_, _01736_);
  and _23626_ (_01765_, _01764_, _01735_);
  and _23627_ (_01766_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or _23628_ (_01768_, _01766_, _01761_);
  and _23629_ (_01769_, _01726_, _11920_);
  and _23630_ (_01770_, _01769_, _11958_);
  or _23631_ (_01771_, _12330_, _12225_);
  or _23632_ (_01772_, _01771_, _12268_);
  nor _23633_ (_01773_, _01772_, _11873_);
  and _23634_ (_01774_, _01773_, _01770_);
  and _23635_ (_01775_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _23636_ (_01776_, _01769_, _11960_);
  and _23637_ (_01777_, _01776_, _01738_);
  and _23638_ (_01778_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _23639_ (_01779_, _01778_, _01775_);
  or _23640_ (_01780_, _01779_, _01768_);
  or _23641_ (_01781_, _01780_, _01758_);
  and _23642_ (_01782_, _01736_, _01748_);
  and _23643_ (_01783_, _01728_, _01782_);
  and _23644_ (_01784_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _23645_ (_01785_, _01764_, _01728_);
  and _23646_ (_01786_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or _23647_ (_01787_, _01786_, _01784_);
  and _23648_ (_01788_, _01753_, _01728_);
  and _23649_ (_01789_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _23650_ (_01790_, _01728_, _01749_);
  and _23651_ (_01791_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _23652_ (_01792_, _01791_, _01789_);
  or _23653_ (_01793_, _01792_, _01787_);
  and _23654_ (_01794_, _01727_, _11958_);
  and _23655_ (_01796_, _01794_, _01782_);
  and _23656_ (_01797_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _23657_ (_01798_, _01738_, _01794_);
  and _23658_ (_01800_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _23659_ (_01802_, _01800_, _01797_);
  and _23660_ (_01803_, _01743_, _01728_);
  and _23661_ (_01805_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _23662_ (_01806_, _01773_, _01728_);
  and _23663_ (_01807_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _23664_ (_01808_, _01807_, _01805_);
  or _23665_ (_01809_, _01808_, _01802_);
  or _23666_ (_01810_, _01809_, _01793_);
  or _23667_ (_01811_, _01810_, _01781_);
  and _23668_ (_01813_, _01737_, _01729_);
  and _23669_ (_01814_, _01813_, _11958_);
  and _23670_ (_01815_, _01733_, _11920_);
  and _23671_ (_01816_, _01815_, _01814_);
  and _23672_ (_01817_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _23673_ (_01818_, _01729_, _01748_);
  and _23674_ (_01819_, _01818_, _01728_);
  and _23675_ (_01820_, _01819_, _11976_);
  or _23676_ (_01821_, _01820_, _01817_);
  and _23677_ (_01823_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _23678_ (_01824_, _01762_, _01729_);
  and _23679_ (_01825_, _01824_, _01728_);
  and _23680_ (_01827_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _23681_ (_01828_, _01827_, _01823_);
  or _23682_ (_01829_, _01828_, _01821_);
  and _23683_ (_01830_, _01770_, _01813_);
  and _23684_ (_01831_, _07079_, _06431_);
  nor _23685_ (_01832_, _01831_, _06817_);
  and _23686_ (_01833_, _01832_, _06834_);
  nor _23687_ (_01834_, _01649_, _07074_);
  and _23688_ (_01835_, _01834_, _01833_);
  nor _23689_ (_01836_, _01665_, _11755_);
  nor _23690_ (_01837_, _06938_, _06823_);
  and _23691_ (_01838_, _07069_, _06810_);
  nor _23692_ (_01839_, _01838_, _07095_);
  and _23693_ (_01840_, _01839_, _01837_);
  and _23694_ (_01841_, _01840_, _11747_);
  and _23695_ (_01842_, _01841_, _01836_);
  and _23696_ (_01843_, _01842_, _01835_);
  and _23697_ (_01844_, _01843_, _11746_);
  nor _23698_ (_01846_, _01844_, _12089_);
  or _23699_ (_01847_, _01846_, p3_in[7]);
  not _23700_ (_01848_, _01846_);
  or _23701_ (_01849_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _23702_ (_01850_, _01849_, _01847_);
  and _23703_ (_01852_, _01850_, _01830_);
  and _23704_ (_01853_, _01776_, _01813_);
  or _23705_ (_01854_, _01846_, p2_in[7]);
  or _23706_ (_01855_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _23707_ (_01856_, _01855_, _01854_);
  and _23708_ (_01857_, _01856_, _01853_);
  or _23709_ (_01858_, _01857_, _01852_);
  and _23710_ (_01859_, _01813_, _01728_);
  or _23711_ (_01861_, _01846_, p0_in[7]);
  or _23712_ (_01862_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _23713_ (_01863_, _01862_, _01861_);
  and _23714_ (_01864_, _01863_, _01859_);
  and _23715_ (_01865_, _01813_, _01794_);
  or _23716_ (_01866_, _01846_, p1_in[7]);
  or _23717_ (_01867_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _23718_ (_01868_, _01867_, _01866_);
  and _23719_ (_01870_, _01868_, _01865_);
  or _23720_ (_01871_, _01870_, _01864_);
  or _23721_ (_01872_, _01871_, _01858_);
  or _23722_ (_01873_, _01872_, _01829_);
  and _23723_ (_01874_, _01814_, _01734_);
  and _23724_ (_01875_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _23725_ (_01876_, _01813_, _11960_);
  and _23726_ (_01877_, _01815_, _01876_);
  and _23727_ (_01878_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _23728_ (_01879_, _01878_, _01875_);
  or _23729_ (_01880_, _01879_, _01873_);
  or _23730_ (_01881_, _01880_, _01811_);
  nand _23731_ (_01882_, _01874_, _12172_);
  nand _23732_ (_01883_, _01877_, _06613_);
  and _23733_ (_01884_, _01883_, _01882_);
  nand _23734_ (_01885_, _01825_, _06471_);
  nand _23735_ (_01886_, _01885_, _01884_);
  nand _23736_ (_01887_, _01886_, _05151_);
  nand _23737_ (_01888_, _01877_, _06617_);
  and _23738_ (_01889_, _01772_, _06150_);
  nand _23739_ (_01890_, _01889_, _12082_);
  and _23740_ (_01891_, _01890_, _01888_);
  and _23741_ (_01892_, _01891_, _12340_);
  and _23742_ (_01893_, _01892_, _01887_);
  and _23743_ (_01894_, _01893_, _01881_);
  nor _23744_ (_01895_, _01877_, _01874_);
  nand _23745_ (_01896_, _01813_, _01726_);
  nor _23746_ (_01897_, _01825_, _01731_);
  nor _23747_ (_01898_, _01819_, _01816_);
  and _23748_ (_01899_, _01898_, _01897_);
  and _23749_ (_01900_, _01899_, _01896_);
  and _23750_ (_01901_, _01900_, _01895_);
  nor _23751_ (_01902_, _01744_, _01739_);
  nand _23752_ (_01903_, _01733_, _11918_);
  or _23753_ (_01904_, _01903_, _11958_);
  not _23754_ (_01906_, _01742_);
  or _23755_ (_01907_, _12330_, _12228_);
  or _23756_ (_01909_, _01907_, _01906_);
  or _23757_ (_01910_, _01909_, _01904_);
  nand _23758_ (_01912_, _01724_, _01736_);
  or _23759_ (_01913_, _01912_, _01904_);
  and _23760_ (_01915_, _01913_, _01910_);
  and _23761_ (_01916_, _01915_, _01902_);
  or _23762_ (_01918_, _12071_, _12020_);
  or _23763_ (_01919_, _01918_, _11920_);
  or _23764_ (_01921_, _01919_, _11958_);
  not _23765_ (_01922_, _01736_);
  or _23766_ (_01923_, _12328_, _12228_);
  or _23767_ (_01924_, _01923_, _01922_);
  or _23768_ (_01925_, _01924_, _01921_);
  or _23769_ (_01926_, _01771_, _01922_);
  or _23770_ (_01927_, _01926_, _01904_);
  and _23771_ (_01928_, _01927_, _01925_);
  nor _23772_ (_01929_, _01777_, _01774_);
  and _23773_ (_01930_, _01929_, _01928_);
  and _23774_ (_01932_, _01930_, _01916_);
  or _23775_ (_01933_, _01922_, _01907_);
  or _23776_ (_01935_, _01921_, _01933_);
  or _23777_ (_01936_, _01926_, _01921_);
  and _23778_ (_01938_, _01936_, _01935_);
  nor _23779_ (_01939_, _01790_, _01788_);
  and _23780_ (_01941_, _01939_, _01938_);
  nor _23781_ (_01942_, _01806_, _01803_);
  nor _23782_ (_01943_, _01798_, _01796_);
  and _23783_ (_01944_, _01943_, _01942_);
  and _23784_ (_01945_, _01944_, _01941_);
  and _23785_ (_01946_, _01945_, _01932_);
  nand _23786_ (_01947_, _01946_, _01901_);
  nand _23787_ (_01948_, _01947_, _01893_);
  and _23788_ (_01949_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or _23789_ (_01950_, _01949_, _01894_);
  or _23790_ (_01951_, _01950_, _01732_);
  nand _23791_ (_01952_, _01732_, _07028_);
  and _23792_ (_01953_, _01952_, _05110_);
  and _23793_ (_02423_, _01953_, _01951_);
  and _23794_ (_01954_, _00523_, _10209_);
  nand _23795_ (_01955_, _00523_, _10208_);
  and _23796_ (_01956_, _01955_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _23797_ (_01957_, _01956_, _01954_);
  and _23798_ (_01958_, _01957_, _05794_);
  and _23799_ (_01959_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _23800_ (_01960_, _00531_, _07235_);
  or _23801_ (_01961_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _23802_ (_01962_, _01961_, _05806_);
  and _23803_ (_01963_, _01962_, _01960_);
  or _23804_ (_01964_, _01963_, _01959_);
  or _23805_ (_01965_, _01964_, _01958_);
  and _23806_ (_02463_, _01965_, _05110_);
  and _23807_ (_01966_, _00523_, _08272_);
  nand _23808_ (_01967_, _01966_, _05872_);
  or _23809_ (_01968_, _01966_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _23810_ (_01969_, _01968_, _05794_);
  and _23811_ (_01970_, _01969_, _01967_);
  and _23812_ (_01971_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _23813_ (_01972_, _00550_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor _23814_ (_01973_, _00550_, _06512_);
  or _23815_ (_01974_, _01973_, _01972_);
  and _23816_ (_01975_, _01974_, _05806_);
  or _23817_ (_01976_, _01975_, _01971_);
  or _23818_ (_01977_, _01976_, _01970_);
  and _23819_ (_02466_, _01977_, _05110_);
  and _23820_ (_02472_, _11976_, _05110_);
  or _23821_ (_01978_, _01732_, rst);
  nor _23822_ (_02476_, _01978_, _01893_);
  and _23823_ (_01979_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _23824_ (_01980_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _23825_ (_02503_, _01980_, _01979_);
  and _23826_ (_01981_, _06625_, _06122_);
  and _23827_ (_01982_, _01981_, _08133_);
  nand _23828_ (_01983_, _01982_, _05872_);
  or _23829_ (_01984_, _01982_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _23830_ (_01985_, _01984_, _05794_);
  and _23831_ (_01986_, _01985_, _01983_);
  and _23832_ (_01987_, _06128_, _05992_);
  not _23833_ (_01988_, _01987_);
  nor _23834_ (_01989_, _01988_, _06054_);
  and _23835_ (_01990_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _23836_ (_01991_, _01990_, _01989_);
  and _23837_ (_01992_, _01991_, _05806_);
  and _23838_ (_01993_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _23839_ (_01994_, _01993_, rst);
  or _23840_ (_01995_, _01994_, _01992_);
  or _23841_ (_02518_, _01995_, _01986_);
  and _23842_ (_01996_, _10154_, _05789_);
  and _23843_ (_01997_, _01996_, _05488_);
  nand _23844_ (_01998_, _01997_, _05872_);
  or _23845_ (_01999_, _01997_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _23846_ (_02000_, _01999_, _05794_);
  and _23847_ (_02001_, _02000_, _01998_);
  and _23848_ (_02002_, _08252_, _05992_);
  nand _23849_ (_02003_, _02002_, _05841_);
  or _23850_ (_02004_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _23851_ (_02005_, _02004_, _05806_);
  and _23852_ (_02006_, _02005_, _02003_);
  and _23853_ (_02007_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _23854_ (_02008_, _02007_, rst);
  or _23855_ (_02009_, _02008_, _02006_);
  or _23856_ (_02520_, _02009_, _02001_);
  and _23857_ (_02011_, _01996_, _08272_);
  nand _23858_ (_02012_, _02011_, _05872_);
  or _23859_ (_02013_, _02011_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _23860_ (_02014_, _02013_, _05794_);
  and _23861_ (_02015_, _02014_, _02012_);
  nand _23862_ (_02016_, _02002_, _05938_);
  or _23863_ (_02017_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _23864_ (_02018_, _02017_, _05806_);
  and _23865_ (_02019_, _02018_, _02016_);
  and _23866_ (_02020_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _23867_ (_02021_, _02020_, rst);
  or _23868_ (_02022_, _02021_, _02019_);
  or _23869_ (_02522_, _02022_, _02015_);
  nand _23870_ (_02023_, _01174_, _11559_);
  and _23871_ (_02024_, _02023_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _23872_ (_02025_, _06173_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _23873_ (_02026_, _02025_, _08245_);
  and _23874_ (_02027_, _02026_, _01174_);
  or _23875_ (_02028_, _02027_, _02024_);
  and _23876_ (_02029_, _02028_, _05794_);
  nand _23877_ (_02030_, _01180_, _06229_);
  or _23878_ (_02031_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _23879_ (_02032_, _02031_, _05806_);
  and _23880_ (_02033_, _02032_, _02030_);
  and _23881_ (_02034_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _23882_ (_02035_, _02034_, rst);
  or _23883_ (_02036_, _02035_, _02033_);
  or _23884_ (_02525_, _02036_, _02029_);
  nor _23885_ (_02037_, _08056_, _06054_);
  and _23886_ (_02038_, _08117_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or _23887_ (_02039_, _02038_, _02037_);
  and _23888_ (_02543_, _02039_, _05110_);
  and _23889_ (_02040_, _10154_, _06122_);
  and _23890_ (_02041_, _02040_, _10208_);
  nand _23891_ (_02042_, _02041_, _05872_);
  or _23892_ (_02043_, _02041_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _23893_ (_02044_, _02043_, _05794_);
  and _23894_ (_02045_, _02044_, _02042_);
  and _23895_ (_02046_, _06145_, _05992_);
  not _23896_ (_02047_, _02046_);
  nor _23897_ (_02049_, _02047_, _05334_);
  and _23898_ (_02050_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _23899_ (_02051_, _02050_, _02049_);
  and _23900_ (_02052_, _02051_, _05806_);
  and _23901_ (_02053_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _23902_ (_02054_, _02053_, rst);
  or _23903_ (_02055_, _02054_, _02052_);
  or _23904_ (_02547_, _02055_, _02045_);
  and _23905_ (_02056_, _01981_, _10208_);
  nand _23906_ (_02057_, _02056_, _05872_);
  or _23907_ (_02058_, _02056_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _23908_ (_02059_, _02058_, _05794_);
  and _23909_ (_02060_, _02059_, _02057_);
  nor _23910_ (_02061_, _01988_, _05334_);
  and _23911_ (_02062_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _23912_ (_02063_, _02062_, _02061_);
  and _23913_ (_02064_, _02063_, _05806_);
  and _23914_ (_02065_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _23915_ (_02066_, _02065_, rst);
  or _23916_ (_02067_, _02066_, _02064_);
  or _23917_ (_02549_, _02067_, _02060_);
  and _23918_ (_02068_, _01996_, _08133_);
  nand _23919_ (_02069_, _02068_, _05872_);
  or _23920_ (_02070_, _02068_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _23921_ (_02071_, _02070_, _05794_);
  and _23922_ (_02072_, _02071_, _02069_);
  nand _23923_ (_02073_, _02002_, _06054_);
  or _23924_ (_02074_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _23925_ (_02075_, _02074_, _05806_);
  and _23926_ (_02076_, _02075_, _02073_);
  and _23927_ (_02077_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _23928_ (_02078_, _02077_, rst);
  or _23929_ (_02079_, _02078_, _02076_);
  or _23930_ (_02553_, _02079_, _02072_);
  not _23931_ (_02080_, _02002_);
  or _23932_ (_02081_, _02080_, _05782_);
  or _23933_ (_02082_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _23934_ (_02083_, _02082_, _05794_);
  and _23935_ (_02084_, _02083_, _02081_);
  nand _23936_ (_02085_, _02002_, _06798_);
  and _23937_ (_02087_, _02082_, _05806_);
  and _23938_ (_02088_, _02087_, _02085_);
  not _23939_ (_02089_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor _23940_ (_02090_, _05793_, _02089_);
  or _23941_ (_02091_, _02090_, rst);
  or _23942_ (_02092_, _02091_, _02088_);
  or _23943_ (_02555_, _02092_, _02084_);
  and _23944_ (_02093_, _01996_, _06631_);
  nand _23945_ (_02094_, _02093_, _05872_);
  or _23946_ (_02095_, _02093_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _23947_ (_02096_, _02095_, _05794_);
  and _23948_ (_02097_, _02096_, _02094_);
  nand _23949_ (_02098_, _02002_, _06088_);
  or _23950_ (_02099_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _23951_ (_02100_, _02099_, _05806_);
  and _23952_ (_02101_, _02100_, _02098_);
  and _23953_ (_02102_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _23954_ (_02103_, _02102_, rst);
  or _23955_ (_02104_, _02103_, _02101_);
  or _23956_ (_02557_, _02104_, _02097_);
  and _23957_ (_02105_, _01174_, _05488_);
  nand _23958_ (_02106_, _02105_, _05872_);
  or _23959_ (_02107_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _23960_ (_02108_, _02107_, _05794_);
  and _23961_ (_02109_, _02108_, _02106_);
  nand _23962_ (_02110_, _01180_, _05841_);
  or _23963_ (_02111_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _23964_ (_02112_, _02111_, _05806_);
  and _23965_ (_02113_, _02112_, _02110_);
  and _23966_ (_02114_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _23967_ (_02115_, _02114_, rst);
  or _23968_ (_02116_, _02115_, _02113_);
  or _23969_ (_02559_, _02116_, _02109_);
  and _23970_ (_02117_, _05804_, _05996_);
  nand _23971_ (_02118_, _02117_, _05872_);
  or _23972_ (_02119_, _02117_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _23973_ (_02120_, _02119_, _05794_);
  and _23974_ (_02121_, _02120_, _02118_);
  nand _23975_ (_02122_, _01180_, _05938_);
  or _23976_ (_02123_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _23977_ (_02124_, _02123_, _05806_);
  and _23978_ (_02125_, _02124_, _02122_);
  and _23979_ (_02126_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _23980_ (_02127_, _02126_, rst);
  or _23981_ (_02128_, _02127_, _02125_);
  or _23982_ (_02562_, _02128_, _02121_);
  and _23983_ (_02129_, _01174_, _10208_);
  nand _23984_ (_02130_, _02129_, _05872_);
  or _23985_ (_02131_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _23986_ (_02132_, _02131_, _05794_);
  and _23987_ (_02133_, _02132_, _02130_);
  nand _23988_ (_02134_, _01180_, _05334_);
  or _23989_ (_02135_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _23990_ (_02136_, _02135_, _05806_);
  and _23991_ (_02137_, _02136_, _02134_);
  and _23992_ (_02138_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _23993_ (_02139_, _02138_, rst);
  or _23994_ (_02140_, _02139_, _02137_);
  or _23995_ (_02565_, _02140_, _02133_);
  nand _23996_ (_02141_, _06560_, _06054_);
  or _23997_ (_02142_, _06560_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _23998_ (_02143_, _02142_, _05110_);
  and _23999_ (_02578_, _02143_, _02141_);
  or _24000_ (_02144_, _07141_, _07125_);
  and _24001_ (_02145_, _02144_, _05474_);
  and _24002_ (_02146_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _24003_ (_02147_, _02146_, _07150_);
  or _24004_ (_02148_, _02147_, _02145_);
  and _24005_ (_02587_, _02148_, _05110_);
  and _24006_ (_02602_, _11954_, _05110_);
  and _24007_ (_02149_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _24008_ (_02150_, _02149_, _07149_);
  and _24009_ (_02151_, _02150_, _05110_);
  and _24010_ (_02152_, _07116_, _06277_);
  or _24011_ (_02153_, _06868_, _07065_);
  or _24012_ (_02154_, _02153_, _07134_);
  or _24013_ (_02155_, _02154_, _02152_);
  and _24014_ (_02156_, _02155_, _06842_);
  or _24015_ (_02607_, _02156_, _02151_);
  not _24016_ (_02157_, _08253_);
  and _24017_ (_02158_, _08243_, _05867_);
  or _24018_ (_02159_, _02158_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _24019_ (_02160_, _02159_, _02157_);
  nand _24020_ (_02161_, _02158_, _05872_);
  and _24021_ (_02162_, _02161_, _02160_);
  nor _24022_ (_02163_, _02157_, _05901_);
  or _24023_ (_02164_, _02163_, _02162_);
  and _24024_ (_02626_, _02164_, _05110_);
  and _24025_ (_02165_, _01981_, _06631_);
  nand _24026_ (_02166_, _02165_, _05872_);
  or _24027_ (_02167_, _02165_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _24028_ (_02168_, _02167_, _05794_);
  and _24029_ (_02169_, _02168_, _02166_);
  nor _24030_ (_02170_, _01988_, _06088_);
  and _24031_ (_02171_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _24032_ (_02172_, _02171_, _02170_);
  and _24033_ (_02173_, _02172_, _05806_);
  and _24034_ (_02174_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _24035_ (_02175_, _02174_, rst);
  or _24036_ (_02176_, _02175_, _02173_);
  or _24037_ (_02655_, _02176_, _02169_);
  and _24038_ (_02177_, _01981_, _06472_);
  nand _24039_ (_02178_, _02177_, _05872_);
  or _24040_ (_02179_, _02177_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _24041_ (_02180_, _02179_, _05794_);
  and _24042_ (_02181_, _02180_, _02178_);
  nor _24043_ (_02182_, _01988_, _06229_);
  and _24044_ (_02183_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _24045_ (_02184_, _02183_, _02182_);
  and _24046_ (_02185_, _02184_, _05806_);
  and _24047_ (_02186_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _24048_ (_02187_, _02186_, rst);
  or _24049_ (_02188_, _02187_, _02185_);
  or _24050_ (_02656_, _02188_, _02181_);
  and _24051_ (_02189_, _01981_, _08272_);
  nand _24052_ (_02190_, _02189_, _05872_);
  or _24053_ (_02191_, _02189_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _24054_ (_02192_, _02191_, _05794_);
  and _24055_ (_02193_, _02192_, _02190_);
  nor _24056_ (_02194_, _01988_, _05938_);
  and _24057_ (_02195_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _24058_ (_02196_, _02195_, _02194_);
  and _24059_ (_02197_, _02196_, _05806_);
  and _24060_ (_02198_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _24061_ (_02199_, _02198_, rst);
  or _24062_ (_02200_, _02199_, _02197_);
  or _24063_ (_02666_, _02200_, _02193_);
  and _24064_ (_02201_, _02040_, _06472_);
  nand _24065_ (_02202_, _02201_, _05872_);
  or _24066_ (_02203_, _02201_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _24067_ (_02204_, _02203_, _05794_);
  and _24068_ (_02205_, _02204_, _02202_);
  nor _24069_ (_02206_, _02047_, _06229_);
  and _24070_ (_02208_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _24071_ (_02209_, _02208_, _02206_);
  and _24072_ (_02210_, _02209_, _05806_);
  and _24073_ (_02211_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _24074_ (_02212_, _02211_, rst);
  or _24075_ (_02213_, _02212_, _02210_);
  or _24076_ (_02668_, _02213_, _02205_);
  and _24077_ (_02214_, _02040_, _08272_);
  nand _24078_ (_02215_, _02214_, _05872_);
  or _24079_ (_02216_, _02214_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _24080_ (_02217_, _02216_, _05794_);
  and _24081_ (_02219_, _02217_, _02215_);
  nor _24082_ (_02220_, _02047_, _05938_);
  and _24083_ (_02221_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _24084_ (_02223_, _02221_, _02220_);
  and _24085_ (_02224_, _02223_, _05806_);
  and _24086_ (_02225_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _24087_ (_02226_, _02225_, rst);
  or _24088_ (_02227_, _02226_, _02224_);
  or _24089_ (_02671_, _02227_, _02219_);
  and _24090_ (_02228_, _02040_, _05488_);
  nand _24091_ (_02229_, _02228_, _05872_);
  or _24092_ (_02230_, _02228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _24093_ (_02231_, _02230_, _05794_);
  and _24094_ (_02232_, _02231_, _02229_);
  nor _24095_ (_02233_, _02047_, _05841_);
  and _24096_ (_02234_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _24097_ (_02235_, _02234_, _02233_);
  and _24098_ (_02236_, _02235_, _05806_);
  and _24099_ (_02237_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _24100_ (_02238_, _02237_, rst);
  or _24101_ (_02239_, _02238_, _02236_);
  or _24102_ (_02677_, _02239_, _02232_);
  or _24103_ (_02240_, _08257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _24104_ (_02241_, _02240_, _05110_);
  nand _24105_ (_02242_, _08257_, _05901_);
  and _24106_ (_02688_, _02242_, _02241_);
  nand _24107_ (_02243_, _01174_, _05805_);
  or _24108_ (_02244_, _02243_, _05782_);
  or _24109_ (_02245_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _24110_ (_02246_, _02245_, _05794_);
  and _24111_ (_02247_, _02246_, _02244_);
  nand _24112_ (_02248_, _01180_, _06798_);
  and _24113_ (_02249_, _02245_, _05806_);
  and _24114_ (_02250_, _02249_, _02248_);
  not _24115_ (_02251_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor _24116_ (_02252_, _05793_, _02251_);
  or _24117_ (_02253_, _02252_, rst);
  or _24118_ (_02254_, _02253_, _02250_);
  or _24119_ (_02690_, _02254_, _02247_);
  and _24120_ (_02256_, _01174_, _08133_);
  nand _24121_ (_02257_, _02256_, _05872_);
  or _24122_ (_02258_, _02256_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _24123_ (_02259_, _02258_, _05794_);
  and _24124_ (_02260_, _02259_, _02257_);
  nand _24125_ (_02261_, _01180_, _06054_);
  or _24126_ (_02262_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _24127_ (_02263_, _02262_, _05806_);
  and _24128_ (_02264_, _02263_, _02261_);
  and _24129_ (_02265_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _24130_ (_02266_, _02265_, rst);
  or _24131_ (_02267_, _02266_, _02264_);
  or _24132_ (_02692_, _02267_, _02260_);
  and _24133_ (_02268_, _01174_, _06631_);
  nand _24134_ (_02269_, _02268_, _05872_);
  or _24135_ (_02270_, _02268_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _24136_ (_02271_, _02270_, _05794_);
  and _24137_ (_02272_, _02271_, _02269_);
  nand _24138_ (_02273_, _01180_, _06088_);
  or _24139_ (_02274_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _24140_ (_02275_, _02274_, _05806_);
  and _24141_ (_02276_, _02275_, _02273_);
  and _24142_ (_02277_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _24143_ (_02278_, _02277_, rst);
  or _24144_ (_02279_, _02278_, _02276_);
  or _24145_ (_02694_, _02279_, _02272_);
  or _24146_ (_02280_, _01988_, _05782_);
  or _24147_ (_02281_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _24148_ (_02282_, _02281_, _05794_);
  and _24149_ (_02283_, _02282_, _02280_);
  and _24150_ (_02284_, _01987_, _06799_);
  not _24151_ (_02285_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor _24152_ (_02286_, _01987_, _02285_);
  or _24153_ (_02287_, _02286_, _02284_);
  and _24154_ (_02288_, _02287_, _05806_);
  nor _24155_ (_02289_, _05793_, _02285_);
  or _24156_ (_02290_, _02289_, rst);
  or _24157_ (_02291_, _02290_, _02288_);
  or _24158_ (_02696_, _02291_, _02283_);
  and _24159_ (_02292_, _01996_, _10208_);
  nand _24160_ (_02293_, _02292_, _05872_);
  or _24161_ (_02294_, _02292_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _24162_ (_02295_, _02294_, _05794_);
  and _24163_ (_02296_, _02295_, _02293_);
  nand _24164_ (_02297_, _02002_, _05334_);
  or _24165_ (_02298_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _24166_ (_02299_, _02298_, _05806_);
  and _24167_ (_02300_, _02299_, _02297_);
  and _24168_ (_02301_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _24169_ (_02302_, _02301_, rst);
  or _24170_ (_02303_, _02302_, _02300_);
  or _24171_ (_02698_, _02303_, _02296_);
  and _24172_ (_02304_, _01996_, _06472_);
  nand _24173_ (_02305_, _02304_, _05872_);
  or _24174_ (_02306_, _02304_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _24175_ (_02307_, _02306_, _05794_);
  and _24176_ (_02308_, _02307_, _02305_);
  nand _24177_ (_02309_, _02002_, _06229_);
  or _24178_ (_02310_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _24179_ (_02311_, _02310_, _05806_);
  and _24180_ (_02312_, _02311_, _02309_);
  and _24181_ (_02313_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _24182_ (_02314_, _02313_, rst);
  or _24183_ (_02315_, _02314_, _02312_);
  or _24184_ (_02700_, _02315_, _02308_);
  nand _24185_ (_02316_, _02040_, _05805_);
  or _24186_ (_02317_, _02316_, _05782_);
  or _24187_ (_02318_, _02046_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _24188_ (_02319_, _02318_, _05794_);
  and _24189_ (_02320_, _02319_, _02317_);
  nand _24190_ (_02321_, _02046_, _06798_);
  and _24191_ (_02322_, _02318_, _05806_);
  and _24192_ (_02323_, _02322_, _02321_);
  not _24193_ (_02324_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor _24194_ (_02325_, _05793_, _02324_);
  or _24195_ (_02326_, _02325_, rst);
  or _24196_ (_02327_, _02326_, _02323_);
  or _24197_ (_02702_, _02327_, _02320_);
  and _24198_ (_02328_, _01981_, _05488_);
  nand _24199_ (_02329_, _02328_, _05872_);
  or _24200_ (_02330_, _02328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _24201_ (_02331_, _02330_, _05794_);
  and _24202_ (_02332_, _02331_, _02329_);
  nor _24203_ (_02333_, _01988_, _05841_);
  and _24204_ (_02334_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _24205_ (_02335_, _02334_, _02333_);
  and _24206_ (_02336_, _02335_, _05806_);
  and _24207_ (_02337_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _24208_ (_02338_, _02337_, rst);
  or _24209_ (_02339_, _02338_, _02336_);
  or _24210_ (_02704_, _02339_, _02332_);
  and _24211_ (_02340_, _02040_, _08133_);
  nand _24212_ (_02341_, _02340_, _05872_);
  or _24213_ (_02342_, _02340_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _24214_ (_02343_, _02342_, _05794_);
  and _24215_ (_02344_, _02343_, _02341_);
  nor _24216_ (_02345_, _02047_, _06054_);
  and _24217_ (_02346_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _24218_ (_02347_, _02346_, _02345_);
  and _24219_ (_02348_, _02347_, _05806_);
  and _24220_ (_02349_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _24221_ (_02350_, _02349_, rst);
  or _24222_ (_02351_, _02350_, _02348_);
  or _24223_ (_02707_, _02351_, _02344_);
  and _24224_ (_02352_, _02040_, _06631_);
  nand _24225_ (_02353_, _02352_, _05872_);
  or _24226_ (_02354_, _02352_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _24227_ (_02355_, _02354_, _05794_);
  and _24228_ (_02356_, _02355_, _02353_);
  nor _24229_ (_02357_, _02047_, _06088_);
  and _24230_ (_02358_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _24231_ (_02359_, _02358_, _02357_);
  and _24232_ (_02360_, _02359_, _05806_);
  and _24233_ (_02361_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _24234_ (_02362_, _02361_, rst);
  or _24235_ (_02363_, _02362_, _02360_);
  or _24236_ (_02709_, _02363_, _02356_);
  and _24237_ (_02364_, _07034_, _05997_);
  nand _24238_ (_02365_, _05997_, _05337_);
  and _24239_ (_02366_, _02365_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or _24240_ (_02367_, _02366_, _02364_);
  and _24241_ (_02738_, _02367_, _05110_);
  and _24242_ (_02368_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not _24243_ (_02369_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _24244_ (_02370_, pc_log_change, _02369_);
  or _24245_ (_02371_, _02370_, _02368_);
  and _24246_ (_02755_, _02371_, _05110_);
  or _24247_ (_02372_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  not _24248_ (_02373_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand _24249_ (_02374_, pc_log_change, _02373_);
  and _24250_ (_02375_, _02374_, _05110_);
  and _24251_ (_02759_, _02375_, _02372_);
  or _24252_ (_02376_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  not _24253_ (_02377_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand _24254_ (_02378_, pc_log_change, _02377_);
  and _24255_ (_02379_, _02378_, _05110_);
  and _24256_ (_02762_, _02379_, _02376_);
  and _24257_ (_02380_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _24258_ (_02381_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _24259_ (_02382_, pc_log_change, _02381_);
  or _24260_ (_02383_, _02382_, _02380_);
  and _24261_ (_02763_, _02383_, _05110_);
  and _24262_ (_02384_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _24263_ (_02385_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _24264_ (_02386_, pc_log_change, _02385_);
  or _24265_ (_02387_, _02386_, _02384_);
  and _24266_ (_02771_, _02387_, _05110_);
  or _24267_ (_02388_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _24268_ (_02389_, pc_log_change, _05264_);
  and _24269_ (_02390_, _02389_, _05110_);
  and _24270_ (_02774_, _02390_, _02388_);
  and _24271_ (_02392_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _24272_ (_02393_, pc_log_change, _06162_);
  or _24273_ (_02394_, _02393_, _02392_);
  and _24274_ (_02776_, _02394_, _05110_);
  and _24275_ (_02395_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not _24276_ (_02396_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _24277_ (_02397_, pc_log_change, _02396_);
  or _24278_ (_02398_, _02397_, _02395_);
  and _24279_ (_02780_, _02398_, _05110_);
  or _24280_ (_02399_, _01668_, _07093_);
  and _24281_ (_02400_, _06463_, _06434_);
  or _24282_ (_02401_, _07052_, _02400_);
  or _24283_ (_02402_, _02401_, _02399_);
  or _24284_ (_02403_, _06849_, _06435_);
  and _24285_ (_02404_, _11727_, _06464_);
  or _24286_ (_02405_, _02404_, _02403_);
  and _24287_ (_02406_, _07139_, _11802_);
  or _24288_ (_02408_, _02406_, _12156_);
  and _24289_ (_02409_, _07107_, _06852_);
  and _24290_ (_02410_, _11729_, _06464_);
  or _24291_ (_02411_, _02410_, _02409_);
  or _24292_ (_02412_, _02411_, _02408_);
  or _24293_ (_02413_, _02412_, _02405_);
  or _24294_ (_02414_, _02413_, _02402_);
  or _24295_ (_02415_, _13078_, _12134_);
  or _24296_ (_02416_, _01664_, _06439_);
  or _24297_ (_02417_, _02416_, _01648_);
  or _24298_ (_02418_, _02417_, _02415_);
  or _24299_ (_02419_, _07126_, _07089_);
  or _24300_ (_02420_, _02419_, _07041_);
  or _24301_ (_02421_, _07131_, _07106_);
  or _24302_ (_02422_, _02421_, _02420_);
  or _24303_ (_02424_, _01665_, _06867_);
  or _24304_ (_02425_, _01670_, _01712_);
  or _24305_ (_02426_, _02425_, _02424_);
  or _24306_ (_02427_, _02426_, _01650_);
  or _24307_ (_02428_, _02427_, _02422_);
  or _24308_ (_02429_, _02428_, _02418_);
  or _24309_ (_02430_, _02429_, _02414_);
  and _24310_ (_02431_, _02430_, _05474_);
  and _24311_ (_02432_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _24312_ (_02433_, _00489_);
  and _24313_ (_02434_, _02433_, _06240_);
  or _24314_ (_02435_, _07056_, _02434_);
  or _24315_ (_02436_, _02435_, _02432_);
  or _24316_ (_02437_, _02436_, _02431_);
  and _24317_ (_02812_, _02437_, _05110_);
  or _24318_ (_02438_, _06453_, _06435_);
  or _24319_ (_02439_, _02438_, _07139_);
  or _24320_ (_02440_, _07108_, _07041_);
  or _24321_ (_02441_, _02440_, _02439_);
  or _24322_ (_02442_, _02441_, _01650_);
  or _24323_ (_02443_, _11756_, _11297_);
  and _24324_ (_02444_, _13086_, _06827_);
  and _24325_ (_02445_, _12149_, _06448_);
  or _24326_ (_02446_, _02445_, _02444_);
  or _24327_ (_02447_, _02446_, _02443_);
  or _24328_ (_02448_, _02447_, _02402_);
  or _24329_ (_02449_, _02448_, _02442_);
  or _24330_ (_02450_, _02449_, _02418_);
  and _24331_ (_02451_, _02450_, _05474_);
  and _24332_ (_02452_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _24333_ (_02453_, _02452_, _02435_);
  or _24334_ (_02454_, _02453_, _02451_);
  and _24335_ (_02814_, _02454_, _05110_);
  and _24336_ (_02455_, _06901_, _08224_);
  and _24337_ (_02456_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _24338_ (_02457_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and _24339_ (_02458_, _02457_, _06011_);
  or _24340_ (_02459_, _02458_, _02456_);
  or _24341_ (_02460_, _02459_, _02455_);
  and _24342_ (_02820_, _02460_, _05110_);
  or _24343_ (_02461_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  not _24344_ (_02462_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _24345_ (_02464_, pc_log_change, _02462_);
  and _24346_ (_02465_, _02464_, _05110_);
  and _24347_ (_02825_, _02465_, _02461_);
  and _24348_ (_02467_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _24349_ (_02468_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _24350_ (_02469_, pc_log_change, _02468_);
  or _24351_ (_02470_, _02469_, _02467_);
  and _24352_ (_02828_, _02470_, _05110_);
  or _24353_ (_02471_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand _24354_ (_02473_, _06205_, _07553_);
  and _24355_ (_02474_, _02473_, _05110_);
  and _24356_ (_02834_, _02474_, _02471_);
  and _24357_ (_02475_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not _24358_ (_02477_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _24359_ (_02478_, pc_log_change, _02477_);
  or _24360_ (_02479_, _02478_, _02475_);
  and _24361_ (_02837_, _02479_, _05110_);
  and _24362_ (_02480_, _06807_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and _24363_ (_02481_, _06825_, _06448_);
  or _24364_ (_02482_, _02481_, _01645_);
  or _24365_ (_02483_, _02482_, _11738_);
  or _24366_ (_02484_, _02483_, _06951_);
  and _24367_ (_02485_, _06820_, _06448_);
  or _24368_ (_02486_, _02485_, _06939_);
  or _24369_ (_02487_, _11742_, _11754_);
  or _24370_ (_02488_, _02487_, _02486_);
  or _24371_ (_02489_, _07045_, _06458_);
  or _24372_ (_02490_, _02489_, _02404_);
  and _24373_ (_02491_, _11727_, _06448_);
  and _24374_ (_02492_, _07044_, _06276_);
  or _24375_ (_02493_, _02492_, _02491_);
  or _24376_ (_02494_, _02493_, _02490_);
  and _24377_ (_02495_, _11727_, _06431_);
  or _24378_ (_02496_, _02495_, _07041_);
  or _24379_ (_02497_, _07111_, _07052_);
  or _24380_ (_02498_, _02497_, _02496_);
  or _24381_ (_02499_, _02498_, _02494_);
  or _24382_ (_02500_, _02499_, _02488_);
  or _24383_ (_02501_, _02500_, _02484_);
  and _24384_ (_02502_, _02501_, _06842_);
  or _24385_ (_02848_, _02502_, _02480_);
  and _24386_ (_02504_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not _24387_ (_02505_, pc_log_change);
  and _24388_ (_02506_, _02505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or _24389_ (_02507_, _02506_, _02504_);
  and _24390_ (_02850_, _02507_, _05110_);
  or _24391_ (_02508_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  not _24392_ (_02509_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _24393_ (_02510_, pc_log_change, _02509_);
  and _24394_ (_02511_, _02510_, _05110_);
  and _24395_ (_02861_, _02511_, _02508_);
  and _24396_ (_02512_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _24397_ (_02513_, pc_log_change, _02509_);
  or _24398_ (_02514_, _02513_, _02512_);
  and _24399_ (_02863_, _02514_, _05110_);
  or _24400_ (_02515_, _06461_, _06457_);
  or _24401_ (_02516_, _07081_, _06465_);
  or _24402_ (_02517_, _02516_, _02515_);
  or _24403_ (_02519_, _11293_, _06449_);
  or _24404_ (_02521_, _02519_, _02517_);
  and _24405_ (_02523_, _07080_, _06460_);
  or _24406_ (_02524_, _01668_, _01645_);
  nor _24407_ (_02526_, _02524_, _02523_);
  nand _24408_ (_02527_, _02526_, _01836_);
  or _24409_ (_02528_, _02527_, _02521_);
  or _24410_ (_02529_, _02491_, _02485_);
  or _24411_ (_02530_, _02410_, _12156_);
  or _24412_ (_02531_, _02530_, _02529_);
  or _24413_ (_02532_, _02531_, _07091_);
  or _24414_ (_02533_, _02532_, _02405_);
  or _24415_ (_02534_, _02533_, _02528_);
  and _24416_ (_02535_, _02534_, _06842_);
  nor _24417_ (_02536_, _06870_, rst);
  and _24418_ (_02537_, _02536_, _06435_);
  and _24419_ (_02538_, _06807_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or _24420_ (_02539_, _02538_, _02537_);
  or _24421_ (_02875_, _02539_, _02535_);
  nand _24422_ (_02540_, _08288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _24423_ (_02541_, _02540_, _08274_);
  and _24424_ (_02542_, _08274_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _24425_ (_02544_, _02542_, _02541_);
  and _24426_ (_02878_, _02544_, _05110_);
  nand _24427_ (_02545_, _01836_, _11299_);
  or _24428_ (_02546_, _01667_, _07092_);
  or _24429_ (_02548_, _02546_, _02415_);
  or _24430_ (_02550_, _02548_, _02545_);
  and _24431_ (_02551_, _07038_, _06448_);
  or _24432_ (_02552_, _02489_, _01649_);
  or _24433_ (_02554_, _02552_, _02551_);
  or _24434_ (_02556_, _07052_, _06828_);
  or _24435_ (_02558_, _11737_, _07097_);
  or _24436_ (_02560_, _02558_, _02556_);
  or _24437_ (_02561_, _02560_, _02554_);
  or _24438_ (_02563_, _01664_, _07121_);
  or _24439_ (_02564_, _02563_, _02481_);
  or _24440_ (_02566_, _02564_, _06822_);
  or _24441_ (_02567_, _02566_, _02561_);
  or _24442_ (_02568_, _02567_, _02550_);
  and _24443_ (_02569_, _02568_, _05474_);
  and _24444_ (_02570_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _24445_ (_02571_, _06435_, _05151_);
  or _24446_ (_02572_, _02571_, _02570_);
  or _24447_ (_02573_, _02572_, _02569_);
  and _24448_ (_02881_, _02573_, _05110_);
  and _24449_ (_02574_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _24450_ (_02575_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or _24451_ (_02576_, _02575_, _02574_);
  and _24452_ (_02885_, _02576_, _05110_);
  and _24453_ (_02577_, _06807_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  or _24454_ (_02579_, _06460_, _06448_);
  and _24455_ (_02580_, _02579_, _06814_);
  or _24456_ (_02581_, _02546_, _02487_);
  or _24457_ (_02582_, _02581_, _02580_);
  or _24458_ (_02583_, _01649_, _06462_);
  and _24459_ (_02584_, _06946_, _06810_);
  or _24460_ (_02585_, _01647_, _02584_);
  or _24461_ (_02586_, _02585_, _02583_);
  or _24462_ (_02588_, _12089_, _06439_);
  or _24463_ (_02589_, _01665_, _07139_);
  or _24464_ (_02590_, _02589_, _02588_);
  or _24465_ (_02591_, _02590_, _06819_);
  or _24466_ (_02592_, _02591_, _02586_);
  or _24467_ (_02593_, _02592_, _02564_);
  or _24468_ (_02594_, _02593_, _02582_);
  or _24469_ (_02595_, _06439_, _05473_);
  nor _24470_ (_02596_, \oc8051_top_1.oc8051_sfr1.wait_data , rst);
  and _24471_ (_02597_, _02596_, _02595_);
  and _24472_ (_02598_, _02597_, _02594_);
  or _24473_ (_02894_, _02598_, _02577_);
  or _24474_ (_02599_, _09328_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand _24475_ (_02600_, _09328_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _24476_ (_02601_, _02600_, _02599_);
  nand _24477_ (_02603_, _02601_, _05110_);
  nor _24478_ (_02897_, _02603_, _08274_);
  nor _24479_ (_02604_, _05901_, _06010_);
  and _24480_ (_02605_, _06010_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _24481_ (_02606_, _02605_, _05995_);
  or _24482_ (_02608_, _02606_, _02604_);
  or _24483_ (_02609_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _24484_ (_02610_, _02609_, _05110_);
  and _24485_ (_02906_, _02610_, _02608_);
  nand _24486_ (_02611_, _06673_, _05901_);
  or _24487_ (_02612_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _24488_ (_02613_, _02612_, _05110_);
  and _24489_ (_02917_, _02613_, _02611_);
  and _24490_ (_02614_, _01996_, _05867_);
  nand _24491_ (_02615_, _02614_, _05872_);
  or _24492_ (_02616_, _02614_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _24493_ (_02617_, _02616_, _05794_);
  and _24494_ (_02618_, _02617_, _02615_);
  nand _24495_ (_02619_, _02002_, _05901_);
  or _24496_ (_02620_, _02002_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _24497_ (_02621_, _02620_, _05806_);
  and _24498_ (_02622_, _02621_, _02619_);
  and _24499_ (_02623_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _24500_ (_02624_, _02623_, rst);
  or _24501_ (_02625_, _02624_, _02622_);
  or _24502_ (_02921_, _02625_, _02618_);
  nand _24503_ (_02627_, _06673_, _05841_);
  or _24504_ (_02628_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _24505_ (_02629_, _02628_, _05110_);
  and _24506_ (_02925_, _02629_, _02627_);
  and _24507_ (_02630_, _06807_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or _24508_ (_02631_, _02556_, _11738_);
  or _24509_ (_02632_, _02631_, _02482_);
  or _24510_ (_02633_, _12134_, _11761_);
  or _24511_ (_02634_, _13072_, _02491_);
  or _24512_ (_02635_, _02634_, _02633_);
  or _24513_ (_02636_, _02635_, _07050_);
  or _24514_ (_02637_, _02636_, _02488_);
  or _24515_ (_02638_, _02637_, _02632_);
  and _24516_ (_02639_, _02638_, _06842_);
  or _24517_ (_02940_, _02639_, _02630_);
  or _24518_ (_02640_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand _24519_ (_02641_, _06205_, _12002_);
  and _24520_ (_02642_, _02641_, _05110_);
  and _24521_ (_02946_, _02642_, _02640_);
  and _24522_ (_02948_, _01725_, _05110_);
  nand _24523_ (_02643_, _06560_, _06088_);
  or _24524_ (_02644_, _06560_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and _24525_ (_02645_, _02644_, _05110_);
  and _24526_ (_02954_, _02645_, _02643_);
  and _24527_ (_02646_, _06901_, _12894_);
  and _24528_ (_02647_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _24529_ (_02648_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and _24530_ (_02649_, _02648_, _06011_);
  or _24531_ (_02650_, _02649_, _02647_);
  or _24532_ (_02651_, _02650_, _02646_);
  and _24533_ (_02963_, _02651_, _05110_);
  and _24534_ (_02652_, _08056_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor _24535_ (_02653_, _08056_, _05901_);
  or _24536_ (_02654_, _02653_, _02652_);
  and _24537_ (_02970_, _02654_, _05110_);
  or _24538_ (_02657_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand _24539_ (_02658_, _06205_, _13066_);
  and _24540_ (_02659_, _02658_, _05110_);
  and _24541_ (_03001_, _02659_, _02657_);
  and _24542_ (_02660_, _08056_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _24543_ (_02661_, _07034_, _06001_);
  or _24544_ (_02662_, _02661_, _02660_);
  and _24545_ (_03033_, _02662_, _05110_);
  nor _24546_ (_02663_, _01320_, _05841_);
  and _24547_ (_02664_, _01320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _24548_ (_02665_, _02664_, _02663_);
  and _24549_ (_03057_, _02665_, _05110_);
  and _24550_ (_02667_, _12841_, _08280_);
  and _24551_ (_02669_, _08286_, _12828_);
  and _24552_ (_02670_, _02669_, _12841_);
  not _24553_ (_02672_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _24554_ (_02673_, _08286_, _02672_);
  or _24555_ (_02674_, _02673_, _02670_);
  and _24556_ (_02675_, _02674_, _08282_);
  nand _24557_ (_02676_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _24558_ (_02678_, _02676_, _08281_);
  nor _24559_ (_02679_, _02678_, _02675_);
  nor _24560_ (_02680_, _02679_, _08280_);
  or _24561_ (_02681_, _02680_, _02667_);
  nand _24562_ (_02682_, _02681_, _05110_);
  nor _24563_ (_03059_, _02682_, _08274_);
  and _24564_ (_03064_, _11832_, _05110_);
  and _24565_ (_03073_, _12252_, _05110_);
  and _24566_ (_03075_, _12220_, _05110_);
  nand _24567_ (_02683_, _02670_, _08281_);
  nand _24568_ (_02684_, _02683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _24569_ (_02685_, _02684_, _02667_);
  or _24570_ (_02686_, _02685_, _08274_);
  and _24571_ (_03085_, _02686_, _05110_);
  and _24572_ (_03089_, _12291_, _05110_);
  nor _24573_ (_03101_, _12014_, rst);
  and _24574_ (_02687_, _10641_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _24575_ (_03108_, _02687_, _10460_);
  and _24576_ (_02689_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _24577_ (_02691_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or _24578_ (_03112_, _02691_, _02689_);
  not _24579_ (_02693_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  and _24580_ (_02695_, _01326_, _02693_);
  and _24581_ (_02697_, _02695_, _08752_);
  or _24582_ (_02699_, _02697_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not _24583_ (_02701_, rxd_i);
  nand _24584_ (_02703_, _02697_, _02701_);
  and _24585_ (_02705_, _02703_, _05110_);
  and _24586_ (_03114_, _02705_, _02699_);
  and _24587_ (_02706_, _01140_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _24588_ (_02708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _05850_);
  nor _24589_ (_02710_, _02708_, _05987_);
  not _24590_ (_02711_, _02710_);
  and _24591_ (_02712_, _02711_, _06099_);
  or _24592_ (_02713_, _02712_, _05986_);
  or _24593_ (_02714_, _02713_, _02706_);
  or _24594_ (_02715_, _02710_, _06137_);
  and _24595_ (_02716_, _02715_, _05110_);
  and _24596_ (_03130_, _02716_, _02714_);
  and _24597_ (_02717_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _24598_ (_02718_, _08235_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _24599_ (_02719_, _02718_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _24600_ (_02720_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _24601_ (_02721_, _02720_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _24602_ (_02722_, _02693_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _24603_ (_02723_, _02722_, _02721_);
  and _24604_ (_02724_, _02723_, _08745_);
  nor _24605_ (_02725_, _02724_, _02719_);
  nor _24606_ (_02726_, _02725_, _01050_);
  nor _24607_ (_02727_, _02723_, _01325_);
  and _24608_ (_02728_, _08742_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _24609_ (_02729_, _08235_, _01057_);
  and _24610_ (_02730_, _02729_, _02728_);
  nor _24611_ (_02731_, _02730_, _08745_);
  not _24612_ (_02732_, _02731_);
  nor _24613_ (_02733_, _02732_, _08748_);
  nor _24614_ (_02734_, _02733_, _02727_);
  not _24615_ (_02735_, _02719_);
  nand _24616_ (_02736_, _02735_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nor _24617_ (_02737_, _02736_, _02734_);
  or _24618_ (_02739_, _02737_, _02726_);
  and _24619_ (_02740_, _02739_, _09325_);
  or _24620_ (_03135_, _02740_, _02717_);
  not _24621_ (_02741_, _02725_);
  and _24622_ (_02742_, _02741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nand _24623_ (_02743_, _02735_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor _24624_ (_02744_, _02743_, _02734_);
  or _24625_ (_02745_, _02744_, _02742_);
  and _24626_ (_02746_, _02745_, _09325_);
  or _24627_ (_03143_, _02746_, _09324_);
  and _24628_ (_02747_, _02741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _24629_ (_02748_, _02727_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _24630_ (_02749_, _08748_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _24631_ (_02750_, _02749_, _02731_);
  or _24632_ (_02751_, _02750_, _02748_);
  and _24633_ (_02752_, _02751_, _02735_);
  or _24634_ (_02753_, _02752_, _02747_);
  and _24635_ (_02754_, _02753_, _09325_);
  or _24636_ (_03145_, _02754_, _01065_);
  or _24637_ (_02756_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _24638_ (_02757_, _02756_, _02734_);
  or _24639_ (_02758_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _24640_ (_02760_, _02758_, _09325_);
  and _24641_ (_02761_, _02760_, _02757_);
  or _24642_ (_03147_, _02761_, _01195_);
  or _24643_ (_02764_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _24644_ (_02765_, _02764_, _02734_);
  or _24645_ (_02766_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _24646_ (_02767_, _02766_, _09325_);
  and _24647_ (_02768_, _02767_, _02765_);
  or _24648_ (_03149_, _02768_, _01197_);
  or _24649_ (_02769_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _24650_ (_02770_, _02769_, _02734_);
  or _24651_ (_02772_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and _24652_ (_02773_, _02772_, _09325_);
  and _24653_ (_02775_, _02773_, _02770_);
  or _24654_ (_03151_, _02775_, _01199_);
  or _24655_ (_02777_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _24656_ (_02778_, _02777_, _02734_);
  or _24657_ (_02779_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _24658_ (_02781_, _02779_, _09325_);
  and _24659_ (_02782_, _02781_, _02778_);
  or _24660_ (_03153_, _02782_, _01979_);
  not _24661_ (_02783_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _24662_ (_02784_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not _24663_ (_02785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _24664_ (_02786_, _05846_, _02785_);
  or _24665_ (_02787_, _02786_, _11265_);
  nor _24666_ (_02788_, _02787_, _02784_);
  nand _24667_ (_02789_, _02788_, _02783_);
  nor _24668_ (_02790_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor _24669_ (_02791_, _02790_, _02788_);
  nand _24670_ (_02792_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _24671_ (_02793_, _02792_, _02791_);
  and _24672_ (_02794_, _02793_, _05110_);
  and _24673_ (_03155_, _02794_, _02789_);
  or _24674_ (_02795_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _24675_ (_02796_, _02795_, _02734_);
  or _24676_ (_02797_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _24677_ (_02798_, _02797_, _09325_);
  and _24678_ (_02799_, _02798_, _02796_);
  or _24679_ (_03165_, _02799_, _02689_);
  or _24680_ (_02800_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _24681_ (_02801_, _02800_, _02734_);
  and _24682_ (_02802_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _24683_ (_02803_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _24684_ (_02804_, _02803_, _09325_);
  or _24685_ (_02805_, _02804_, _02802_);
  and _24686_ (_03167_, _02805_, _02801_);
  or _24687_ (_02806_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _24688_ (_02807_, _02806_, _02734_);
  and _24689_ (_02808_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _24690_ (_02809_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  and _24691_ (_02810_, _02809_, _09325_);
  or _24692_ (_02811_, _02810_, _02808_);
  and _24693_ (_03170_, _02811_, _02807_);
  or _24694_ (_02813_, _02719_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _24695_ (_02815_, _02813_, _02734_);
  and _24696_ (_02816_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _24697_ (_02817_, _02725_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  and _24698_ (_02818_, _02817_, _09325_);
  or _24699_ (_02819_, _02818_, _02816_);
  and _24700_ (_03173_, _02819_, _02815_);
  and _24701_ (_03186_, _02791_, _05110_);
  nor _24702_ (_02821_, _02734_, _01050_);
  and _24703_ (_02822_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  or _24704_ (_02823_, _02822_, rxd_i);
  or _24705_ (_02824_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  and _24706_ (_02826_, _02824_, _02724_);
  or _24707_ (_02827_, _02826_, _02719_);
  and _24708_ (_02829_, _02827_, _02823_);
  or _24709_ (_02830_, _02829_, _02821_);
  nand _24710_ (_02831_, _02719_, _02701_);
  and _24711_ (_02832_, _02831_, _09325_);
  and _24712_ (_02833_, _02832_, _02830_);
  and _24713_ (_02835_, _09323_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _24714_ (_03191_, _02835_, _02833_);
  and _24715_ (_02836_, _09325_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or _24716_ (_03193_, _02836_, _02717_);
  or _24717_ (_02838_, _12171_, _05782_);
  nor _24718_ (_02839_, _12172_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _24719_ (_02840_, _02839_, _10157_);
  and _24720_ (_02841_, _02840_, _02838_);
  or _24721_ (_02842_, _02841_, _10162_);
  and _24722_ (_02843_, _12083_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _24723_ (_02844_, _02843_, _01548_);
  and _24724_ (_02845_, _02844_, _10157_);
  or _24725_ (_02846_, _02845_, _02842_);
  nand _24726_ (_02847_, _10162_, _05901_);
  and _24727_ (_02849_, _02847_, _05110_);
  and _24728_ (_03196_, _02849_, _02846_);
  and _24729_ (_03198_, _12049_, _05110_);
  and _24730_ (_03203_, _11909_, _05110_);
  and _24731_ (_02851_, _07204_, _06613_);
  nor _24732_ (_02852_, _10208_, _05142_);
  or _24733_ (_02853_, _02852_, _10209_);
  and _24734_ (_02854_, _06638_, _08132_);
  nand _24735_ (_02855_, _02854_, _02853_);
  nor _24736_ (_02856_, _07235_, _06622_);
  and _24737_ (_02857_, _12179_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _24738_ (_02858_, _02857_, _02856_);
  nand _24739_ (_02859_, _02858_, _02855_);
  and _24740_ (_02860_, _02859_, _06637_);
  or _24741_ (_02862_, _02860_, _02851_);
  and _24742_ (_03309_, _02862_, _05110_);
  and _24743_ (_02864_, _06007_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _24744_ (_02865_, _05337_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and _24745_ (_02866_, _02865_, _06011_);
  and _24746_ (_02867_, _06799_, _06901_);
  or _24747_ (_02868_, _02867_, _02866_);
  or _24748_ (_02869_, _02868_, _02864_);
  and _24749_ (_03316_, _02869_, _05110_);
  or _24750_ (_02870_, _01327_, _08750_);
  and _24751_ (_02871_, _02870_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _24752_ (_02872_, _02871_, _02697_);
  and _24753_ (_03532_, _02872_, _05110_);
  and _24754_ (_02873_, _08615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _24755_ (_02874_, _08617_, _06183_);
  or _24756_ (_02876_, _02874_, _02873_);
  and _24757_ (_03534_, _02876_, _05110_);
  not _24758_ (_02877_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _24759_ (_02879_, _02722_, _08753_);
  and _24760_ (_02880_, _02879_, _08752_);
  nor _24761_ (_02882_, _02880_, _02877_);
  and _24762_ (_02883_, _02880_, rxd_i);
  or _24763_ (_02884_, _02883_, _02882_);
  and _24764_ (_03571_, _02884_, _05110_);
  and _24765_ (_02886_, _01981_, _05867_);
  nand _24766_ (_02887_, _02886_, _05872_);
  or _24767_ (_02888_, _02886_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _24768_ (_02889_, _02888_, _05794_);
  and _24769_ (_02890_, _02889_, _02887_);
  nor _24770_ (_02891_, _01988_, _05901_);
  and _24771_ (_02892_, _01988_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _24772_ (_02893_, _02892_, _02891_);
  and _24773_ (_02895_, _02893_, _05806_);
  and _24774_ (_02896_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _24775_ (_02898_, _02896_, rst);
  or _24776_ (_02899_, _02898_, _02895_);
  or _24777_ (_03593_, _02899_, _02890_);
  and _24778_ (_02900_, _02040_, _05867_);
  nand _24779_ (_02901_, _02900_, _05872_);
  or _24780_ (_02902_, _02900_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _24781_ (_02903_, _02902_, _05794_);
  and _24782_ (_02904_, _02903_, _02901_);
  nor _24783_ (_02905_, _02047_, _05901_);
  and _24784_ (_02907_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _24785_ (_02908_, _02907_, _02905_);
  and _24786_ (_02909_, _02908_, _05806_);
  and _24787_ (_02910_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _24788_ (_02911_, _02910_, rst);
  or _24789_ (_02912_, _02911_, _02909_);
  or _24790_ (_03596_, _02912_, _02904_);
  not _24791_ (_02913_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _24792_ (_02914_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and _24793_ (_02915_, _02914_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  not _24794_ (_02916_, _02915_);
  nor _24795_ (_02918_, _08235_, _08741_);
  and _24796_ (_02919_, _02918_, _02916_);
  and _24797_ (_02920_, _02919_, _01325_);
  nor _24798_ (_02922_, _02920_, _02913_);
  and _24799_ (_02923_, _02920_, rxd_i);
  or _24800_ (_02924_, _02923_, rst);
  or _24801_ (_03599_, _02924_, _02922_);
  nor _24802_ (_02926_, _08235_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _24803_ (_02927_, _02926_, _08745_);
  nor _24804_ (_02928_, _02724_, _08741_);
  or _24805_ (_02929_, _02928_, _02927_);
  and _24806_ (_02930_, _02929_, _02735_);
  nand _24807_ (_02931_, _02741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _24808_ (_02932_, _02931_, _09325_);
  or _24809_ (_03659_, _02932_, _02930_);
  or _24810_ (_02933_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nand _24811_ (_02934_, pc_log_change, _00990_);
  and _24812_ (_02935_, _02934_, _05110_);
  and _24813_ (_03660_, _02935_, _02933_);
  and _24814_ (_02936_, _08617_, _08224_);
  nor _24815_ (_02937_, _06004_, _05995_);
  or _24816_ (_02938_, _02937_, _08614_);
  and _24817_ (_02939_, _02938_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or _24818_ (_02941_, _02939_, _02936_);
  and _24819_ (_03663_, _02941_, _05110_);
  and _24820_ (_02942_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _24821_ (_02943_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _24822_ (_02944_, pc_log_change, _02943_);
  or _24823_ (_02945_, _02944_, _02942_);
  and _24824_ (_03670_, _02945_, _05110_);
  and _24825_ (_02947_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _24826_ (_02949_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _24827_ (_02950_, _02949_, _02947_);
  and _24828_ (_02951_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _24829_ (_02952_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _24830_ (_02953_, _02952_, _02951_);
  or _24831_ (_02955_, _02953_, _02950_);
  and _24832_ (_02956_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _24833_ (_02957_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _24834_ (_02958_, _02957_, _02956_);
  and _24835_ (_02959_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _24836_ (_02960_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _24837_ (_02961_, _02960_, _02959_);
  or _24838_ (_02962_, _02961_, _02958_);
  or _24839_ (_02964_, _02962_, _02955_);
  and _24840_ (_02965_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _24841_ (_02966_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _24842_ (_02967_, _02966_, _02965_);
  and _24843_ (_02968_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _24844_ (_02969_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _24845_ (_02971_, _02969_, _02968_);
  or _24846_ (_02972_, _02971_, _02967_);
  and _24847_ (_02973_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _24848_ (_02974_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _24849_ (_02975_, _02974_, _02973_);
  and _24850_ (_02976_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _24851_ (_02977_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or _24852_ (_02978_, _02977_, _02976_);
  or _24853_ (_02979_, _02978_, _02975_);
  or _24854_ (_02980_, _02979_, _02972_);
  or _24855_ (_02981_, _02980_, _02964_);
  and _24856_ (_02982_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _24857_ (_02983_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _24858_ (_02984_, _02983_, _02982_);
  and _24859_ (_02985_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _24860_ (_02986_, _01819_, _12029_);
  or _24861_ (_02987_, _02986_, _02985_);
  or _24862_ (_02988_, _02987_, _02984_);
  or _24863_ (_02989_, _01846_, p2_in[6]);
  or _24864_ (_02990_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _24865_ (_02991_, _02990_, _02989_);
  and _24866_ (_02992_, _02991_, _01853_);
  or _24867_ (_02993_, _01846_, p3_in[6]);
  or _24868_ (_02994_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _24869_ (_02995_, _02994_, _02993_);
  and _24870_ (_02996_, _02995_, _01830_);
  or _24871_ (_02997_, _02996_, _02992_);
  or _24872_ (_02998_, _01846_, p1_in[6]);
  or _24873_ (_02999_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _24874_ (_03000_, _02999_, _02998_);
  and _24875_ (_03002_, _03000_, _01865_);
  or _24876_ (_03003_, _01846_, p0_in[6]);
  or _24877_ (_03004_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _24878_ (_03005_, _03004_, _03003_);
  and _24879_ (_03006_, _03005_, _01859_);
  or _24880_ (_03007_, _03006_, _03002_);
  or _24881_ (_03008_, _03007_, _02997_);
  or _24882_ (_03009_, _03008_, _02988_);
  and _24883_ (_03010_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _24884_ (_03011_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _24885_ (_03012_, _03011_, _03010_);
  or _24886_ (_03013_, _03012_, _03009_);
  or _24887_ (_03014_, _03013_, _02981_);
  and _24888_ (_03015_, _03014_, _01893_);
  and _24889_ (_03016_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or _24890_ (_03017_, _03016_, _03015_);
  or _24891_ (_03018_, _03017_, _01732_);
  nand _24892_ (_03019_, _01732_, _06780_);
  and _24893_ (_03020_, _03019_, _05110_);
  and _24894_ (_03684_, _03020_, _03018_);
  or _24895_ (_03021_, _02913_, rxd_i);
  nand _24896_ (_03022_, _03021_, _08746_);
  or _24897_ (_03023_, _08748_, _08743_);
  and _24898_ (_03024_, _03023_, _03022_);
  or _24899_ (_03025_, _02732_, _02718_);
  or _24900_ (_03026_, _03025_, _03024_);
  and _24901_ (_03686_, _03026_, _09325_);
  not _24902_ (_03027_, _06239_);
  and _24903_ (_03028_, _12095_, _03027_);
  or _24904_ (_03029_, _11730_, _07111_);
  or _24905_ (_03030_, _03029_, _11761_);
  or _24906_ (_03031_, _03030_, _02487_);
  or _24907_ (_03032_, _03031_, _11740_);
  and _24908_ (_03034_, _03032_, _06870_);
  or _24909_ (_03035_, _03034_, _03028_);
  and _24910_ (_03704_, _03035_, _05110_);
  nor _24911_ (_03036_, _01722_, rst);
  nand _24912_ (_03037_, _01721_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or _24913_ (_03038_, _01721_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _24914_ (_03039_, _03038_, _03037_);
  and _24915_ (_03706_, _03039_, _03036_);
  nor _24916_ (_03040_, _06229_, _05465_);
  and _24917_ (_03041_, _08329_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or _24918_ (_03042_, _03041_, _03040_);
  and _24919_ (_03709_, _03042_, _05110_);
  nor _24920_ (_03724_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  nand _24921_ (_03043_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand _24922_ (_03044_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _24923_ (_03045_, _03044_, _03043_);
  or _24924_ (_03046_, _01910_, _11600_);
  or _24925_ (_03047_, _01913_, _06897_);
  and _24926_ (_03048_, _03047_, _03046_);
  and _24927_ (_03049_, _03048_, _03045_);
  or _24928_ (_03050_, _01927_, _11628_);
  or _24929_ (_03051_, _01925_, _05904_);
  and _24930_ (_03052_, _03051_, _03050_);
  nand _24931_ (_03053_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nand _24932_ (_03054_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _24933_ (_03055_, _03054_, _03053_);
  and _24934_ (_03056_, _03055_, _03052_);
  and _24935_ (_03058_, _03056_, _03049_);
  or _24936_ (_03060_, _01936_, _13275_);
  or _24937_ (_03061_, _01935_, _00059_);
  and _24938_ (_03062_, _03061_, _03060_);
  nand _24939_ (_03063_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand _24940_ (_03065_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _24941_ (_03066_, _03065_, _03063_);
  and _24942_ (_03067_, _03066_, _03062_);
  nand _24943_ (_03068_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _24944_ (_03069_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _24945_ (_03070_, _03069_, _03068_);
  nand _24946_ (_03071_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand _24947_ (_03072_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and _24948_ (_03074_, _03072_, _03071_);
  and _24949_ (_03076_, _03074_, _03070_);
  and _24950_ (_03077_, _03076_, _03067_);
  and _24951_ (_03078_, _03077_, _03058_);
  nand _24952_ (_03079_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand _24953_ (_03080_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _24954_ (_03081_, _03080_, _03079_);
  nand _24955_ (_03082_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not _24956_ (_03083_, _12324_);
  nand _24957_ (_03084_, _01819_, _03083_);
  and _24958_ (_03086_, _03084_, _03082_);
  and _24959_ (_03087_, _03086_, _03081_);
  nor _24960_ (_03088_, _01846_, p3_in[0]);
  and _24961_ (_03090_, _01846_, _02324_);
  nor _24962_ (_03091_, _03090_, _03088_);
  nand _24963_ (_03092_, _03091_, _01830_);
  nor _24964_ (_03093_, _01846_, p2_in[0]);
  and _24965_ (_03094_, _01846_, _02285_);
  nor _24966_ (_03095_, _03094_, _03093_);
  nand _24967_ (_03096_, _03095_, _01853_);
  and _24968_ (_03097_, _03096_, _03092_);
  nor _24969_ (_03098_, _01846_, p0_in[0]);
  and _24970_ (_03100_, _01846_, _02251_);
  nor _24971_ (_03102_, _03100_, _03098_);
  nand _24972_ (_03103_, _03102_, _01859_);
  nor _24973_ (_03104_, _01846_, p1_in[0]);
  and _24974_ (_03105_, _01846_, _02089_);
  nor _24975_ (_03106_, _03105_, _03104_);
  nand _24976_ (_03107_, _03106_, _01865_);
  and _24977_ (_03109_, _03107_, _03103_);
  and _24978_ (_03110_, _03109_, _03097_);
  and _24979_ (_03111_, _03110_, _03087_);
  and _24980_ (_03113_, _12179_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _24981_ (_03115_, _06622_, _06512_);
  nor _24982_ (_03116_, _03115_, _03113_);
  and _24983_ (_03117_, _03116_, _06637_);
  nor _24984_ (_03118_, _08272_, _05269_);
  or _24985_ (_03119_, _03118_, _00998_);
  nand _24986_ (_03120_, _03119_, _02854_);
  nand _24987_ (_03121_, _03120_, _03117_);
  or _24988_ (_03122_, _07364_, _06637_);
  nand _24989_ (_03123_, _03122_, _03121_);
  nand _24990_ (_03124_, _03123_, _08312_);
  or _24991_ (_03125_, _03123_, _08312_);
  nand _24992_ (_03126_, _03125_, _03124_);
  not _24993_ (_03127_, _08155_);
  nand _24994_ (_03128_, _03127_, _06672_);
  or _24995_ (_03129_, _03127_, _06672_);
  and _24996_ (_03131_, _03129_, _03128_);
  nand _24997_ (_03132_, _03131_, _03126_);
  or _24998_ (_03133_, _03131_, _03126_);
  nand _24999_ (_03134_, _03133_, _03132_);
  nor _25000_ (_03136_, _06784_, _06746_);
  nand _25001_ (_03137_, _08144_, _03136_);
  or _25002_ (_03138_, _08144_, _03136_);
  and _25003_ (_03139_, _03138_, _03137_);
  nand _25004_ (_03140_, _03139_, _03134_);
  or _25005_ (_03141_, _03139_, _03134_);
  and _25006_ (_03142_, _03141_, _03140_);
  or _25007_ (_03144_, _02862_, _07032_);
  nand _25008_ (_03146_, _02862_, _07032_);
  and _25009_ (_03148_, _03146_, _03144_);
  nand _25010_ (_03150_, _03148_, _03142_);
  or _25011_ (_03152_, _03148_, _03142_);
  nand _25012_ (_03154_, _03152_, _03150_);
  nand _25013_ (_03156_, _03154_, _01874_);
  nand _25014_ (_03157_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _25015_ (_03158_, _03157_, _03156_);
  and _25016_ (_03159_, _03158_, _03111_);
  nand _25017_ (_03160_, _03159_, _03078_);
  and _25018_ (_03161_, _03160_, _01893_);
  and _25019_ (_03162_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or _25020_ (_03163_, _03162_, _01732_);
  or _25021_ (_03164_, _03163_, _03161_);
  nand _25022_ (_03166_, _01732_, _07418_);
  and _25023_ (_03168_, _03166_, _05110_);
  and _25024_ (_03748_, _03168_, _03164_);
  and _25025_ (_03169_, _08615_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and _25026_ (_03171_, _08617_, _12874_);
  or _25027_ (_03172_, _03171_, _03169_);
  and _25028_ (_03755_, _03172_, _05110_);
  and _25029_ (_03174_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _25030_ (_03175_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _25031_ (_03176_, _03175_, _03174_);
  and _25032_ (_03177_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _25033_ (_03178_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _25034_ (_03179_, _03178_, _03177_);
  or _25035_ (_03180_, _03179_, _03176_);
  and _25036_ (_03181_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _25037_ (_03182_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _25038_ (_03183_, _03182_, _03181_);
  and _25039_ (_03184_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _25040_ (_03185_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _25041_ (_03187_, _03185_, _03184_);
  or _25042_ (_03188_, _03187_, _03183_);
  or _25043_ (_03189_, _03188_, _03180_);
  and _25044_ (_03190_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _25045_ (_03192_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _25046_ (_03194_, _03192_, _03190_);
  and _25047_ (_03195_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _25048_ (_03197_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _25049_ (_03199_, _03197_, _03195_);
  or _25050_ (_03200_, _03199_, _03194_);
  and _25051_ (_03201_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and _25052_ (_03202_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _25053_ (_03204_, _03202_, _03201_);
  and _25054_ (_03205_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _25055_ (_03206_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or _25056_ (_03207_, _03206_, _03205_);
  or _25057_ (_03208_, _03207_, _03204_);
  or _25058_ (_03209_, _03208_, _03200_);
  or _25059_ (_03210_, _03209_, _03189_);
  and _25060_ (_03211_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _25061_ (_03212_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or _25062_ (_03213_, _03212_, _03211_);
  and _25063_ (_03214_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _25064_ (_03215_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _25065_ (_03216_, _03215_, _03214_);
  and _25066_ (_03217_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _25067_ (_03218_, _01819_, _12194_);
  or _25068_ (_03219_, _03218_, _03217_);
  or _25069_ (_03220_, _03219_, _03216_);
  or _25070_ (_03221_, _01846_, p3_in[1]);
  or _25071_ (_03223_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _25072_ (_03224_, _03223_, _03221_);
  and _25073_ (_03225_, _03224_, _01830_);
  or _25074_ (_03226_, _01846_, p2_in[1]);
  or _25075_ (_03227_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _25076_ (_03228_, _03227_, _03226_);
  and _25077_ (_03229_, _03228_, _01853_);
  or _25078_ (_03230_, _03229_, _03225_);
  or _25079_ (_03231_, _01846_, p1_in[1]);
  or _25080_ (_03232_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _25081_ (_03233_, _03232_, _03231_);
  and _25082_ (_03234_, _03233_, _01865_);
  or _25083_ (_03235_, _01846_, p0_in[1]);
  or _25084_ (_03236_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _25085_ (_03237_, _03236_, _03235_);
  and _25086_ (_03238_, _03237_, _01859_);
  or _25087_ (_03239_, _03238_, _03234_);
  or _25088_ (_03240_, _03239_, _03230_);
  or _25089_ (_03241_, _03240_, _03220_);
  or _25090_ (_03242_, _03241_, _03213_);
  or _25091_ (_03243_, _03242_, _03210_);
  and _25092_ (_03244_, _03243_, _01893_);
  and _25093_ (_03245_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  or _25094_ (_03246_, _03245_, _03244_);
  or _25095_ (_03247_, _03246_, _01732_);
  nand _25096_ (_03248_, _01732_, _06512_);
  and _25097_ (_03249_, _03248_, _05110_);
  and _25098_ (_03766_, _03249_, _03247_);
  or _25099_ (_03250_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor _25100_ (_03251_, _01721_, rst);
  and _25101_ (_03769_, _03251_, _03250_);
  and _25102_ (_03252_, _11871_, _11960_);
  and _25103_ (_03253_, _01815_, _03252_);
  and _25104_ (_03254_, _03253_, _06617_);
  nor _25105_ (_03255_, _03254_, _12086_);
  and _25106_ (_03256_, _01748_, _06183_);
  or _25107_ (_03257_, _03256_, _12268_);
  and _25108_ (_03258_, _01737_, _12874_);
  and _25109_ (_03259_, _01762_, _12894_);
  and _25110_ (_03260_, _01724_, _08224_);
  or _25111_ (_03261_, _03260_, _03259_);
  or _25112_ (_03262_, _03261_, _03258_);
  or _25113_ (_03263_, _03262_, _03257_);
  and _25114_ (_03264_, _01748_, _06559_);
  or _25115_ (_03265_, _03264_, _12270_);
  and _25116_ (_03266_, _01737_, _06799_);
  and _25117_ (_03267_, _01762_, _06194_);
  and _25118_ (_03268_, _01724_, _06230_);
  or _25119_ (_03269_, _03268_, _03267_);
  or _25120_ (_03270_, _03269_, _03266_);
  or _25121_ (_03271_, _03270_, _03265_);
  nand _25122_ (_03272_, _03271_, _03263_);
  nor _25123_ (_03273_, _03272_, _03255_);
  or _25124_ (_03274_, _11873_, _11960_);
  or _25125_ (_03275_, _03274_, _01903_);
  or _25126_ (_03276_, _03154_, _12270_);
  or _25127_ (_03277_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _25128_ (_03278_, _03277_, _01737_);
  and _25129_ (_03279_, _03278_, _03276_);
  and _25130_ (_03280_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _25131_ (_03281_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _25132_ (_03282_, _03281_, _03280_);
  and _25133_ (_03283_, _03282_, _12270_);
  and _25134_ (_03284_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _25135_ (_03285_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _25136_ (_03286_, _03285_, _03284_);
  and _25137_ (_03287_, _03286_, _01762_);
  and _25138_ (_03288_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _25139_ (_03289_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _25140_ (_03290_, _03289_, _03288_);
  and _25141_ (_03291_, _03290_, _12268_);
  or _25142_ (_03292_, _03291_, _03287_);
  or _25143_ (_03293_, _03292_, _03283_);
  nor _25144_ (_03294_, _03293_, _03279_);
  nor _25145_ (_03295_, _03294_, _03275_);
  and _25146_ (_03296_, _01769_, _11871_);
  or _25147_ (_03297_, _01846_, p3_in[5]);
  or _25148_ (_03298_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _25149_ (_03299_, _03298_, _03297_);
  and _25150_ (_03300_, _03299_, _12270_);
  and _25151_ (_03301_, _03224_, _12268_);
  or _25152_ (_03302_, _03301_, _03300_);
  and _25153_ (_03303_, _03302_, _01748_);
  and _25154_ (_03304_, _01850_, _12270_);
  or _25155_ (_03305_, _01846_, p3_in[3]);
  or _25156_ (_03306_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _25157_ (_03307_, _03306_, _03305_);
  and _25158_ (_03308_, _03307_, _12268_);
  or _25159_ (_03310_, _03308_, _03304_);
  and _25160_ (_03311_, _03310_, _01762_);
  or _25161_ (_03312_, _01846_, p3_in[4]);
  or _25162_ (_03313_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _25163_ (_03314_, _03313_, _03312_);
  and _25164_ (_03315_, _03314_, _12270_);
  and _25165_ (_03317_, _03091_, _12268_);
  or _25166_ (_03318_, _03317_, _03315_);
  and _25167_ (_03319_, _03318_, _01737_);
  and _25168_ (_03320_, _02995_, _12270_);
  or _25169_ (_03321_, _01846_, p3_in[2]);
  or _25170_ (_03322_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _25171_ (_03323_, _03322_, _03321_);
  and _25172_ (_03324_, _03323_, _12268_);
  or _25173_ (_03325_, _03324_, _03320_);
  and _25174_ (_03326_, _03325_, _01724_);
  or _25175_ (_03327_, _03326_, _03319_);
  or _25176_ (_03328_, _03327_, _03311_);
  or _25177_ (_03329_, _03328_, _03303_);
  and _25178_ (_03330_, _03329_, _11958_);
  and _25179_ (_03331_, _01856_, _12270_);
  or _25180_ (_03332_, _01846_, p2_in[3]);
  or _25181_ (_03333_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _25182_ (_03334_, _03333_, _03332_);
  and _25183_ (_03335_, _03334_, _12268_);
  or _25184_ (_03336_, _03335_, _03331_);
  and _25185_ (_03337_, _03336_, _01762_);
  or _25186_ (_03338_, _01846_, p2_in[2]);
  or _25187_ (_03339_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _25188_ (_03340_, _03339_, _03338_);
  or _25189_ (_03341_, _03340_, _12270_);
  or _25190_ (_03342_, _02991_, _12268_);
  and _25191_ (_03343_, _03342_, _03341_);
  and _25192_ (_03344_, _03343_, _01724_);
  or _25193_ (_03345_, _01846_, p2_in[4]);
  or _25194_ (_03346_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _25195_ (_03347_, _03346_, _03345_);
  and _25196_ (_03348_, _03347_, _12270_);
  and _25197_ (_03349_, _03095_, _12268_);
  or _25198_ (_03350_, _03349_, _03348_);
  and _25199_ (_03351_, _03350_, _01737_);
  or _25200_ (_03352_, _03351_, _03344_);
  or _25201_ (_03353_, _01846_, p2_in[5]);
  or _25202_ (_03354_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _25203_ (_03355_, _03354_, _03353_);
  and _25204_ (_03356_, _03355_, _12270_);
  and _25205_ (_03357_, _03228_, _12268_);
  or _25206_ (_03358_, _03357_, _03356_);
  and _25207_ (_03359_, _03358_, _01748_);
  or _25208_ (_03360_, _03359_, _03352_);
  or _25209_ (_03361_, _03360_, _03337_);
  and _25210_ (_03362_, _03361_, _11960_);
  nor _25211_ (_03363_, _03362_, _03330_);
  nand _25212_ (_03364_, _03363_, _03296_);
  and _25213_ (_03365_, _01815_, _11871_);
  nand _25214_ (_03366_, _03252_, _01727_);
  nand _25215_ (_03367_, _03275_, _03366_);
  nor _25216_ (_03368_, _03367_, _03365_);
  nand _25217_ (_03369_, _01794_, _11871_);
  and _25218_ (_03370_, _11918_, _12071_);
  and _25219_ (_03371_, _11873_, _01725_);
  and _25220_ (_03372_, _03371_, _11960_);
  and _25221_ (_03373_, _03372_, _03370_);
  or _25222_ (_03374_, _01918_, _11871_);
  nand _25223_ (_03375_, _03374_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _25224_ (_03376_, _03375_, _03373_);
  and _25225_ (_03377_, _03376_, _03369_);
  and _25226_ (_03378_, _03377_, _03368_);
  or _25227_ (_03379_, _03378_, _03296_);
  and _25228_ (_03380_, _03379_, _03364_);
  and _25229_ (_03381_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _25230_ (_03382_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _25231_ (_03383_, _03382_, _03381_);
  and _25232_ (_03384_, _03383_, _01737_);
  and _25233_ (_03385_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _25234_ (_03386_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _25235_ (_03387_, _03386_, _03385_);
  and _25236_ (_03388_, _03387_, _01762_);
  or _25237_ (_03389_, _03388_, _03384_);
  and _25238_ (_03390_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _25239_ (_03391_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _25240_ (_03392_, _03391_, _03390_);
  and _25241_ (_03393_, _03392_, _01724_);
  and _25242_ (_03394_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _25243_ (_03395_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _25244_ (_03396_, _03395_, _03394_);
  and _25245_ (_03397_, _03396_, _01748_);
  or _25246_ (_03398_, _03397_, _03393_);
  or _25247_ (_03399_, _03398_, _03389_);
  and _25248_ (_03400_, _03399_, _01728_);
  and _25249_ (_03401_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _25250_ (_03402_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _25251_ (_03403_, _03402_, _03401_);
  and _25252_ (_03404_, _03403_, _01737_);
  and _25253_ (_03405_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _25254_ (_03406_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _25255_ (_03407_, _03406_, _03405_);
  and _25256_ (_03408_, _03407_, _01748_);
  or _25257_ (_03409_, _03408_, _03404_);
  and _25258_ (_03410_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _25259_ (_03411_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _25260_ (_03412_, _03411_, _03410_);
  and _25261_ (_03413_, _03412_, _01724_);
  and _25262_ (_03414_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _25263_ (_03415_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _25264_ (_03416_, _03415_, _03414_);
  and _25265_ (_03417_, _03416_, _01762_);
  or _25266_ (_03418_, _03417_, _03413_);
  or _25267_ (_03419_, _03418_, _03409_);
  and _25268_ (_03420_, _03419_, _01776_);
  or _25269_ (_03421_, _03420_, _03400_);
  and _25270_ (_03422_, _03421_, _11873_);
  and _25271_ (_03423_, _01737_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _25272_ (_03424_, _03423_, _12268_);
  and _25273_ (_03425_, _01762_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _25274_ (_03426_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _25275_ (_03427_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or _25276_ (_03428_, _03427_, _03426_);
  or _25277_ (_03429_, _03428_, _03425_);
  or _25278_ (_03430_, _03429_, _03424_);
  and _25279_ (_03431_, _03365_, _11958_);
  and _25280_ (_03432_, _01737_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _25281_ (_03433_, _03432_, _12270_);
  and _25282_ (_03434_, _01762_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _25283_ (_03435_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _25284_ (_03436_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _25285_ (_03437_, _03436_, _03435_);
  or _25286_ (_03438_, _03437_, _03434_);
  or _25287_ (_03439_, _03438_, _03433_);
  and _25288_ (_03440_, _03439_, _03431_);
  and _25289_ (_03441_, _03440_, _03430_);
  and _25290_ (_03442_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _25291_ (_03443_, _03442_, _12270_);
  and _25292_ (_03444_, _01737_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _25293_ (_03445_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _25294_ (_03446_, _01762_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _25295_ (_03447_, _03446_, _03445_);
  or _25296_ (_03448_, _03447_, _03444_);
  or _25297_ (_03449_, _03448_, _03443_);
  and _25298_ (_03450_, _01748_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _25299_ (_03451_, _03450_, _12268_);
  and _25300_ (_03452_, _01737_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _25301_ (_03453_, _01724_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _25302_ (_03454_, _01762_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _25303_ (_03455_, _03454_, _03453_);
  or _25304_ (_03456_, _03455_, _03452_);
  or _25305_ (_03457_, _03456_, _03451_);
  and _25306_ (_03458_, _03457_, _03253_);
  and _25307_ (_03459_, _03458_, _03449_);
  or _25308_ (_03460_, _03459_, _03441_);
  or _25309_ (_03461_, _03460_, _03422_);
  and _25310_ (_03462_, _03106_, _01737_);
  or _25311_ (_03463_, _03462_, _12270_);
  or _25312_ (_03464_, _01846_, p1_in[3]);
  or _25313_ (_03465_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _25314_ (_03466_, _03465_, _03464_);
  and _25315_ (_03467_, _03466_, _01762_);
  or _25316_ (_03468_, _01846_, p1_in[2]);
  or _25317_ (_03469_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _25318_ (_03470_, _03469_, _03468_);
  and _25319_ (_03471_, _03470_, _01724_);
  and _25320_ (_03472_, _03233_, _01748_);
  or _25321_ (_03473_, _03472_, _03471_);
  or _25322_ (_03474_, _03473_, _03467_);
  or _25323_ (_03475_, _03474_, _03463_);
  and _25324_ (_03476_, _03000_, _01724_);
  or _25325_ (_03477_, _03476_, _12268_);
  or _25326_ (_03478_, _01846_, p1_in[4]);
  or _25327_ (_03479_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _25328_ (_03480_, _03479_, _03478_);
  and _25329_ (_03481_, _03480_, _01737_);
  or _25330_ (_03482_, _01846_, p1_in[5]);
  or _25331_ (_03483_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _25332_ (_03484_, _03483_, _03482_);
  and _25333_ (_03485_, _03484_, _01748_);
  and _25334_ (_03486_, _01868_, _01762_);
  or _25335_ (_03487_, _03486_, _03485_);
  or _25336_ (_03488_, _03487_, _03481_);
  or _25337_ (_03489_, _03488_, _03477_);
  and _25338_ (_03490_, _03489_, _03475_);
  or _25339_ (_03491_, _03490_, _11873_);
  and _25340_ (_03492_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _25341_ (_03493_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _25342_ (_03494_, _03493_, _03492_);
  and _25343_ (_03495_, _03494_, _01724_);
  and _25344_ (_03496_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _25345_ (_03497_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _25346_ (_03498_, _03497_, _03496_);
  and _25347_ (_03499_, _03498_, _01737_);
  or _25348_ (_03500_, _03499_, _03495_);
  and _25349_ (_03501_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _25350_ (_03502_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _25351_ (_03503_, _03502_, _03501_);
  and _25352_ (_03504_, _03503_, _01762_);
  or _25353_ (_03505_, _03504_, _03500_);
  and _25354_ (_03506_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _25355_ (_03507_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _25356_ (_03508_, _03507_, _03506_);
  and _25357_ (_03509_, _03508_, _01748_);
  or _25358_ (_03510_, _03509_, _11871_);
  or _25359_ (_03511_, _03510_, _03505_);
  and _25360_ (_03512_, _03511_, _01794_);
  and _25361_ (_03513_, _03512_, _03491_);
  nand _25362_ (_03514_, _12338_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _25363_ (_03515_, _01770_, _11873_);
  and _25364_ (_03516_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _25365_ (_03517_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _25366_ (_03518_, _03517_, _03516_);
  and _25367_ (_03519_, _03518_, _01737_);
  and _25368_ (_03520_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _25369_ (_03521_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _25370_ (_03522_, _03521_, _03520_);
  and _25371_ (_03523_, _03522_, _01748_);
  or _25372_ (_03524_, _03523_, _03519_);
  and _25373_ (_03525_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _25374_ (_03526_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _25375_ (_03527_, _03526_, _03525_);
  and _25376_ (_03528_, _03527_, _01724_);
  and _25377_ (_03529_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _25378_ (_03530_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _25379_ (_03531_, _03530_, _03529_);
  and _25380_ (_03533_, _03531_, _01762_);
  or _25381_ (_03535_, _03533_, _03528_);
  or _25382_ (_03536_, _03535_, _03524_);
  and _25383_ (_03537_, _03536_, _03515_);
  and _25384_ (_03538_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _25385_ (_03539_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _25386_ (_03540_, _03539_, _03538_);
  and _25387_ (_03541_, _03540_, _01724_);
  and _25388_ (_03542_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _25389_ (_03543_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _25390_ (_03544_, _03543_, _03542_);
  and _25391_ (_03545_, _03544_, _01748_);
  or _25392_ (_03546_, _03545_, _03541_);
  and _25393_ (_03547_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _25394_ (_03548_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _25395_ (_03549_, _03548_, _03547_);
  and _25396_ (_03550_, _03549_, _01737_);
  and _25397_ (_03551_, _12270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _25398_ (_03552_, _12268_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _25399_ (_03553_, _03552_, _03551_);
  and _25400_ (_03554_, _03553_, _01762_);
  or _25401_ (_03555_, _03554_, _03550_);
  or _25402_ (_03556_, _03555_, _03546_);
  and _25403_ (_03557_, _03556_, _03373_);
  or _25404_ (_03558_, _01846_, p0_in[4]);
  or _25405_ (_03559_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _25406_ (_03560_, _03559_, _03558_);
  and _25407_ (_03561_, _03560_, _12270_);
  and _25408_ (_03562_, _03102_, _12268_);
  or _25409_ (_03563_, _03562_, _03561_);
  and _25410_ (_03564_, _03563_, _01737_);
  and _25411_ (_03565_, _01863_, _12270_);
  or _25412_ (_03566_, _01846_, p0_in[3]);
  or _25413_ (_03567_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _25414_ (_03568_, _03567_, _03566_);
  and _25415_ (_03569_, _03568_, _12268_);
  or _25416_ (_03570_, _03569_, _03565_);
  and _25417_ (_03572_, _03570_, _01762_);
  or _25418_ (_03573_, _03572_, _03564_);
  and _25419_ (_03574_, _03005_, _12270_);
  or _25420_ (_03575_, _01846_, p0_in[2]);
  or _25421_ (_03576_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _25422_ (_03577_, _03576_, _03575_);
  and _25423_ (_03578_, _03577_, _12268_);
  or _25424_ (_03579_, _03578_, _03574_);
  and _25425_ (_03580_, _03579_, _01724_);
  or _25426_ (_03581_, _01846_, p0_in[5]);
  or _25427_ (_03582_, _01848_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _25428_ (_03583_, _03582_, _03581_);
  and _25429_ (_03584_, _03583_, _12270_);
  and _25430_ (_03585_, _03237_, _12268_);
  or _25431_ (_03586_, _03585_, _03584_);
  and _25432_ (_03587_, _03586_, _01748_);
  or _25433_ (_03588_, _03587_, _03580_);
  nor _25434_ (_03589_, _03588_, _03573_);
  nor _25435_ (_03590_, _03589_, _03366_);
  or _25436_ (_03591_, _03590_, _03557_);
  nor _25437_ (_03592_, _03591_, _03537_);
  nand _25438_ (_03594_, _03592_, _03514_);
  or _25439_ (_03595_, _03594_, _03513_);
  or _25440_ (_03597_, _03595_, _03461_);
  or _25441_ (_03598_, _03597_, _03380_);
  or _25442_ (_03600_, _03598_, _03295_);
  or _25443_ (_03601_, _03514_, _05782_);
  and _25444_ (_03602_, _03601_, _03255_);
  and _25445_ (_03603_, _03602_, _03600_);
  or _25446_ (_03604_, _03603_, _03273_);
  and _25447_ (_03797_, _03604_, _05110_);
  and _25448_ (_03605_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _25449_ (_03606_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  or _25450_ (_03607_, _03606_, _03605_);
  and _25451_ (_03834_, _03607_, _05110_);
  or _25452_ (_03608_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand _25453_ (_03609_, _06205_, _12984_);
  and _25454_ (_03610_, _03609_, _05110_);
  and _25455_ (_03849_, _03610_, _03608_);
  and _25456_ (_03611_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _25457_ (_03612_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  or _25458_ (_03613_, _03612_, _03611_);
  and _25459_ (_03857_, _03613_, _05110_);
  nor _25460_ (_03614_, _01721_, _01720_);
  or _25461_ (_03615_, _03614_, _01722_);
  and _25462_ (_03616_, _03037_, _05110_);
  and _25463_ (_03866_, _03616_, _03615_);
  and _25464_ (_03617_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _25465_ (_03618_, pc_log_change, _01639_);
  or _25466_ (_03619_, _03618_, _03617_);
  and _25467_ (_03868_, _03619_, _05110_);
  nor _25468_ (_03877_, _03123_, rst);
  or _25469_ (_03620_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand _25470_ (_03621_, _06205_, _13092_);
  and _25471_ (_03622_, _03621_, _05110_);
  and _25472_ (_03895_, _03622_, _03620_);
  and _25473_ (_03623_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _25474_ (_03624_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  or _25475_ (_03625_, _03624_, _03623_);
  and _25476_ (_03899_, _03625_, _05110_);
  and _25477_ (_03626_, _01320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _25478_ (_03627_, _07034_, _06002_);
  or _25479_ (_03628_, _03627_, _03626_);
  and _25480_ (_03907_, _03628_, _05110_);
  and _25481_ (_03629_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _25482_ (_03630_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or _25483_ (_03631_, _03630_, _03629_);
  and _25484_ (_03910_, _03631_, _05110_);
  and _25485_ (_03632_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _25486_ (_03633_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or _25487_ (_03634_, _03633_, _03632_);
  and _25488_ (_03912_, _03634_, _05110_);
  or _25489_ (_03635_, _06205_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand _25490_ (_03636_, _06205_, _12904_);
  and _25491_ (_03637_, _03636_, _05110_);
  and _25492_ (_03914_, _03637_, _03635_);
  nand _25493_ (_03638_, _06798_, _06673_);
  or _25494_ (_03639_, _06673_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _25495_ (_03640_, _03639_, _03638_);
  and _25496_ (_03919_, _03640_, _05110_);
  nand _25497_ (_03641_, _00531_, _07028_);
  or _25498_ (_03642_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _25499_ (_03643_, _03642_, _05806_);
  and _25500_ (_03644_, _03643_, _03641_);
  and _25501_ (_03645_, _00529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _25502_ (_03646_, _00523_, _05867_);
  nand _25503_ (_03647_, _03646_, _05872_);
  or _25504_ (_03648_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _25505_ (_03649_, _03648_, _05794_);
  and _25506_ (_03650_, _03649_, _03647_);
  or _25507_ (_03651_, _03650_, _03645_);
  or _25508_ (_03652_, _03651_, _03644_);
  and _25509_ (_03929_, _03652_, _05110_);
  nor _25510_ (_03653_, _08056_, _05841_);
  and _25511_ (_03654_, _08117_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or _25512_ (_03655_, _03654_, _03653_);
  and _25513_ (_03972_, _03655_, _05110_);
  nor _25514_ (_03656_, _01320_, _05334_);
  and _25515_ (_03657_, _01320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or _25516_ (_03658_, _03657_, _03656_);
  and _25517_ (_03985_, _03658_, _05110_);
  and _25518_ (_03661_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _25519_ (_03662_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or _25520_ (_03664_, _03662_, _03661_);
  and _25521_ (_03665_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _25522_ (_03666_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _25523_ (_03667_, _03666_, _03665_);
  or _25524_ (_03668_, _03667_, _03664_);
  and _25525_ (_03669_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _25526_ (_03671_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or _25527_ (_03672_, _03671_, _03669_);
  and _25528_ (_03673_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _25529_ (_03674_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _25530_ (_03675_, _03674_, _03673_);
  or _25531_ (_03676_, _03675_, _03672_);
  or _25532_ (_03677_, _03676_, _03668_);
  and _25533_ (_03678_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _25534_ (_03679_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or _25535_ (_03680_, _03679_, _03678_);
  and _25536_ (_03681_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _25537_ (_03682_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _25538_ (_03683_, _03682_, _03681_);
  or _25539_ (_03685_, _03683_, _03680_);
  and _25540_ (_03687_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and _25541_ (_03688_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _25542_ (_03689_, _03688_, _03687_);
  and _25543_ (_03690_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _25544_ (_03691_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or _25545_ (_03692_, _03691_, _03690_);
  or _25546_ (_03693_, _03692_, _03689_);
  or _25547_ (_03694_, _03693_, _03685_);
  or _25548_ (_03695_, _03694_, _03677_);
  and _25549_ (_03696_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _25550_ (_03697_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _25551_ (_03698_, _03697_, _03696_);
  and _25552_ (_03699_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _25553_ (_03700_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _25554_ (_03701_, _03700_, _03699_);
  and _25555_ (_03702_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not _25556_ (_03703_, _11866_);
  and _25557_ (_03705_, _01819_, _03703_);
  or _25558_ (_03707_, _03705_, _03702_);
  or _25559_ (_03708_, _03707_, _03701_);
  and _25560_ (_03710_, _03334_, _01853_);
  and _25561_ (_03711_, _03307_, _01830_);
  or _25562_ (_03712_, _03711_, _03710_);
  and _25563_ (_03713_, _03466_, _01865_);
  and _25564_ (_03714_, _03568_, _01859_);
  or _25565_ (_03715_, _03714_, _03713_);
  or _25566_ (_03716_, _03715_, _03712_);
  or _25567_ (_03717_, _03716_, _03708_);
  or _25568_ (_03718_, _03717_, _03698_);
  or _25569_ (_03719_, _03718_, _03695_);
  and _25570_ (_03720_, _03719_, _01893_);
  and _25571_ (_03721_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  or _25572_ (_03722_, _03721_, _03720_);
  or _25573_ (_03723_, _03722_, _01732_);
  nand _25574_ (_03725_, _01732_, _06668_);
  and _25575_ (_03726_, _03725_, _05110_);
  and _25576_ (_03992_, _03726_, _03723_);
  or _25577_ (_03727_, _08750_, _02720_);
  or _25578_ (_03728_, _08752_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _25579_ (_03729_, _03728_, _05110_);
  and _25580_ (_03994_, _03729_, _03727_);
  and _25581_ (_03730_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _25582_ (_03731_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _25583_ (_03732_, _03731_, _03730_);
  and _25584_ (_03733_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _25585_ (_03734_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _25586_ (_03735_, _03734_, _03733_);
  or _25587_ (_03736_, _03735_, _03732_);
  and _25588_ (_03737_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _25589_ (_03738_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _25590_ (_03739_, _03738_, _03737_);
  and _25591_ (_03740_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _25592_ (_03741_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _25593_ (_03742_, _03741_, _03740_);
  or _25594_ (_03743_, _03742_, _03739_);
  or _25595_ (_03744_, _03743_, _03736_);
  and _25596_ (_03745_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _25597_ (_03746_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _25598_ (_03747_, _03746_, _03745_);
  and _25599_ (_03749_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _25600_ (_03750_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _25601_ (_03751_, _03750_, _03749_);
  or _25602_ (_03752_, _03751_, _03747_);
  and _25603_ (_03753_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and _25604_ (_03754_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _25605_ (_03756_, _03754_, _03753_);
  and _25606_ (_03757_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _25607_ (_03758_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or _25608_ (_03759_, _03758_, _03757_);
  or _25609_ (_03760_, _03759_, _03756_);
  or _25610_ (_03761_, _03760_, _03752_);
  or _25611_ (_03762_, _03761_, _03744_);
  and _25612_ (_03763_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and _25613_ (_03764_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _25614_ (_03765_, _03764_, _03763_);
  and _25615_ (_03767_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _25616_ (_03768_, _01819_, _12262_);
  or _25617_ (_03770_, _03768_, _03767_);
  and _25618_ (_03771_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _25619_ (_03772_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _25620_ (_03773_, _03772_, _03771_);
  or _25621_ (_03774_, _03773_, _03770_);
  and _25622_ (_03775_, _03340_, _01853_);
  and _25623_ (_03776_, _03323_, _01830_);
  or _25624_ (_03777_, _03776_, _03775_);
  and _25625_ (_03778_, _03577_, _01859_);
  and _25626_ (_03779_, _03470_, _01865_);
  or _25627_ (_03780_, _03779_, _03778_);
  or _25628_ (_03781_, _03780_, _03777_);
  or _25629_ (_03782_, _03781_, _03774_);
  or _25630_ (_03783_, _03782_, _03765_);
  or _25631_ (_03784_, _03783_, _03762_);
  and _25632_ (_03785_, _03784_, _01893_);
  and _25633_ (_03786_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  or _25634_ (_03787_, _03786_, _03785_);
  or _25635_ (_03788_, _03787_, _01732_);
  nand _25636_ (_03789_, _01732_, _07337_);
  and _25637_ (_03790_, _03789_, _05110_);
  and _25638_ (_03996_, _03790_, _03788_);
  and _25639_ (_03791_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _25640_ (_03792_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or _25641_ (_03793_, _03792_, _03791_);
  and _25642_ (_03999_, _03793_, _05110_);
  and _25643_ (_03794_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _25644_ (_03795_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  or _25645_ (_03796_, _03795_, _03794_);
  and _25646_ (_04001_, _03796_, _05110_);
  or _25647_ (_03798_, _01892_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _25648_ (_03799_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _25649_ (_03800_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _25650_ (_03801_, _03800_, _03799_);
  and _25651_ (_03802_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _25652_ (_03803_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _25653_ (_03804_, _03803_, _03802_);
  or _25654_ (_03805_, _03804_, _03801_);
  and _25655_ (_03806_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _25656_ (_03807_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _25657_ (_03808_, _03807_, _03806_);
  and _25658_ (_03809_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _25659_ (_03810_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _25660_ (_03811_, _03810_, _03809_);
  or _25661_ (_03812_, _03811_, _03808_);
  or _25662_ (_03813_, _03812_, _03805_);
  and _25663_ (_03814_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _25664_ (_03815_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _25665_ (_03816_, _03815_, _03814_);
  and _25666_ (_03817_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _25667_ (_03818_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _25668_ (_03819_, _03818_, _03817_);
  or _25669_ (_03820_, _03819_, _03816_);
  and _25670_ (_03821_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _25671_ (_03822_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _25672_ (_03823_, _03822_, _03821_);
  and _25673_ (_03824_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _25674_ (_03825_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _25675_ (_03826_, _03825_, _03824_);
  or _25676_ (_03827_, _03826_, _03823_);
  or _25677_ (_03828_, _03827_, _03820_);
  or _25678_ (_03829_, _03828_, _03813_);
  and _25679_ (_03830_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _25680_ (_03831_, _01819_, _11890_);
  or _25681_ (_03833_, _03831_, _03830_);
  and _25682_ (_03835_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _25683_ (_03836_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _25684_ (_03837_, _03836_, _03835_);
  or _25685_ (_03838_, _03837_, _03833_);
  and _25686_ (_03839_, _03299_, _01830_);
  and _25687_ (_03840_, _03355_, _01853_);
  or _25688_ (_03841_, _03840_, _03839_);
  and _25689_ (_03842_, _03484_, _01865_);
  and _25690_ (_03843_, _03583_, _01859_);
  or _25691_ (_03844_, _03843_, _03842_);
  or _25692_ (_03845_, _03844_, _03841_);
  or _25693_ (_03846_, _03845_, _03838_);
  and _25694_ (_03847_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _25695_ (_03848_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or _25696_ (_03850_, _03848_, _03847_);
  or _25697_ (_03851_, _03850_, _03846_);
  or _25698_ (_03852_, _03851_, _03829_);
  and _25699_ (_03853_, _03852_, _01887_);
  and _25700_ (_03854_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or _25701_ (_03855_, _03854_, _03853_);
  and _25702_ (_03856_, _03855_, _03798_);
  or _25703_ (_03858_, _03856_, _01732_);
  nand _25704_ (_03859_, _01732_, _06548_);
  and _25705_ (_03860_, _03859_, _05110_);
  and _25706_ (_04003_, _03860_, _03858_);
  and _25707_ (_03861_, _01739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _25708_ (_03862_, _01744_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _25709_ (_03863_, _03862_, _03861_);
  and _25710_ (_03864_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _25711_ (_03865_, _01750_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _25712_ (_03867_, _03865_, _03864_);
  or _25713_ (_03869_, _03867_, _03863_);
  and _25714_ (_03870_, _01760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _25715_ (_03871_, _01765_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _25716_ (_03872_, _03871_, _03870_);
  and _25717_ (_03873_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _25718_ (_03874_, _01777_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _25719_ (_03875_, _03874_, _03873_);
  or _25720_ (_03876_, _03875_, _03872_);
  or _25721_ (_03878_, _03876_, _03869_);
  and _25722_ (_03879_, _01783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _25723_ (_03880_, _01785_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or _25724_ (_03881_, _03880_, _03879_);
  and _25725_ (_03882_, _01790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _25726_ (_03883_, _01788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _25727_ (_03884_, _03883_, _03882_);
  or _25728_ (_03885_, _03884_, _03881_);
  and _25729_ (_03886_, _01796_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and _25730_ (_03887_, _01798_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _25731_ (_03888_, _03887_, _03886_);
  and _25732_ (_03889_, _01803_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _25733_ (_03890_, _01806_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or _25734_ (_03891_, _03890_, _03889_);
  or _25735_ (_03892_, _03891_, _03888_);
  or _25736_ (_03893_, _03892_, _03885_);
  or _25737_ (_03894_, _03893_, _03878_);
  and _25738_ (_03896_, _01877_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _25739_ (_03897_, _01874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _25740_ (_03898_, _03897_, _03896_);
  and _25741_ (_03900_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _25742_ (_03901_, _01819_, _11954_);
  or _25743_ (_03902_, _03901_, _03900_);
  and _25744_ (_03903_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _25745_ (_03904_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _25746_ (_03905_, _03904_, _03903_);
  or _25747_ (_03906_, _03905_, _03902_);
  and _25748_ (_03908_, _03347_, _01853_);
  and _25749_ (_03909_, _03314_, _01830_);
  or _25750_ (_03911_, _03909_, _03908_);
  and _25751_ (_03913_, _03560_, _01859_);
  and _25752_ (_03915_, _03480_, _01865_);
  or _25753_ (_03916_, _03915_, _03913_);
  or _25754_ (_03917_, _03916_, _03911_);
  or _25755_ (_03918_, _03917_, _03906_);
  or _25756_ (_03920_, _03918_, _03898_);
  or _25757_ (_03921_, _03920_, _03894_);
  and _25758_ (_03922_, _03921_, _01893_);
  and _25759_ (_03923_, _01948_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  or _25760_ (_03924_, _03923_, _03922_);
  or _25761_ (_03925_, _03924_, _01732_);
  nand _25762_ (_03926_, _01732_, _07235_);
  and _25763_ (_03927_, _03926_, _05110_);
  and _25764_ (_04065_, _03927_, _03925_);
  and _25765_ (_03928_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _25766_ (_03930_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or _25767_ (_03931_, _03930_, _03928_);
  and _25768_ (_04067_, _03931_, _05110_);
  and _25769_ (_03932_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _25770_ (_03933_, pc_log_change, _02462_);
  or _25771_ (_03934_, _03933_, _03932_);
  and _25772_ (_04070_, _03934_, _05110_);
  and _25773_ (_03935_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _25774_ (_03936_, pc_log_change, _02373_);
  or _25775_ (_03937_, _03936_, _03935_);
  and _25776_ (_04112_, _03937_, _05110_);
  and _25777_ (_03938_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _25778_ (_03939_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or _25779_ (_03940_, _03939_, _03938_);
  and _25780_ (_04114_, _03940_, _05110_);
  and _25781_ (_03941_, pc_log_change, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _25782_ (_03942_, pc_log_change, _02377_);
  or _25783_ (_03943_, _03942_, _03941_);
  and _25784_ (_04166_, _03943_, _05110_);
  not _25785_ (_03944_, cy_reg);
  and _25786_ (_03945_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _25787_ (_03946_, _03945_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or _25788_ (_03947_, _03946_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nand _25789_ (_03948_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _25790_ (_03949_, _03948_, _05482_);
  or _25791_ (_03951_, _03949_, _00664_);
  and _25792_ (_03952_, _03951_, _03947_);
  or _25793_ (_03953_, _03952_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _25794_ (_03954_, _03945_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _25795_ (_03955_, _03954_, _03949_);
  and _25796_ (_03956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _07627_);
  not _25797_ (_03957_, _03956_);
  and _25798_ (_03958_, _03957_, _03955_);
  nand _25799_ (_03959_, _03958_, _03953_);
  not _25800_ (_03960_, _03955_);
  or _25801_ (_03961_, _03952_, _07604_);
  nand _25802_ (_03962_, _03952_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nand _25803_ (_03963_, _03962_, _03961_);
  nand _25804_ (_03964_, _03963_, _03960_);
  nand _25805_ (_03965_, _03964_, _03959_);
  nor _25806_ (_03966_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nand _25807_ (_03967_, _03966_, _03965_);
  or _25808_ (_03968_, _03952_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _25809_ (_03969_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _02468_);
  or _25810_ (_03970_, _00664_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _25811_ (_03971_, _03970_, _03969_);
  and _25812_ (_03973_, _03971_, _03968_);
  nand _25813_ (_03974_, _03951_, _03947_);
  or _25814_ (_03975_, _03974_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _25815_ (_03976_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and _25816_ (_03977_, _03976_, _03945_);
  and _25817_ (_03978_, _03977_, _03975_);
  or _25818_ (_03979_, _03978_, _03973_);
  and _25819_ (_03980_, _03979_, _03955_);
  or _25820_ (_03981_, _03952_, _07666_);
  nand _25821_ (_03982_, _03952_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _25822_ (_03983_, _03982_, _03981_);
  and _25823_ (_03984_, _03983_, _03946_);
  not _25824_ (_03986_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _25825_ (_03987_, _03952_, _03986_);
  or _25826_ (_03988_, _03974_, _08206_);
  nand _25827_ (_03989_, _03988_, _03987_);
  not _25828_ (_03990_, _03969_);
  nor _25829_ (_03991_, _03990_, _03955_);
  and _25830_ (_03993_, _03991_, _03989_);
  or _25831_ (_03995_, _03993_, _03984_);
  nor _25832_ (_03997_, _03995_, _03980_);
  and _25833_ (_03998_, _02381_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _25834_ (_04000_, _03974_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _25835_ (_04002_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  not _25836_ (_04004_, _04002_);
  and _25837_ (_04005_, _04004_, _03955_);
  nand _25838_ (_04006_, _04005_, _04000_);
  or _25839_ (_04007_, _03952_, _07638_);
  nand _25840_ (_04008_, _03952_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nand _25841_ (_04009_, _04008_, _04007_);
  nand _25842_ (_04010_, _04009_, _03960_);
  nand _25843_ (_04011_, _04010_, _04006_);
  nand _25844_ (_04012_, _04011_, _03998_);
  and _25845_ (_04013_, _04012_, _03997_);
  and _25846_ (_04014_, _04013_, _03967_);
  and _25847_ (_04015_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _25848_ (_04016_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _25849_ (_04017_, _04016_, _04015_);
  and _25850_ (_04018_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _25851_ (_04019_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _25852_ (_04020_, _04019_, _04018_);
  and _25853_ (_04021_, _04020_, _04017_);
  and _25854_ (_04022_, _04021_, _03960_);
  and _25855_ (_04023_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _25856_ (_04024_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _25857_ (_04025_, _04024_, _04023_);
  and _25858_ (_04026_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _25859_ (_04027_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _25860_ (_04028_, _04027_, _04026_);
  and _25861_ (_04029_, _04028_, _04025_);
  and _25862_ (_04030_, _04029_, _03955_);
  or _25863_ (_04031_, _04030_, _03952_);
  nor _25864_ (_04032_, _04031_, _04022_);
  and _25865_ (_04033_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _25866_ (_04034_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _25867_ (_04035_, _04034_, _04033_);
  and _25868_ (_04036_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _25869_ (_04037_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor _25870_ (_04038_, _04037_, _04036_);
  and _25871_ (_04039_, _04038_, _04035_);
  nor _25872_ (_04040_, _04039_, _03955_);
  and _25873_ (_04041_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _25874_ (_04042_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _25875_ (_04043_, _04042_, _04041_);
  and _25876_ (_04044_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _25877_ (_04045_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _25878_ (_04046_, _04045_, _04044_);
  and _25879_ (_04047_, _04046_, _04043_);
  nor _25880_ (_04048_, _04047_, _03960_);
  or _25881_ (_04049_, _04048_, _04040_);
  and _25882_ (_04050_, _04049_, _03952_);
  nor _25883_ (_04051_, _04050_, _04032_);
  nor _25884_ (_04052_, _04051_, _04014_);
  and _25885_ (_04053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _25886_ (_04054_, _04053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _25887_ (_04055_, _04054_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and _25888_ (_04056_, _04055_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and _25889_ (_04057_, _04056_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and _25890_ (_04058_, _04057_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _25891_ (_04059_, _04058_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _25892_ (_04060_, _04059_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and _25893_ (_04061_, _04060_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _25894_ (_04062_, _04061_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _25895_ (_04063_, _04062_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _25896_ (_04064_, _04063_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _25897_ (_04066_, _04064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _25898_ (_04068_, _04064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _25899_ (_04069_, _04068_, _04066_);
  and _25900_ (_04071_, _04069_, _04052_);
  nor _25901_ (_04072_, _04063_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _25902_ (_04073_, _04072_, _04064_);
  and _25903_ (_04074_, _04073_, _04052_);
  nor _25904_ (_04075_, _04073_, _04052_);
  nor _25905_ (_04076_, _04075_, _04074_);
  not _25906_ (_04077_, _04076_);
  nor _25907_ (_04078_, _04061_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _25908_ (_04079_, _04078_, _04062_);
  and _25909_ (_04080_, _04079_, _04052_);
  nor _25910_ (_04081_, _04060_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _25911_ (_04082_, _04081_, _04061_);
  and _25912_ (_04083_, _04082_, _04052_);
  and _25913_ (_04084_, _04083_, _13096_);
  nor _25914_ (_04085_, _04084_, _04080_);
  nor _25915_ (_04086_, _04079_, _04052_);
  nor _25916_ (_04087_, _04086_, _04080_);
  not _25917_ (_04088_, _04087_);
  nor _25918_ (_04089_, _04082_, _04052_);
  nor _25919_ (_04090_, _04089_, _04083_);
  nor _25920_ (_04091_, _04059_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _25921_ (_04092_, _04091_, _04060_);
  and _25922_ (_04093_, _04092_, _04052_);
  nor _25923_ (_04094_, _04058_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _25924_ (_04095_, _04094_, _04059_);
  and _25925_ (_04096_, _04095_, _04052_);
  nor _25926_ (_04097_, _04096_, _04093_);
  nor _25927_ (_04098_, _04092_, _04052_);
  nor _25928_ (_04099_, _04098_, _04093_);
  not _25929_ (_04100_, _04099_);
  nor _25930_ (_04101_, _04057_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _25931_ (_04102_, _04101_, _04058_);
  and _25932_ (_04103_, _04102_, _04052_);
  nor _25933_ (_04104_, _04102_, _04052_);
  and _25934_ (_04105_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _25935_ (_04106_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _25936_ (_04107_, _04106_, _04105_);
  and _25937_ (_04108_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _25938_ (_04109_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _25939_ (_04110_, _04109_, _04108_);
  and _25940_ (_04111_, _04110_, _04107_);
  and _25941_ (_04113_, _04111_, _03960_);
  and _25942_ (_04115_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _25943_ (_04116_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _25944_ (_04117_, _04116_, _04115_);
  and _25945_ (_04118_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _25946_ (_04119_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _25947_ (_04120_, _04119_, _04118_);
  and _25948_ (_04121_, _04120_, _04117_);
  and _25949_ (_04122_, _04121_, _03955_);
  or _25950_ (_04123_, _04122_, _03952_);
  nor _25951_ (_04124_, _04123_, _04113_);
  and _25952_ (_04125_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _25953_ (_04126_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _25954_ (_04127_, _04126_, _04125_);
  and _25955_ (_04128_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _25956_ (_04129_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _25957_ (_04130_, _04129_, _04128_);
  and _25958_ (_04131_, _04130_, _04127_);
  and _25959_ (_04132_, _04131_, _03960_);
  and _25960_ (_04133_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _25961_ (_04134_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _25962_ (_04135_, _04134_, _04133_);
  and _25963_ (_04136_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _25964_ (_04137_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _25965_ (_04138_, _04137_, _04136_);
  and _25966_ (_04139_, _04138_, _04135_);
  and _25967_ (_04140_, _04139_, _03955_);
  or _25968_ (_04141_, _04140_, _03974_);
  nor _25969_ (_04142_, _04141_, _04132_);
  nor _25970_ (_04143_, _04142_, _04124_);
  nor _25971_ (_04144_, _04143_, _04014_);
  nor _25972_ (_04145_, _04056_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _25973_ (_04146_, _04145_, _04057_);
  and _25974_ (_04147_, _04146_, _04144_);
  nor _25975_ (_04148_, _04146_, _04144_);
  nor _25976_ (_04149_, _04148_, _04147_);
  and _25977_ (_04150_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _25978_ (_04151_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _25979_ (_04152_, _04151_, _04150_);
  and _25980_ (_04153_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _25981_ (_04154_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _25982_ (_04155_, _04154_, _04153_);
  and _25983_ (_04156_, _04155_, _04152_);
  and _25984_ (_04157_, _04156_, _03960_);
  and _25985_ (_04158_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _25986_ (_04159_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _25987_ (_04160_, _04159_, _04158_);
  and _25988_ (_04161_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _25989_ (_04162_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _25990_ (_04163_, _04162_, _04161_);
  and _25991_ (_04164_, _04163_, _04160_);
  and _25992_ (_04165_, _04164_, _03955_);
  or _25993_ (_04167_, _04165_, _03952_);
  nor _25994_ (_04168_, _04167_, _04157_);
  and _25995_ (_04169_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _25996_ (_04170_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _25997_ (_04171_, _04170_, _04169_);
  and _25998_ (_04172_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _25999_ (_04173_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _26000_ (_04174_, _04173_, _04172_);
  and _26001_ (_04175_, _04174_, _04171_);
  and _26002_ (_04176_, _04175_, _03960_);
  and _26003_ (_04177_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _26004_ (_04178_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _26005_ (_04179_, _04178_, _04177_);
  and _26006_ (_04180_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _26007_ (_04181_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _26008_ (_04182_, _04181_, _04180_);
  and _26009_ (_04183_, _04182_, _04179_);
  and _26010_ (_04184_, _04183_, _03955_);
  or _26011_ (_04186_, _04184_, _03974_);
  nor _26012_ (_04187_, _04186_, _04176_);
  nor _26013_ (_04188_, _04187_, _04168_);
  nor _26014_ (_04189_, _04188_, _04014_);
  nor _26015_ (_04190_, _04055_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _26016_ (_04191_, _04190_, _04056_);
  and _26017_ (_04192_, _04191_, _04189_);
  nor _26018_ (_04193_, _04191_, _04189_);
  nor _26019_ (_04194_, _04193_, _04192_);
  and _26020_ (_04195_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _26021_ (_04196_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _26022_ (_04197_, _04196_, _04195_);
  and _26023_ (_04198_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _26024_ (_04199_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _26025_ (_04200_, _04199_, _04198_);
  and _26026_ (_04201_, _04200_, _04197_);
  and _26027_ (_04202_, _04201_, _03960_);
  and _26028_ (_04203_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _26029_ (_04204_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _26030_ (_04205_, _04204_, _04203_);
  and _26031_ (_04206_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _26032_ (_04207_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _26033_ (_04208_, _04207_, _04206_);
  and _26034_ (_04209_, _04208_, _04205_);
  and _26035_ (_04210_, _04209_, _03955_);
  or _26036_ (_04211_, _04210_, _03952_);
  nor _26037_ (_04212_, _04211_, _04202_);
  and _26038_ (_04213_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _26039_ (_04214_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _26040_ (_04215_, _04214_, _04213_);
  and _26041_ (_04216_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _26042_ (_04217_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _26043_ (_04218_, _04217_, _04216_);
  and _26044_ (_04219_, _04218_, _04215_);
  and _26045_ (_04220_, _04219_, _03955_);
  and _26046_ (_04221_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _26047_ (_04222_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _26048_ (_04223_, _04222_, _04221_);
  and _26049_ (_04224_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _26050_ (_04225_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _26051_ (_04226_, _04225_, _04224_);
  and _26052_ (_04227_, _04226_, _04223_);
  and _26053_ (_04228_, _04227_, _03960_);
  nor _26054_ (_04229_, _04228_, _04220_);
  and _26055_ (_04230_, _04229_, _03952_);
  nor _26056_ (_04231_, _04230_, _04212_);
  nor _26057_ (_04232_, _04231_, _04014_);
  nor _26058_ (_04233_, _04054_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _26059_ (_04234_, _04233_, _04055_);
  and _26060_ (_04235_, _04234_, _04232_);
  and _26061_ (_04236_, _04235_, _04194_);
  nor _26062_ (_04237_, _04236_, _04192_);
  and _26063_ (_04238_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _26064_ (_04239_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _26065_ (_04240_, _04239_, _04238_);
  and _26066_ (_04241_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _26067_ (_04242_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _26068_ (_04243_, _04242_, _04241_);
  and _26069_ (_04244_, _04243_, _04240_);
  and _26070_ (_04245_, _04244_, _03960_);
  and _26071_ (_04246_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _26072_ (_04247_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _26073_ (_04248_, _04247_, _04246_);
  and _26074_ (_04249_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _26075_ (_04250_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _26076_ (_04251_, _04250_, _04249_);
  and _26077_ (_04252_, _04251_, _04248_);
  and _26078_ (_04253_, _04252_, _03955_);
  or _26079_ (_04254_, _04253_, _03952_);
  nor _26080_ (_04255_, _04254_, _04245_);
  and _26081_ (_04256_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _26082_ (_04257_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _26083_ (_04258_, _04257_, _04256_);
  and _26084_ (_04259_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _26085_ (_04260_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _26086_ (_04261_, _04260_, _04259_);
  and _26087_ (_04262_, _04261_, _04258_);
  nor _26088_ (_04263_, _04262_, _03955_);
  and _26089_ (_04264_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _26090_ (_04265_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _26091_ (_04266_, _04265_, _04264_);
  and _26092_ (_04267_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _26093_ (_04268_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _26094_ (_04269_, _04268_, _04267_);
  and _26095_ (_04270_, _04269_, _04266_);
  nor _26096_ (_04271_, _04270_, _03960_);
  or _26097_ (_04272_, _04271_, _04263_);
  and _26098_ (_04273_, _04272_, _03952_);
  nor _26099_ (_04274_, _04273_, _04255_);
  nor _26100_ (_04275_, _04274_, _04014_);
  nor _26101_ (_04276_, _04053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _26102_ (_04277_, _04276_, _04054_);
  nand _26103_ (_04278_, _04277_, _04275_);
  or _26104_ (_04279_, _04277_, _04275_);
  and _26105_ (_04280_, _04279_, _04278_);
  not _26106_ (_04281_, _04280_);
  and _26107_ (_04282_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _05482_);
  and _26108_ (_04283_, _02468_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _26109_ (_04284_, _04283_, _04282_);
  not _26110_ (_04285_, _04284_);
  and _26111_ (_04286_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _26112_ (_04287_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _26113_ (_04288_, _04287_, _04286_);
  and _26114_ (_04289_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _26115_ (_04290_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _26116_ (_04291_, _04290_, _04289_);
  and _26117_ (_04292_, _04291_, _04288_);
  and _26118_ (_04293_, _04292_, _03960_);
  and _26119_ (_04294_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _26120_ (_04295_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _26121_ (_04297_, _04295_, _04294_);
  and _26122_ (_04298_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _26123_ (_04299_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _26124_ (_04300_, _04299_, _04298_);
  and _26125_ (_04301_, _04300_, _04297_);
  and _26126_ (_04302_, _04301_, _03955_);
  or _26127_ (_04303_, _04302_, _03952_);
  nor _26128_ (_04304_, _04303_, _04293_);
  and _26129_ (_04305_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _26130_ (_04306_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _26131_ (_04307_, _04306_, _04305_);
  and _26132_ (_04308_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _26133_ (_04309_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _26134_ (_04310_, _04309_, _04308_);
  and _26135_ (_04311_, _04310_, _04307_);
  nor _26136_ (_04312_, _04311_, _03955_);
  and _26137_ (_04313_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _26138_ (_04314_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _26139_ (_04315_, _04314_, _04313_);
  and _26140_ (_04316_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _26141_ (_04317_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _26142_ (_04318_, _04317_, _04316_);
  and _26143_ (_04319_, _04318_, _04315_);
  nor _26144_ (_04320_, _04319_, _03960_);
  or _26145_ (_04321_, _04320_, _04312_);
  and _26146_ (_04322_, _04321_, _03952_);
  nor _26147_ (_04323_, _04322_, _04304_);
  nor _26148_ (_04324_, _04323_, _04014_);
  nand _26149_ (_04325_, _04324_, _04285_);
  not _26150_ (_04326_, _04014_);
  and _26151_ (_04327_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _26152_ (_04328_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _26153_ (_04329_, _04328_, _04327_);
  and _26154_ (_04330_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _26155_ (_04331_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _26156_ (_04332_, _04331_, _04330_);
  and _26157_ (_04333_, _04332_, _04329_);
  and _26158_ (_04334_, _04333_, _03955_);
  nand _26159_ (_04335_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nand _26160_ (_04336_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _26161_ (_04337_, _04336_, _04335_);
  and _26162_ (_04338_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _26163_ (_04339_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _26164_ (_04340_, _04339_, _04338_);
  and _26165_ (_04341_, _04340_, _04337_);
  nand _26166_ (_04342_, _04341_, _03960_);
  nand _26167_ (_04343_, _04342_, _03952_);
  or _26168_ (_04344_, _04343_, _04334_);
  and _26169_ (_04345_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _26170_ (_04346_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _26171_ (_04347_, _04346_, _04345_);
  and _26172_ (_04348_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _26173_ (_04349_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _26174_ (_04350_, _04349_, _04348_);
  and _26175_ (_04351_, _04350_, _04347_);
  and _26176_ (_04352_, _04351_, _03955_);
  nand _26177_ (_04353_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nand _26178_ (_04354_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _26179_ (_04355_, _04354_, _04353_);
  and _26180_ (_04356_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _26181_ (_04357_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _26182_ (_04358_, _04357_, _04356_);
  and _26183_ (_04359_, _04358_, _04355_);
  nand _26184_ (_04360_, _04359_, _03960_);
  nand _26185_ (_04361_, _04360_, _03974_);
  or _26186_ (_04362_, _04361_, _04352_);
  nand _26187_ (_04363_, _04362_, _04344_);
  and _26188_ (_04364_, _04363_, _04326_);
  nand _26189_ (_04365_, _04364_, _02468_);
  and _26190_ (_04366_, _03969_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _26191_ (_04367_, _03945_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _26192_ (_04368_, _04367_, _04366_);
  and _26193_ (_04369_, _03998_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _26194_ (_04370_, _03966_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor _26195_ (_04371_, _04370_, _04369_);
  and _26196_ (_04372_, _04371_, _04368_);
  and _26197_ (_04373_, _04372_, _03960_);
  and _26198_ (_04374_, _03998_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _26199_ (_04375_, _03966_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _26200_ (_04376_, _04375_, _04374_);
  and _26201_ (_04378_, _03969_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _26202_ (_04379_, _03945_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _26203_ (_04380_, _04379_, _04378_);
  and _26204_ (_04381_, _04380_, _04376_);
  and _26205_ (_04382_, _04381_, _03955_);
  or _26206_ (_04383_, _04382_, _03952_);
  nor _26207_ (_04384_, _04383_, _04373_);
  and _26208_ (_04385_, _03969_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _26209_ (_04386_, _03998_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor _26210_ (_04387_, _04386_, _04385_);
  and _26211_ (_04388_, _03966_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _26212_ (_04389_, _03945_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _26213_ (_04390_, _04389_, _04388_);
  and _26214_ (_04391_, _04390_, _04387_);
  and _26215_ (_04392_, _04391_, _03960_);
  and _26216_ (_04393_, _03969_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _26217_ (_04394_, _03945_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _26218_ (_04395_, _04394_, _04393_);
  and _26219_ (_04396_, _03998_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _26220_ (_04397_, _03966_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _26221_ (_04398_, _04397_, _04396_);
  and _26222_ (_04399_, _04398_, _04395_);
  and _26223_ (_04400_, _04399_, _03955_);
  or _26224_ (_04401_, _04400_, _03974_);
  nor _26225_ (_04402_, _04401_, _04392_);
  nor _26226_ (_04403_, _04402_, _04384_);
  nor _26227_ (_04404_, _04403_, _04014_);
  and _26228_ (_04405_, _04404_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _26229_ (_04406_, _04364_, _02468_);
  nand _26230_ (_04407_, _04406_, _04365_);
  not _26231_ (_04408_, _04407_);
  nand _26232_ (_04409_, _04408_, _04405_);
  and _26233_ (_04410_, _04409_, _04365_);
  or _26234_ (_04411_, _04324_, _04285_);
  and _26235_ (_04412_, _04411_, _04325_);
  not _26236_ (_04413_, _04412_);
  or _26237_ (_04414_, _04413_, _04410_);
  and _26238_ (_04415_, _04414_, _04325_);
  or _26239_ (_04416_, _04415_, _04281_);
  nand _26240_ (_04417_, _04416_, _04278_);
  nor _26241_ (_04418_, _04234_, _04232_);
  nor _26242_ (_04419_, _04418_, _04235_);
  and _26243_ (_04420_, _04419_, _04194_);
  nand _26244_ (_04421_, _04420_, _04417_);
  nand _26245_ (_04422_, _04421_, _04237_);
  and _26246_ (_04423_, _04422_, _04149_);
  nor _26247_ (_04424_, _04423_, _04147_);
  nor _26248_ (_04425_, _04424_, _04104_);
  or _26249_ (_04426_, _04425_, _04103_);
  nor _26250_ (_04427_, _04095_, _04052_);
  nor _26251_ (_04428_, _04427_, _04096_);
  nand _26252_ (_04429_, _04428_, _04426_);
  or _26253_ (_04430_, _04429_, _04100_);
  nand _26254_ (_04431_, _04430_, _04097_);
  nand _26255_ (_04432_, _04431_, _04090_);
  or _26256_ (_04433_, _04432_, _04088_);
  nand _26257_ (_04434_, _04433_, _04085_);
  nor _26258_ (_04435_, _04062_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _26259_ (_04436_, _04435_, _04063_);
  and _26260_ (_04437_, _04436_, _04052_);
  nor _26261_ (_04438_, _04436_, _04052_);
  nor _26262_ (_04439_, _04438_, _04437_);
  nand _26263_ (_04440_, _04439_, _04434_);
  or _26264_ (_04441_, _04440_, _04077_);
  and _26265_ (_04442_, _04437_, _02369_);
  nor _26266_ (_04443_, _04442_, _04074_);
  nand _26267_ (_04444_, _04443_, _04441_);
  nor _26268_ (_04445_, _04069_, _04052_);
  nor _26269_ (_04446_, _04445_, _04071_);
  and _26270_ (_04447_, _04446_, _04444_);
  nor _26271_ (_04448_, _04447_, _04071_);
  or _26272_ (_04449_, _04066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand _26273_ (_04450_, _04066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and _26274_ (_04451_, _04450_, _04449_);
  nor _26275_ (_04452_, _04451_, _04052_);
  and _26276_ (_04453_, _04451_, _04052_);
  nor _26277_ (_04454_, _04453_, _04452_);
  or _26278_ (_04455_, _04454_, _04448_);
  nand _26279_ (_04456_, _04454_, _04448_);
  and _26280_ (_04457_, _04456_, _04455_);
  and _26281_ (_04458_, _04457_, _03944_);
  nor _26282_ (_04459_, _04451_, _03944_);
  or _26283_ (_04460_, _04459_, _04458_);
  nor _26284_ (_04461_, _04460_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _26285_ (_04462_, _04460_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _26286_ (_04463_, _04439_, _04434_);
  nor _26287_ (_04464_, _04463_, _04437_);
  nand _26288_ (_04465_, _04464_, _04077_);
  or _26289_ (_04466_, _04464_, _04077_);
  nand _26290_ (_04467_, _04466_, _04465_);
  and _26291_ (_04468_, _04467_, _03944_);
  nor _26292_ (_04469_, _04073_, _03944_);
  nor _26293_ (_04470_, _04469_, _04468_);
  nor _26294_ (_04471_, _04470_, _02385_);
  and _26295_ (_04472_, _04470_, _02385_);
  nor _26296_ (_04473_, _04079_, _03944_);
  and _26297_ (_04474_, _04431_, _04090_);
  nor _26298_ (_04475_, _04474_, _04083_);
  nand _26299_ (_04476_, _04475_, _04088_);
  or _26300_ (_04477_, _04475_, _04088_);
  nand _26301_ (_04478_, _04477_, _04476_);
  and _26302_ (_04479_, _04478_, _03944_);
  nor _26303_ (_04480_, _04479_, _04473_);
  nor _26304_ (_04481_, _04480_, _12879_);
  and _26305_ (_04482_, _04480_, _12879_);
  and _26306_ (_04483_, _04092_, cy_reg);
  and _26307_ (_04484_, _04428_, _04426_);
  nor _26308_ (_04485_, _04484_, _04096_);
  nand _26309_ (_04486_, _04485_, _04099_);
  or _26310_ (_04487_, _04485_, _04099_);
  nand _26311_ (_04488_, _04487_, _04486_);
  and _26312_ (_04489_, _04488_, _03944_);
  nor _26313_ (_04490_, _04489_, _04483_);
  nor _26314_ (_04491_, _04490_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _26315_ (_04492_, _04490_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  or _26316_ (_04493_, _04428_, _04426_);
  nand _26317_ (_04494_, _04493_, _04429_);
  and _26318_ (_04495_, _04494_, _03944_);
  nor _26319_ (_04496_, _04095_, _03944_);
  nor _26320_ (_04497_, _04496_, _04495_);
  nor _26321_ (_04498_, _04497_, _02462_);
  and _26322_ (_04499_, _04497_, _02462_);
  nor _26323_ (_04500_, _04102_, _03944_);
  nor _26324_ (_04501_, _04103_, _04104_);
  nand _26325_ (_04502_, _04501_, _04424_);
  or _26326_ (_04503_, _04501_, _04424_);
  and _26327_ (_04504_, _04503_, _03944_);
  and _26328_ (_04505_, _04504_, _04502_);
  or _26329_ (_04506_, _04505_, _04500_);
  nor _26330_ (_04507_, _04506_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _26331_ (_04508_, _04422_, _04149_);
  or _26332_ (_04509_, _04508_, _04423_);
  and _26333_ (_04510_, _04509_, _03944_);
  nor _26334_ (_04511_, _04146_, _03944_);
  or _26335_ (_04512_, _04511_, _04510_);
  nor _26336_ (_04513_, _04512_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not _26337_ (_04514_, _04235_);
  nand _26338_ (_04515_, _04419_, _04417_);
  nand _26339_ (_04516_, _04515_, _04514_);
  nand _26340_ (_04517_, _04516_, _04194_);
  or _26341_ (_04518_, _04516_, _04194_);
  nand _26342_ (_04519_, _04518_, _04517_);
  and _26343_ (_04520_, _04519_, _03944_);
  nor _26344_ (_04521_, _04191_, _03944_);
  or _26345_ (_04522_, _04521_, _04520_);
  nor _26346_ (_04523_, _04522_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _26347_ (_04524_, _04234_, cy_reg);
  or _26348_ (_04525_, _04419_, _04417_);
  and _26349_ (_04526_, _04525_, _04515_);
  and _26350_ (_04527_, _04526_, _03944_);
  or _26351_ (_04528_, _04527_, _04524_);
  and _26352_ (_04529_, _04528_, _02377_);
  and _26353_ (_04530_, _04277_, cy_reg);
  nand _26354_ (_04531_, _04415_, _04281_);
  and _26355_ (_04532_, _04531_, _04416_);
  and _26356_ (_04533_, _04532_, _03944_);
  nor _26357_ (_04534_, _04533_, _04530_);
  nor _26358_ (_04535_, _04534_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _26359_ (_04536_, _04284_, _03944_);
  nand _26360_ (_04537_, _04413_, _04410_);
  and _26361_ (_04538_, _04537_, _04414_);
  and _26362_ (_04539_, _04538_, _03944_);
  nor _26363_ (_04540_, _04539_, _04536_);
  nor _26364_ (_04541_, _04540_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26365_ (_04542_, _04404_, _03944_);
  nor _26366_ (_04543_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _26367_ (_04544_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _26368_ (_04545_, _04544_, _04543_);
  nand _26369_ (_04546_, _04545_, _04542_);
  or _26370_ (_04547_, _04545_, _04542_);
  and _26371_ (_04548_, _04547_, _04546_);
  or _26372_ (_04549_, _04548_, _04541_);
  or _26373_ (_04550_, _04549_, _04535_);
  or _26374_ (_04551_, _04550_, _04529_);
  or _26375_ (_04552_, _04551_, _04523_);
  or _26376_ (_04553_, _04552_, _04513_);
  and _26377_ (_04554_, _04506_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _26378_ (_04555_, _04512_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _26379_ (_04556_, _04522_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor _26380_ (_04557_, _04528_, _02377_);
  and _26381_ (_04558_, _04534_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _26382_ (_04559_, _04540_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26383_ (_04560_, cy_reg, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _26384_ (_04561_, _04408_, _04405_);
  nand _26385_ (_04562_, _04561_, _04409_);
  and _26386_ (_04563_, _04562_, _03944_);
  or _26387_ (_04564_, _04563_, _04560_);
  nor _26388_ (_04565_, _04564_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _26389_ (_04566_, _04564_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _26390_ (_04567_, _04566_, _04565_);
  or _26391_ (_04568_, _04567_, _04559_);
  or _26392_ (_04569_, _04568_, _04558_);
  or _26393_ (_04570_, _04569_, _04557_);
  or _26394_ (_04571_, _04570_, _04556_);
  or _26395_ (_04572_, _04571_, _04555_);
  or _26396_ (_04573_, _04572_, _04554_);
  or _26397_ (_04574_, _04573_, _04553_);
  or _26398_ (_04575_, _04574_, _04507_);
  or _26399_ (_04576_, _04575_, _04499_);
  or _26400_ (_04577_, _04576_, _04498_);
  or _26401_ (_04578_, _04577_, _04492_);
  or _26402_ (_04579_, _04578_, _04491_);
  and _26403_ (_04580_, _04082_, cy_reg);
  or _26404_ (_04581_, _04431_, _04090_);
  and _26405_ (_04582_, _04581_, _04432_);
  and _26406_ (_04583_, _04582_, _03944_);
  or _26407_ (_04584_, _04583_, _04580_);
  nor _26408_ (_04585_, _04584_, _02509_);
  and _26409_ (_04586_, _04584_, _02509_);
  or _26410_ (_04587_, _04586_, _04585_);
  or _26411_ (_04588_, _04587_, _04579_);
  or _26412_ (_04589_, _04588_, _04482_);
  or _26413_ (_04590_, _04589_, _04481_);
  and _26414_ (_04591_, _04436_, cy_reg);
  or _26415_ (_04592_, _04439_, _04434_);
  and _26416_ (_04593_, _04592_, _04440_);
  and _26417_ (_04594_, _04593_, _03944_);
  or _26418_ (_04595_, _04594_, _04591_);
  nor _26419_ (_04596_, _04595_, _01639_);
  and _26420_ (_04597_, _04595_, _01639_);
  or _26421_ (_04598_, _04597_, _04596_);
  or _26422_ (_04599_, _04598_, _04590_);
  or _26423_ (_04600_, _04599_, _04472_);
  or _26424_ (_04601_, _04600_, _04471_);
  and _26425_ (_04602_, _04069_, cy_reg);
  nor _26426_ (_04603_, _04446_, _04444_);
  nor _26427_ (_04604_, _04603_, _04447_);
  and _26428_ (_04605_, _04604_, _03944_);
  or _26429_ (_04606_, _04605_, _04602_);
  nor _26430_ (_04607_, _04606_, _00990_);
  and _26431_ (_04608_, _04606_, _00990_);
  or _26432_ (_04609_, _04608_, _04607_);
  or _26433_ (_04610_, _04609_, _04601_);
  or _26434_ (_04611_, _04610_, _04462_);
  or _26435_ (_04612_, _04611_, _04461_);
  nor _26436_ (_04613_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _26437_ (_04614_, _04613_, _02396_);
  nor _26438_ (_04615_, _04614_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _26439_ (_04616_, _04614_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _26440_ (_04617_, _04616_, _04615_);
  or _26441_ (_04618_, _01339_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _26442_ (_04619_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and _26443_ (_04620_, _04619_, _04618_);
  or _26444_ (_04621_, _04620_, _04617_);
  and _26445_ (_04622_, _04613_, _02396_);
  nor _26446_ (_04623_, _04622_, _04614_);
  or _26447_ (_04624_, _01339_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _26448_ (_04625_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _26449_ (_04626_, _04625_, _04624_);
  and _26450_ (_04627_, _04626_, _04617_);
  nor _26451_ (_04628_, _04627_, _04623_);
  and _26452_ (_04629_, _04628_, _04621_);
  and _26453_ (_04630_, _04617_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _26454_ (_04631_, _02477_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _26455_ (_04632_, _04631_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _26456_ (_04633_, _04632_, _04630_);
  and _26457_ (_04634_, _04617_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _26458_ (_04635_, _02477_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _26459_ (_04636_, _04635_, _01339_);
  or _26460_ (_04637_, _04636_, _04634_);
  and _26461_ (_04638_, _04637_, _04623_);
  and _26462_ (_04639_, _04638_, _04633_);
  or _26463_ (_04640_, _04639_, _04629_);
  and _26464_ (_04641_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _26465_ (_04642_, _04641_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _26466_ (_04643_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _26467_ (_04644_, _04643_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _26468_ (_04645_, _04644_, _04642_);
  not _26469_ (_04646_, _04645_);
  nor _26470_ (_04647_, _04642_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _26471_ (_04648_, _04642_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _26472_ (_04649_, _04648_, _04647_);
  or _26473_ (_04650_, _04649_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _26474_ (_04651_, _02477_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _26475_ (_04652_, _04651_, _04650_);
  or _26476_ (_04653_, _04652_, _04646_);
  nand _26477_ (_04654_, _04649_, _08206_);
  or _26478_ (_04655_, _04649_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _26479_ (_04656_, _04655_, _04654_);
  or _26480_ (_04657_, _04656_, _04645_);
  and _26481_ (_04658_, _04657_, _04653_);
  or _26482_ (_04659_, _04658_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _26483_ (_04660_, _04649_, _07666_);
  and _26484_ (_04661_, _04649_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _26485_ (_04662_, _04661_, _04660_);
  and _26486_ (_04663_, _04662_, _04646_);
  or _26487_ (_04664_, _04649_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _26488_ (_04665_, _02477_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _26489_ (_04666_, _04665_, _04645_);
  and _26490_ (_04667_, _04666_, _04664_);
  or _26491_ (_04668_, _04667_, _01339_);
  or _26492_ (_04669_, _04668_, _04663_);
  or _26493_ (_04670_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  or _26494_ (_04671_, _02477_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _26495_ (_04672_, _04671_, _04670_);
  or _26496_ (_04673_, _04672_, _02396_);
  or _26497_ (_04674_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  or _26498_ (_04675_, _02477_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _26499_ (_04676_, _04675_, _04674_);
  or _26500_ (_04677_, _04676_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26501_ (_04678_, _04677_, _04673_);
  and _26502_ (_04679_, _04678_, _04643_);
  and _26503_ (_04680_, _01339_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _26504_ (_04681_, _02477_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or _26505_ (_04682_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and _26506_ (_04683_, _04682_, _04681_);
  or _26507_ (_04684_, _04683_, _02396_);
  or _26508_ (_04685_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or _26509_ (_04686_, _02477_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _26510_ (_04687_, _04686_, _04685_);
  or _26511_ (_04688_, _04687_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26512_ (_04689_, _04688_, _04684_);
  and _26513_ (_04690_, _04689_, _04680_);
  or _26514_ (_04691_, _04690_, _04679_);
  and _26515_ (_04692_, _04678_, _01339_);
  and _26516_ (_04693_, _02396_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _26517_ (_04694_, _04693_, _04683_);
  or _26518_ (_04695_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  or _26519_ (_04696_, _02477_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _26520_ (_04697_, _04696_, _04641_);
  and _26521_ (_04698_, _04697_, _04695_);
  or _26522_ (_04699_, _04698_, _04694_);
  or _26523_ (_04700_, _04699_, _04692_);
  and _26524_ (_04701_, _04700_, _04691_);
  and _26525_ (_04702_, _04701_, _04669_);
  and _26526_ (_04703_, _04702_, _04659_);
  and _26527_ (_04704_, _04703_, _04640_);
  and _26528_ (_04705_, _04617_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand _26529_ (_04706_, _02477_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand _26530_ (_04707_, _04706_, _04623_);
  or _26531_ (_04708_, _04707_, _04705_);
  and _26532_ (_04709_, _04708_, _01339_);
  nor _26533_ (_04710_, _04617_, _07638_);
  and _26534_ (_04711_, _04617_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _26535_ (_04712_, _04711_, _04710_);
  or _26536_ (_04713_, _04712_, _04623_);
  and _26537_ (_04714_, _04713_, _04709_);
  or _26538_ (_04715_, _04714_, _04699_);
  and _26539_ (_04716_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _26540_ (_04717_, _02477_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _26541_ (_04718_, _04717_, _04716_);
  and _26542_ (_04719_, _04718_, _02396_);
  and _26543_ (_04720_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or _26544_ (_04721_, _04720_, _04631_);
  and _26545_ (_04722_, _04721_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _26546_ (_04723_, _04722_, _04719_);
  and _26547_ (_04724_, _04723_, _01339_);
  or _26548_ (_04725_, _04649_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _26549_ (_04726_, _04681_, _04645_);
  and _26550_ (_04727_, _04726_, _04725_);
  not _26551_ (_04728_, _04649_);
  or _26552_ (_04729_, _04728_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _26553_ (_04730_, _04649_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _26554_ (_04731_, _04730_, _04646_);
  and _26555_ (_04732_, _04731_, _04729_);
  or _26556_ (_04733_, _04732_, _04727_);
  and _26557_ (_04734_, _04733_, _04724_);
  or _26558_ (_04735_, _04649_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _26559_ (_04736_, _04671_, _04645_);
  and _26560_ (_04737_, _04736_, _04735_);
  or _26561_ (_04738_, _04728_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _26562_ (_04739_, _04649_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _26563_ (_04740_, _04739_, _04646_);
  and _26564_ (_04741_, _04740_, _04738_);
  or _26565_ (_04742_, _04741_, _04737_);
  and _26566_ (_04743_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  or _26567_ (_04744_, _04635_, _02396_);
  or _26568_ (_04745_, _04744_, _04743_);
  or _26569_ (_04746_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or _26570_ (_04747_, _02477_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _26571_ (_04748_, _04747_, _04746_);
  or _26572_ (_04749_, _04748_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _26573_ (_04750_, _04749_, _04745_);
  and _26574_ (_04751_, _04750_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _26575_ (_04752_, _04721_, _04693_);
  or _26576_ (_04753_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or _26577_ (_04754_, _02477_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _26578_ (_04755_, _04754_, _04641_);
  and _26579_ (_04756_, _04755_, _04753_);
  or _26580_ (_04757_, _04756_, _04752_);
  and _26581_ (_04758_, _04757_, _04751_);
  and _26582_ (_04759_, _04758_, _04742_);
  or _26583_ (_04760_, _04759_, _04734_);
  or _26584_ (_04761_, _04757_, _04750_);
  and _26585_ (_04762_, _04761_, _02943_);
  and _26586_ (_04763_, _04762_, _04760_);
  and _26587_ (_04764_, _04763_, _04715_);
  or _26588_ (_04765_, _04764_, _04704_);
  not _26589_ (_04766_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _26590_ (_04767_, _03966_, _05482_);
  nor _26591_ (_04768_, _04767_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _26592_ (_04769_, _04767_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _26593_ (_04770_, _04769_, _04768_);
  nand _26594_ (_04771_, _04770_, _04766_);
  nor _26595_ (_04772_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _26596_ (_04773_, _04772_, _02381_);
  nor _26597_ (_04774_, _04773_, _04767_);
  or _26598_ (_04775_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and _26599_ (_04776_, _04775_, _04774_);
  and _26600_ (_04777_, _04776_, _04771_);
  not _26601_ (_04778_, _04774_);
  and _26602_ (_04779_, _04770_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _26603_ (_04780_, _04770_, _03986_);
  or _26604_ (_04781_, _04780_, _04779_);
  and _26605_ (_04782_, _04781_, _04778_);
  or _26606_ (_04783_, _04782_, _04777_);
  and _26607_ (_04784_, _04783_, _03945_);
  nand _26608_ (_04785_, _04770_, _07627_);
  or _26609_ (_04786_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and _26610_ (_04787_, _04786_, _04774_);
  and _26611_ (_04788_, _04787_, _04785_);
  and _26612_ (_04789_, _04770_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _26613_ (_04790_, _04770_, _07604_);
  or _26614_ (_04791_, _04790_, _04789_);
  and _26615_ (_04792_, _04791_, _04778_);
  or _26616_ (_04793_, _04792_, _04788_);
  and _26617_ (_04794_, _04793_, _03998_);
  or _26618_ (_04795_, _04794_, _04784_);
  nand _26619_ (_04796_, _04770_, _07647_);
  and _26620_ (_04797_, _04774_, _04004_);
  and _26621_ (_04798_, _04797_, _04796_);
  and _26622_ (_04799_, _04770_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _26623_ (_04800_, _04770_, _07638_);
  or _26624_ (_04801_, _04800_, _04799_);
  and _26625_ (_04802_, _04801_, _04778_);
  or _26626_ (_04803_, _04802_, _04798_);
  and _26627_ (_04804_, _04803_, _03966_);
  nand _26628_ (_04805_, _04770_, _07675_);
  and _26629_ (_04806_, _04774_, _03976_);
  and _26630_ (_04807_, _04806_, _04805_);
  and _26631_ (_04808_, _04770_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _26632_ (_04809_, _04770_, _07666_);
  or _26633_ (_04810_, _04809_, _04808_);
  and _26634_ (_04811_, _04810_, _04778_);
  or _26635_ (_04812_, _04811_, _04807_);
  and _26636_ (_04813_, _04812_, _03969_);
  or _26637_ (_04814_, _04813_, _04804_);
  or _26638_ (_04815_, _04814_, _04795_);
  or _26639_ (_04816_, \oc8051_symbolic_cxrom1.regarray[5] [1], \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand _26640_ (_04817_, _04816_, _03969_);
  or _26641_ (_04818_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand _26642_ (_04819_, _04818_, _03998_);
  and _26643_ (_04820_, _04819_, _04817_);
  or _26644_ (_04821_, _03948_, _09288_);
  nand _26645_ (_04822_, _03969_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _26646_ (_04823_, _04822_, _04821_);
  and _26647_ (_04824_, _04823_, _04820_);
  nand _26648_ (_04825_, _03998_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  or _26649_ (_04826_, _03948_, _07721_);
  and _26650_ (_04827_, _04826_, _04825_);
  nor _26651_ (_04828_, \oc8051_symbolic_cxrom1.regarray[7] [1], \oc8051_symbolic_cxrom1.regarray[7] [0]);
  or _26652_ (_04829_, _04828_, _03948_);
  nand _26653_ (_04830_, _03966_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _26654_ (_04831_, _04830_, _04829_);
  and _26655_ (_04832_, _04831_, _04827_);
  and _26656_ (_04833_, _04832_, _04824_);
  nand _26657_ (_04834_, _03966_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _26658_ (_04835_, \oc8051_symbolic_cxrom1.regarray[7] [3], \oc8051_symbolic_cxrom1.regarray[7] [2]);
  or _26659_ (_04836_, _04835_, _03948_);
  and _26660_ (_04837_, _04836_, _04834_);
  or _26661_ (_04838_, \oc8051_symbolic_cxrom1.regarray[5] [3], \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand _26662_ (_04839_, _04838_, _03969_);
  or _26663_ (_04840_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand _26664_ (_04841_, _04840_, _03998_);
  and _26665_ (_04842_, _04841_, _04839_);
  and _26666_ (_04843_, _04842_, _04837_);
  or _26667_ (_04844_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand _26668_ (_04845_, _04844_, _03966_);
  or _26669_ (_04846_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nand _26670_ (_04847_, _04846_, _03966_);
  and _26671_ (_04848_, _04847_, _04845_);
  nand _26672_ (_04849_, _03998_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nand _26673_ (_04850_, _03969_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _26674_ (_04851_, _04850_, _04849_);
  and _26675_ (_04852_, _04851_, _04848_);
  and _26676_ (_04853_, _04852_, _04843_);
  and _26677_ (_04854_, _03998_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _26678_ (_04855_, _03969_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  or _26679_ (_04856_, _04855_, _04854_);
  and _26680_ (_04857_, _03945_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _26681_ (_04858_, _03966_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  or _26682_ (_04859_, _04858_, _04857_);
  or _26683_ (_04860_, _04859_, _04856_);
  and _26684_ (_04861_, _03969_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _26685_ (_04862_, _03966_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  or _26686_ (_04863_, _04862_, _04861_);
  and _26687_ (_04864_, _03945_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _26688_ (_04865_, _03998_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  or _26689_ (_04866_, _04865_, _04864_);
  or _26690_ (_04867_, _04866_, _04863_);
  and _26691_ (_04868_, _04867_, _04860_);
  and _26692_ (_04869_, _04868_, _04853_);
  and _26693_ (_04870_, _04869_, _04833_);
  or _26694_ (_04871_, _04870_, _05482_);
  or _26695_ (_04872_, _03948_, _07716_);
  nand _26696_ (_04873_, _03966_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _26697_ (_04874_, _04873_, _04872_);
  nor _26698_ (_04875_, \oc8051_symbolic_cxrom1.regarray[3] [1], \oc8051_symbolic_cxrom1.regarray[3] [0]);
  or _26699_ (_04876_, _04875_, _03948_);
  or _26700_ (_04877_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand _26701_ (_04878_, _04877_, _03966_);
  and _26702_ (_04879_, _04878_, _04876_);
  and _26703_ (_04880_, _04879_, _04874_);
  nand _26704_ (_04881_, _03998_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  or _26705_ (_04882_, _03948_, _08830_);
  and _26706_ (_04883_, _04882_, _04881_);
  or _26707_ (_04884_, \oc8051_symbolic_cxrom1.regarray[1] [1], \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nand _26708_ (_04885_, _04884_, _03969_);
  or _26709_ (_04886_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nand _26710_ (_04887_, _04886_, _03998_);
  and _26711_ (_04888_, _04887_, _04885_);
  and _26712_ (_04889_, _04888_, _04883_);
  and _26713_ (_04890_, _04889_, _04880_);
  nand _26714_ (_04891_, _03969_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _26715_ (_04892_, \oc8051_symbolic_cxrom1.regarray[3] [3], \oc8051_symbolic_cxrom1.regarray[3] [2]);
  or _26716_ (_04893_, _04892_, _03948_);
  and _26717_ (_04894_, _04893_, _04891_);
  or _26718_ (_04895_, \oc8051_symbolic_cxrom1.regarray[1] [3], \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand _26719_ (_04896_, _04895_, _03969_);
  or _26720_ (_04897_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nand _26721_ (_04898_, _04897_, _03998_);
  and _26722_ (_04899_, _04898_, _04896_);
  and _26723_ (_04900_, _04899_, _04894_);
  nand _26724_ (_04901_, _03969_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  or _26725_ (_04902_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nand _26726_ (_04903_, _04902_, _03966_);
  and _26727_ (_04904_, _04903_, _04901_);
  nand _26728_ (_04905_, _03998_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _26729_ (_04906_, _03966_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _26730_ (_04907_, _04906_, _04905_);
  and _26731_ (_04908_, _04907_, _04904_);
  and _26732_ (_04909_, _04908_, _04900_);
  and _26733_ (_04910_, _03998_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _26734_ (_04911_, _03969_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  or _26735_ (_04912_, _04911_, _04910_);
  and _26736_ (_04913_, _03945_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _26737_ (_04914_, _03966_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  or _26738_ (_04915_, _04914_, _04913_);
  or _26739_ (_04916_, _04915_, _04912_);
  and _26740_ (_04917_, _03966_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _26741_ (_04918_, _03969_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  or _26742_ (_04919_, _04918_, _04917_);
  and _26743_ (_04920_, _03998_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _26744_ (_04921_, _03945_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  or _26745_ (_04922_, _04921_, _04920_);
  or _26746_ (_04923_, _04922_, _04919_);
  and _26747_ (_04924_, _04923_, _04916_);
  and _26748_ (_04925_, _04924_, _04909_);
  and _26749_ (_04926_, _04925_, _04890_);
  or _26750_ (_04927_, _04926_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _26751_ (_04928_, _04927_, _04871_);
  or _26752_ (_04929_, _04928_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _26753_ (_04930_, _03998_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _26754_ (_04931_, _03969_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  or _26755_ (_04932_, _04931_, _04930_);
  and _26756_ (_04933_, _03945_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _26757_ (_04934_, _03966_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  or _26758_ (_04935_, _04934_, _04933_);
  or _26759_ (_04936_, _04935_, _04932_);
  and _26760_ (_04937_, _03969_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _26761_ (_04938_, _03966_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  or _26762_ (_04939_, _04938_, _04937_);
  and _26763_ (_04940_, _03945_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _26764_ (_04941_, _03998_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  or _26765_ (_04942_, _04941_, _04940_);
  or _26766_ (_04943_, _04942_, _04939_);
  nand _26767_ (_04944_, _03998_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  or _26768_ (_04945_, _03948_, _09716_);
  and _26769_ (_04946_, _04945_, _04944_);
  nand _26770_ (_04947_, _03966_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _26771_ (_04948_, _04947_, _04946_);
  and _26772_ (_04949_, _04948_, _04943_);
  and _26773_ (_04950_, _04949_, _04936_);
  nor _26774_ (_04951_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor _26775_ (_04952_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nand _26776_ (_04953_, _04952_, _04951_);
  nand _26777_ (_04954_, _04953_, _03998_);
  not _26778_ (_04955_, _03966_);
  nor _26779_ (_04956_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _26780_ (_04957_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _26781_ (_04958_, _04957_, _04956_);
  or _26782_ (_04959_, _04958_, _04955_);
  nor _26783_ (_04960_, \oc8051_symbolic_cxrom1.regarray[9] [1], \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _26784_ (_04961_, \oc8051_symbolic_cxrom1.regarray[9] [3], \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand _26785_ (_04962_, _04961_, _04960_);
  nand _26786_ (_04963_, _04962_, _03969_);
  and _26787_ (_04964_, _04963_, _04959_);
  and _26788_ (_04965_, _04964_, _04954_);
  nand _26789_ (_04966_, _03998_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _26790_ (_04967_, _03969_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _26791_ (_04968_, _04967_, _04966_);
  or _26792_ (_04969_, _03948_, _07691_);
  nand _26793_ (_04970_, _03969_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _26794_ (_04971_, _04970_, _04969_);
  and _26795_ (_04972_, _04971_, _04968_);
  nor _26796_ (_04973_, \oc8051_symbolic_cxrom1.regarray[11] [3], \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _26797_ (_04974_, \oc8051_symbolic_cxrom1.regarray[11] [1], \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _26798_ (_04975_, _04974_, _04973_);
  or _26799_ (_04976_, _04975_, _03948_);
  nand _26800_ (_04977_, _03966_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _26801_ (_04978_, _04977_, _05482_);
  and _26802_ (_04979_, _04978_, _04976_);
  and _26803_ (_04980_, _04979_, _04972_);
  and _26804_ (_04981_, _04980_, _04965_);
  and _26805_ (_04982_, _04981_, _04950_);
  and _26806_ (_04983_, _03998_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _26807_ (_04984_, _03969_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  or _26808_ (_04985_, _04984_, _04983_);
  and _26809_ (_04986_, _03945_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _26810_ (_04987_, _03966_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  or _26811_ (_04988_, _04987_, _04986_);
  or _26812_ (_04989_, _04988_, _04985_);
  and _26813_ (_04990_, _03969_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _26814_ (_04991_, _03966_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  or _26815_ (_04992_, _04991_, _04990_);
  and _26816_ (_04993_, _03945_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _26817_ (_04994_, _03998_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  or _26818_ (_04995_, _04994_, _04993_);
  or _26819_ (_04996_, _04995_, _04992_);
  nand _26820_ (_04997_, _03966_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _26821_ (_04998_, _03998_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _26822_ (_04999_, _03969_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _26823_ (_05000_, _04999_, _04998_);
  and _26824_ (_05001_, _05000_, _04997_);
  and _26825_ (_05002_, _05001_, _04996_);
  and _26826_ (_05003_, _05002_, _04989_);
  nor _26827_ (_05004_, \oc8051_symbolic_cxrom1.regarray[13] [1], \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _26828_ (_05005_, \oc8051_symbolic_cxrom1.regarray[13] [3], \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand _26829_ (_05006_, _05005_, _05004_);
  nand _26830_ (_05007_, _05006_, _03969_);
  nor _26831_ (_05008_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _26832_ (_05009_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _26833_ (_05010_, _05009_, _05008_);
  or _26834_ (_05011_, _05010_, _04955_);
  nor _26835_ (_05012_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor _26836_ (_05013_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand _26837_ (_05014_, _05013_, _05012_);
  nand _26838_ (_05015_, _05014_, _03998_);
  and _26839_ (_05016_, _05015_, _05011_);
  and _26840_ (_05017_, _05016_, _05007_);
  nand _26841_ (_05018_, _03998_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  or _26842_ (_05019_, _03948_, _10131_);
  and _26843_ (_05020_, _05019_, _05018_);
  or _26844_ (_05021_, _03948_, _07684_);
  nand _26845_ (_05022_, _03966_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _26846_ (_05023_, _05022_, _05021_);
  and _26847_ (_05024_, _05023_, _05020_);
  nor _26848_ (_05025_, \oc8051_symbolic_cxrom1.regarray[15] [3], \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _26849_ (_05026_, \oc8051_symbolic_cxrom1.regarray[15] [1], \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _26850_ (_05027_, _05026_, _05025_);
  or _26851_ (_05028_, _05027_, _03948_);
  nand _26852_ (_05029_, _03969_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _26853_ (_05030_, _05029_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _26854_ (_05031_, _05030_, _05028_);
  and _26855_ (_05032_, _05031_, _05024_);
  and _26856_ (_05033_, _05032_, _05017_);
  and _26857_ (_05034_, _05033_, _05003_);
  or _26858_ (_05035_, _05034_, _00664_);
  or _26859_ (_05036_, _05035_, _04982_);
  and _26860_ (_05037_, _04775_, _03970_);
  or _26861_ (_05038_, _05037_, _05482_);
  or _26862_ (_05039_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or _26863_ (_05040_, _00664_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _26864_ (_05041_, _05040_, _05039_);
  or _26865_ (_05042_, _05041_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _26866_ (_05043_, _05042_, _05038_);
  and _26867_ (_05044_, _05043_, _02468_);
  or _26868_ (_05045_, _00664_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _26869_ (_05046_, _05045_, _03976_);
  and _26870_ (_05047_, _05046_, _04282_);
  or _26871_ (_05048_, _00664_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _26872_ (_05049_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _26873_ (_05050_, _05049_, _04053_);
  and _26874_ (_05051_, _05050_, _05048_);
  or _26875_ (_05052_, _05051_, _05047_);
  or _26876_ (_05053_, _05052_, _05044_);
  and _26877_ (_05054_, _05053_, _02381_);
  or _26878_ (_05055_, _00664_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _26879_ (_05056_, _04002_, _05482_);
  and _26880_ (_05057_, _05056_, _05055_);
  or _26881_ (_05058_, _00664_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _26882_ (_05059_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and _26883_ (_05060_, _05059_, _05482_);
  and _26884_ (_05061_, _05060_, _05058_);
  or _26885_ (_05062_, _05061_, _05057_);
  and _26886_ (_05063_, _05062_, _03969_);
  or _26887_ (_05064_, _00664_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _26888_ (_05065_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _26889_ (_05066_, _05065_, _05064_);
  and _26890_ (_05067_, _05066_, _03946_);
  and _26891_ (_05068_, _03945_, _05482_);
  and _26892_ (_05069_, _04786_, _03957_);
  and _26893_ (_05070_, _05069_, _05068_);
  or _26894_ (_05071_, _05070_, _05067_);
  or _26895_ (_05072_, _05071_, _05063_);
  and _26896_ (_05073_, _05062_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _26897_ (_05074_, _05069_, _04283_);
  or _26898_ (_05075_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or _26899_ (_05076_, _00664_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _26900_ (_05077_, _05076_, _05075_);
  and _26901_ (_05078_, _05077_, _04772_);
  or _26902_ (_05079_, _05078_, _02381_);
  or _26903_ (_05080_, _05079_, _05074_);
  or _26904_ (_05081_, _05080_, _05073_);
  and _26905_ (_05082_, _05081_, _05072_);
  or _26906_ (_05083_, _05082_, _05054_);
  and _26907_ (_05084_, _05043_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _26908_ (_05085_, _05046_, _04283_);
  and _26909_ (_05086_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _26910_ (_05087_, _00664_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _26911_ (_05088_, _05087_, _05086_);
  and _26912_ (_05089_, _05088_, _04772_);
  or _26913_ (_05090_, _05089_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _26914_ (_05091_, _05090_, _05085_);
  or _26915_ (_05092_, _05091_, _05084_);
  nor _26916_ (_05093_, _02505_, first_instr);
  and _26917_ (_05094_, _05093_, _05092_);
  and _26918_ (_05095_, _05094_, _05083_);
  and _26919_ (_05096_, _05095_, _05036_);
  and _26920_ (_05097_, _05096_, _04929_);
  and _26921_ (_05098_, _05097_, _04326_);
  and _26922_ (_05099_, _05098_, _04815_);
  and _26923_ (_05100_, _05099_, _04765_);
  and _26924_ (property_invalid_jnc, _05100_, _04612_);
  and _26925_ (_05101_, _06205_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _26926_ (_05102_, _12543_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  or _26927_ (_05103_, _05102_, _05101_);
  and _26928_ (_04185_, _05103_, _05110_);
  or _26929_ (_05104_, pc_log_change_r, _03944_);
  nand _26930_ (_05105_, pc_log_change_r, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand _26931_ (_00000_, _05105_, _05104_);
  and _26932_ (_05106_, _02505_, first_instr);
  or _26933_ (_00001_, _05106_, rst);
  dff _26934_ (cy_reg, _00000_, clk);
  dff _26935_ (pc_log_change_r, pc_log_change, clk);
  dff _26936_ (first_instr, _00001_, clk);
  dff _26937_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _08906_, clk);
  dff _26938_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _08909_, clk);
  dff _26939_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _08913_, clk);
  dff _26940_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _08916_, clk);
  dff _26941_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _08920_, clk);
  dff _26942_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _08923_, clk);
  dff _26943_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _08926_, clk);
  dff _26944_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _06039_, clk);
  dff _26945_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _08823_, clk);
  dff _26946_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _08826_, clk);
  dff _26947_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _08829_, clk);
  dff _26948_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _08832_, clk);
  dff _26949_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _08835_, clk);
  dff _26950_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _08839_, clk);
  dff _26951_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _08843_, clk);
  dff _26952_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _08846_, clk);
  dff _26953_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _13437_, clk);
  dff _26954_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _13438_, clk);
  dff _26955_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _13439_, clk);
  dff _26956_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _08744_, clk);
  dff _26957_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _13440_, clk);
  dff _26958_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _13441_, clk);
  dff _26959_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _13442_, clk);
  dff _26960_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _13443_, clk);
  dff _26961_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _08636_, clk);
  dff _26962_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _08640_, clk);
  dff _26963_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _08645_, clk);
  dff _26964_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _08650_, clk);
  dff _26965_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _13433_, clk);
  dff _26966_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _13434_, clk);
  dff _26967_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _13435_, clk);
  dff _26968_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _13436_, clk);
  dff _26969_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _08550_, clk);
  dff _26970_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _08552_, clk);
  dff _26971_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _08556_, clk);
  dff _26972_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _08559_, clk);
  dff _26973_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _08562_, clk);
  dff _26974_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _08566_, clk);
  dff _26975_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _08568_, clk);
  dff _26976_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _08571_, clk);
  dff _26977_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _08465_, clk);
  dff _26978_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _08468_, clk);
  dff _26979_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _08472_, clk);
  dff _26980_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _08475_, clk);
  dff _26981_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _08477_, clk);
  dff _26982_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _08479_, clk);
  dff _26983_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _08482_, clk);
  dff _26984_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _08485_, clk);
  dff _26985_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _08374_, clk);
  dff _26986_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _08377_, clk);
  dff _26987_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _08382_, clk);
  dff _26988_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _08386_, clk);
  dff _26989_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _08389_, clk);
  dff _26990_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _08392_, clk);
  dff _26991_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _08396_, clk);
  dff _26992_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _08399_, clk);
  dff _26993_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _13449_, clk);
  dff _26994_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _08271_, clk);
  dff _26995_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _08275_, clk);
  dff _26996_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _08279_, clk);
  dff _26997_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _08284_, clk);
  dff _26998_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _08289_, clk);
  dff _26999_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _08295_, clk);
  dff _27000_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _08299_, clk);
  dff _27001_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _08171_, clk);
  dff _27002_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _08175_, clk);
  dff _27003_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _13444_, clk);
  dff _27004_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _13445_, clk);
  dff _27005_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _13446_, clk);
  dff _27006_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _13447_, clk);
  dff _27007_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _13448_, clk);
  dff _27008_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _08185_, clk);
  dff _27009_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _08077_, clk);
  dff _27010_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _08080_, clk);
  dff _27011_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _08084_, clk);
  dff _27012_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _08089_, clk);
  dff _27013_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _08091_, clk);
  dff _27014_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _08094_, clk);
  dff _27015_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _08098_, clk);
  dff _27016_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _08103_, clk);
  dff _27017_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _07991_, clk);
  dff _27018_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _07994_, clk);
  dff _27019_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _07997_, clk);
  dff _27020_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _08000_, clk);
  dff _27021_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _08003_, clk);
  dff _27022_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _08006_, clk);
  dff _27023_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _08009_, clk);
  dff _27024_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _08012_, clk);
  dff _27025_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _07573_, clk);
  dff _27026_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _07577_, clk);
  dff _27027_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _07581_, clk);
  dff _27028_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _07584_, clk);
  dff _27029_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _07587_, clk);
  dff _27030_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _07590_, clk);
  dff _27031_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _07593_, clk);
  dff _27032_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _07597_, clk);
  dff _27033_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _07468_, clk);
  dff _27034_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _07472_, clk);
  dff _27035_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _07476_, clk);
  dff _27036_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _07481_, clk);
  dff _27037_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _07484_, clk);
  dff _27038_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _07488_, clk);
  dff _27039_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _07491_, clk);
  dff _27040_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _07495_, clk);
  dff _27041_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _07792_, clk);
  dff _27042_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _07795_, clk);
  dff _27043_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _07798_, clk);
  dff _27044_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _07803_, clk);
  dff _27045_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _07807_, clk);
  dff _27046_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _07812_, clk);
  dff _27047_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _07817_, clk);
  dff _27048_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _07822_, clk);
  dff _27049_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _07686_, clk);
  dff _27050_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _07689_, clk);
  dff _27051_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _07692_, clk);
  dff _27052_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _07697_, clk);
  dff _27053_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _07700_, clk);
  dff _27054_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _07703_, clk);
  dff _27055_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _07708_, clk);
  dff _27056_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _07713_, clk);
  dff _27057_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _07911_, clk);
  dff _27058_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _07915_, clk);
  dff _27059_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _07919_, clk);
  dff _27060_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _07922_, clk);
  dff _27061_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _07924_, clk);
  dff _27062_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _07928_, clk);
  dff _27063_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _07932_, clk);
  dff _27064_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _07934_, clk);
  dff _27065_ (\oc8051_symbolic_cxrom1.regvalid [0], _06060_, clk);
  dff _27066_ (\oc8051_symbolic_cxrom1.regvalid [1], _06090_, clk);
  dff _27067_ (\oc8051_symbolic_cxrom1.regvalid [2], _06133_, clk);
  dff _27068_ (\oc8051_symbolic_cxrom1.regvalid [3], _06181_, clk);
  dff _27069_ (\oc8051_symbolic_cxrom1.regvalid [4], _06236_, clk);
  dff _27070_ (\oc8051_symbolic_cxrom1.regvalid [5], _06299_, clk);
  dff _27071_ (\oc8051_symbolic_cxrom1.regvalid [6], _06361_, clk);
  dff _27072_ (\oc8051_symbolic_cxrom1.regvalid [7], _06441_, clk);
  dff _27073_ (\oc8051_symbolic_cxrom1.regvalid [8], _06527_, clk);
  dff _27074_ (\oc8051_symbolic_cxrom1.regvalid [9], _06614_, clk);
  dff _27075_ (\oc8051_symbolic_cxrom1.regvalid [10], _06715_, clk);
  dff _27076_ (\oc8051_symbolic_cxrom1.regvalid [11], _06806_, clk);
  dff _27077_ (\oc8051_symbolic_cxrom1.regvalid [12], _06900_, clk);
  dff _27078_ (\oc8051_symbolic_cxrom1.regvalid [13], _06995_, clk);
  dff _27079_ (\oc8051_symbolic_cxrom1.regvalid [14], _07112_, clk);
  dff _27080_ (\oc8051_symbolic_cxrom1.regvalid [15], _06013_, clk);
  dff _27081_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _05695_, clk);
  dff _27082_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _05698_, clk);
  dff _27083_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _05701_, clk);
  dff _27084_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _05704_, clk);
  dff _27085_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _05706_, clk);
  dff _27086_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _05709_, clk);
  dff _27087_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _05712_, clk);
  dff _27088_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _05565_, clk);
  dff _27089_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _10979_, clk);
  dff _27090_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _05721_, clk);
  dff _27091_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _05724_, clk);
  dff _27092_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _05727_, clk);
  dff _27093_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _05730_, clk);
  dff _27094_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _05733_, clk);
  dff _27095_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _12746_, clk);
  dff _27096_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _05745_, clk);
  dff _27097_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _05748_, clk);
  dff _27098_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _05750_, clk);
  dff _27099_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _12081_, clk);
  dff _27100_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _05757_, clk);
  dff _27101_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _05569_, clk);
  dff _27102_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _11725_, clk);
  dff _27103_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _12506_, clk);
  dff _27104_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _11704_, clk);
  dff _27105_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _12511_, clk);
  dff _27106_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _05342_, clk);
  dff _27107_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _11694_, clk);
  dff _27108_ (\oc8051_top_1.oc8051_decoder1.state [0], _05315_, clk);
  dff _27109_ (\oc8051_top_1.oc8051_decoder1.state [1], _11718_, clk);
  dff _27110_ (\oc8051_top_1.oc8051_decoder1.op [0], _05525_, clk);
  dff _27111_ (\oc8051_top_1.oc8051_decoder1.op [1], _09737_, clk);
  dff _27112_ (\oc8051_top_1.oc8051_decoder1.op [2], _09877_, clk);
  dff _27113_ (\oc8051_top_1.oc8051_decoder1.op [3], _09900_, clk);
  dff _27114_ (\oc8051_top_1.oc8051_decoder1.op [4], _09902_, clk);
  dff _27115_ (\oc8051_top_1.oc8051_decoder1.op [5], _09897_, clk);
  dff _27116_ (\oc8051_top_1.oc8051_decoder1.op [6], _09905_, clk);
  dff _27117_ (\oc8051_top_1.oc8051_decoder1.op [7], _02086_, clk);
  dff _27118_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _11679_, clk);
  dff _27119_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _02048_, clk);
  dff _27120_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _01001_, clk);
  dff _27121_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _02391_, clk);
  dff _27122_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _05179_, clk);
  dff _27123_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _02587_, clk);
  dff _27124_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _02607_, clk);
  dff _27125_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _05205_, clk);
  dff _27126_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _02812_, clk);
  dff _27127_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _02814_, clk);
  dff _27128_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _05208_, clk);
  dff _27129_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _02848_, clk);
  dff _27130_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _05331_, clk);
  dff _27131_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _02875_, clk);
  dff _27132_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _02881_, clk);
  dff _27133_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _02894_, clk);
  dff _27134_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _05477_, clk);
  dff _27135_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _02940_, clk);
  dff _27136_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _05430_, clk);
  dff _27137_ (\oc8051_top_1.oc8051_decoder1.wr , _05513_, clk);
  dff _27138_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _03919_, clk);
  dff _27139_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _02218_, clk);
  dff _27140_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _11913_, clk);
  dff _27141_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _03950_, clk);
  dff _27142_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _05107_, clk);
  dff _27143_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _04296_, clk);
  dff _27144_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _02925_, clk);
  dff _27145_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _02917_, clk);
  dff _27146_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _02738_, clk);
  dff _27147_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _02207_, clk);
  dff _27148_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _07166_, clk);
  dff _27149_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _02222_, clk);
  dff _27150_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _04377_, clk);
  dff _27151_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _01746_, clk);
  dff _27152_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _01905_, clk);
  dff _27153_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _02906_, clk);
  dff _27154_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _03907_, clk);
  dff _27155_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _03222_, clk);
  dff _27156_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _05108_, clk);
  dff _27157_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _02954_, clk);
  dff _27158_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _03985_, clk);
  dff _27159_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _02578_, clk);
  dff _27160_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _03057_, clk);
  dff _27161_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _01604_, clk);
  dff _27162_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _03033_, clk);
  dff _27163_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _06408_, clk);
  dff _27164_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _06372_, clk);
  dff _27165_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _06192_, clk);
  dff _27166_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _06684_, clk);
  dff _27167_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _02543_, clk);
  dff _27168_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _03972_, clk);
  dff _27169_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _02970_, clk);
  dff _27170_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _03316_, clk);
  dff _27171_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _08933_, clk);
  dff _27172_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _10862_, clk);
  dff _27173_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _00018_, clk);
  dff _27174_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _00921_, clk);
  dff _27175_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _05289_, clk);
  dff _27176_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _02820_, clk);
  dff _27177_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _02963_, clk);
  dff _27178_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _13169_, clk);
  dff _27179_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _07653_, clk);
  dff _27180_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _00648_, clk);
  dff _27181_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _07648_, clk);
  dff _27182_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _03755_, clk);
  dff _27183_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _03534_, clk);
  dff _27184_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _03663_, clk);
  dff _27185_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _01577_, clk);
  dff _27186_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _05173_, clk);
  dff _27187_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _07639_, clk);
  dff _27188_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _03709_, clk);
  dff _27189_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _07665_, clk);
  dff _27190_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _05161_, clk);
  dff _27191_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _10144_, clk);
  dff _27192_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _01540_, clk);
  dff _27193_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _07102_, clk);
  dff _27194_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _05428_, clk);
  dff _27195_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _12941_, clk);
  dff _27196_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _13173_, clk);
  dff _27197_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _12945_, clk);
  dff _27198_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _12614_, clk);
  dff _27199_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _12886_, clk);
  dff _27200_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _06855_, clk);
  dff _27201_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _11392_, clk);
  dff _27202_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _01561_, clk);
  dff _27203_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _01531_, clk);
  dff _27204_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _00824_, clk);
  dff _27205_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _00590_, clk);
  dff _27206_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _10714_, clk);
  dff _27207_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _03670_, clk);
  dff _27208_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _01646_, clk);
  dff _27209_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _02780_, clk);
  dff _27210_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _02837_, clk);
  dff _27211_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _04166_, clk);
  dff _27212_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _01869_, clk);
  dff _27213_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _02776_, clk);
  dff _27214_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _04112_, clk);
  dff _27215_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _04070_, clk);
  dff _27216_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _02774_, clk);
  dff _27217_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _02863_, clk);
  dff _27218_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _11004_, clk);
  dff _27219_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _03868_, clk);
  dff _27220_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _02771_, clk);
  dff _27221_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _00915_, clk);
  dff _27222_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _13027_, clk);
  dff _27223_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _02763_, clk);
  dff _27224_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _02828_, clk);
  dff _27225_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _06919_, clk);
  dff _27226_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _00377_, clk);
  dff _27227_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _02762_, clk);
  dff _27228_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _06782_, clk);
  dff _27229_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _10427_, clk);
  dff _27230_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _02759_, clk);
  dff _27231_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _02825_, clk);
  dff _27232_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _02850_, clk);
  dff _27233_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _02861_, clk);
  dff _27234_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _11702_, clk);
  dff _27235_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _02010_, clk);
  dff _27236_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _02755_, clk);
  dff _27237_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _03660_, clk);
  dff _27238_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _13022_, clk);
  dff _27239_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _10724_, clk);
  dff _27240_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _10883_, clk);
  dff _27241_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _11198_, clk);
  dff _27242_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _02834_, clk);
  dff _27243_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _02255_, clk);
  dff _27244_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _13108_, clk);
  dff _27245_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _11991_, clk);
  dff _27246_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _08747_, clk);
  dff _27247_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _08380_, clk);
  dff _27248_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _12124_, clk);
  dff _27249_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _03849_, clk);
  dff _27250_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _03001_, clk);
  dff _27251_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _11980_, clk);
  dff _27252_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _10720_, clk);
  dff _27253_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _03895_, clk);
  dff _27254_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _03914_, clk);
  dff _27255_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _03912_, clk);
  dff _27256_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _03910_, clk);
  dff _27257_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _03899_, clk);
  dff _27258_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _12019_, clk);
  dff _27259_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _04185_, clk);
  dff _27260_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _04114_, clk);
  dff _27261_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _04067_, clk);
  dff _27262_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _04001_, clk);
  dff _27263_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _03999_, clk);
  dff _27264_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _12015_, clk);
  dff _27265_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _10717_, clk);
  dff _27266_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _10880_, clk);
  dff _27267_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _10935_, clk);
  dff _27268_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _03834_, clk);
  dff _27269_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _03857_, clk);
  dff _27270_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _02885_, clk);
  dff _27271_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _02948_, clk);
  dff _27272_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _03089_, clk);
  dff _27273_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _03075_, clk);
  dff _27274_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _03073_, clk);
  dff _27275_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _03064_, clk);
  dff _27276_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _12047_, clk);
  dff _27277_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _03203_, clk);
  dff _27278_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _03198_, clk);
  dff _27279_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _10712_, clk);
  dff _27280_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _12055_, clk);
  dff _27281_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _03101_, clk);
  dff _27282_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _12593_, clk);
  dff _27283_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _10813_, clk);
  dff _27284_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _10803_, clk);
  dff _27285_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _00796_, clk);
  dff _27286_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _00792_, clk);
  dff _27287_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _00785_, clk);
  dff _27288_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _00769_, clk);
  dff _27289_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _00767_, clk);
  dff _27290_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _12143_, clk);
  dff _27291_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _00933_, clk);
  dff _27292_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _00931_, clk);
  dff _27293_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _00884_, clk);
  dff _27294_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _00871_, clk);
  dff _27295_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _12139_, clk);
  dff _27296_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _10697_, clk);
  dff _27297_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _00483_, clk);
  dff _27298_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _00467_, clk);
  dff _27299_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _00462_, clk);
  dff _27300_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _10789_, clk);
  dff _27301_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _00253_, clk);
  dff _27302_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _00306_, clk);
  dff _27303_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _00302_, clk);
  dff _27304_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _00273_, clk);
  dff _27305_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _12157_, clk);
  dff _27306_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _10679_, clk);
  dff _27307_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _11164_, clk);
  dff _27308_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _11210_, clk);
  dff _27309_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _11201_, clk);
  dff _27310_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _11195_, clk);
  dff _27311_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _12202_, clk);
  dff _27312_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _00004_, clk);
  dff _27313_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _00038_, clk);
  dff _27314_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _00035_, clk);
  dff _27315_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _00028_, clk);
  dff _27316_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _10784_, clk);
  dff _27317_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _10517_, clk);
  dff _27318_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _10562_, clk);
  dff _27319_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _10567_, clk);
  dff _27320_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _12129_, clk);
  dff _27321_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _12107_, clk);
  dff _27322_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _12079_, clk);
  dff _27323_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _12076_, clk);
  dff _27324_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _12069_, clk);
  dff _27325_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _12685_, clk);
  dff _27326_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _12644_, clk);
  dff _27327_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _10558_, clk);
  dff _27328_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _11739_, clk);
  dff _27329_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _11733_, clk);
  dff _27330_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _10539_, clk);
  dff _27331_ (\oc8051_top_1.oc8051_memory_interface1.reti , _10663_, clk);
  dff _27332_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _11534_, clk);
  dff _27333_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _11531_, clk);
  dff _27334_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _11522_, clk);
  dff _27335_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _12600_, clk);
  dff _27336_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _12582_, clk);
  dff _27337_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _12721_, clk);
  dff _27338_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _11496_, clk);
  dff _27339_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _10654_, clk);
  dff _27340_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _10641_, clk);
  dff _27341_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _10620_, clk);
  dff _27342_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _11514_, clk);
  dff _27343_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _11509_, clk);
  dff _27344_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _11126_, clk);
  dff _27345_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _03099_, clk);
  dff _27346_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _11624_, clk);
  dff _27347_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _11121_, clk);
  dff _27348_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _11229_, clk);
  dff _27349_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _11270_, clk);
  dff _27350_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _11649_, clk);
  dff _27351_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _11643_, clk);
  dff _27352_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _11115_, clk);
  dff _27353_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _11663_, clk);
  dff _27354_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _11659_, clk);
  dff _27355_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _11112_, clk);
  dff _27356_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _11224_, clk);
  dff _27357_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _11674_, clk);
  dff _27358_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _11668_, clk);
  dff _27359_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _11707_, clk);
  dff _27360_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _11697_, clk);
  dff _27361_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _11095_, clk);
  dff _27362_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _11221_, clk);
  dff _27363_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _11267_, clk);
  dff _27364_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _11291_, clk);
  dff _27365_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _11364_, clk);
  dff _27366_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11361_, clk);
  dff _27367_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _11150_, clk);
  dff _27368_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _11390_, clk);
  dff _27369_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _11375_, clk);
  dff _27370_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _11148_, clk);
  dff _27371_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _11244_, clk);
  dff _27372_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _11352_, clk);
  dff _27373_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _11318_, clk);
  dff _27374_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _11154_, clk);
  dff _27375_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _11278_, clk);
  dff _27376_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _11413_, clk);
  dff _27377_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _02946_, clk);
  dff _27378_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _10400_, clk);
  dff _27379_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _03108_, clk);
  dff _27380_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _10460_, clk);
  dff _27381_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _11058_, clk);
  dff _27382_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _11285_, clk);
  dff _27383_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _11947_, clk);
  dff _27384_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _11940_, clk);
  dff _27385_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _10472_, clk);
  dff _27386_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0], clk);
  dff _27387_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1], clk);
  dff _27388_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2], clk);
  dff _27389_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3], clk);
  dff _27390_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4], clk);
  dff _27391_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5], clk);
  dff _27392_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6], clk);
  dff _27393_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7], clk);
  dff _27394_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8], clk);
  dff _27395_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9], clk);
  dff _27396_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10], clk);
  dff _27397_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11], clk);
  dff _27398_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12], clk);
  dff _27399_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13], clk);
  dff _27400_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14], clk);
  dff _27401_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15], clk);
  dff _27402_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16], clk);
  dff _27403_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17], clk);
  dff _27404_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18], clk);
  dff _27405_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19], clk);
  dff _27406_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20], clk);
  dff _27407_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21], clk);
  dff _27408_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22], clk);
  dff _27409_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23], clk);
  dff _27410_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24], clk);
  dff _27411_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25], clk);
  dff _27412_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26], clk);
  dff _27413_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27], clk);
  dff _27414_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28], clk);
  dff _27415_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29], clk);
  dff _27416_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30], clk);
  dff _27417_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31], clk);
  dff _27418_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _02407_, clk);
  dff _27419_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _03724_, clk);
  dff _27420_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _03769_, clk);
  dff _27421_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _03866_, clk);
  dff _27422_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _03706_, clk);
  dff _27423_ (\oc8051_top_1.oc8051_sfr1.bit_out , _03797_, clk);
  dff _27424_ (\oc8051_top_1.oc8051_sfr1.wait_data , _02476_, clk);
  dff _27425_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _03748_, clk);
  dff _27426_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _03766_, clk);
  dff _27427_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _03996_, clk);
  dff _27428_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _03992_, clk);
  dff _27429_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _04065_, clk);
  dff _27430_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _04003_, clk);
  dff _27431_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _03684_, clk);
  dff _27432_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _02423_, clk);
  dff _27433_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _03704_, clk);
  dff _27434_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _06484_, clk);
  dff _27435_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _03877_, clk);
  dff _27436_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _07042_, clk);
  dff _27437_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _03832_, clk);
  dff _27438_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _03309_, clk);
  dff _27439_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _06474_, clk);
  dff _27440_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _05109_, clk);
  dff _27441_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _05360_, clk);
  dff _27442_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _13347_, clk);
  dff _27443_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _02466_, clk);
  dff _27444_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _13360_, clk);
  dff _27445_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _13357_, clk);
  dff _27446_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _02463_, clk);
  dff _27447_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _13307_, clk);
  dff _27448_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _13293_, clk);
  dff _27449_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _03929_, clk);
  dff _27450_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _05691_, clk);
  dff _27451_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _05688_, clk);
  dff _27452_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _05680_, clk);
  dff _27453_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _05660_, clk);
  dff _27454_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _05657_, clk);
  dff _27455_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _05670_, clk);
  dff _27456_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _05665_, clk);
  dff _27457_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _01636_, clk);
  dff _27458_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _05775_, clk);
  dff _27459_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _01593_, clk);
  dff _27460_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _07867_, clk);
  dff _27461_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _05780_, clk);
  dff _27462_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _05772_, clk);
  dff _27463_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _01615_, clk);
  dff _27464_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _05783_, clk);
  dff _27465_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _01669_, clk);
  dff _27466_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _08294_, clk);
  dff _27467_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _01574_, clk);
  dff _27468_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _01571_, clk);
  dff _27469_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _01479_, clk);
  dff _27470_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _01590_, clk);
  dff _27471_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _01581_, clk);
  dff _27472_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _01478_, clk);
  dff _27473_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _01520_, clk);
  dff _27474_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _08055_, clk);
  dff _27475_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _01475_, clk);
  dff _27476_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _03130_, clk);
  dff _27477_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _07918_, clk);
  dff _27478_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _01527_, clk);
  dff _27479_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _01756_, clk);
  dff _27480_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _10256_, clk);
  dff _27481_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _01759_, clk);
  dff _27482_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _01471_, clk);
  dff _27483_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _10385_, clk);
  dff _27484_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _01763_, clk);
  dff _27485_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _01767_, clk);
  dff _27486_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _09243_, clk);
  dff _27487_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _07655_, clk);
  dff _27488_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _08980_, clk);
  dff _27489_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _07357_, clk);
  dff _27490_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _01522_, clk);
  dff _27491_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _01567_, clk);
  dff _27492_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _01565_, clk);
  dff _27493_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _07249_, clk);
  dff _27494_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _01795_, clk);
  dff _27495_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _01465_, clk);
  dff _27496_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _01801_, clk);
  dff _27497_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _01799_, clk);
  dff _27498_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _01463_, clk);
  dff _27499_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _01516_, clk);
  dff _27500_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _01804_, clk);
  dff _27501_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _10306_, clk);
  dff _27502_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _01812_, clk);
  dff _27503_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _01460_, clk);
  dff _27504_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _01826_, clk);
  dff _27505_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _01822_, clk);
  dff _27506_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _01459_, clk);
  dff _27507_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _01494_, clk);
  dff _27508_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _01845_, clk);
  dff _27509_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _10406_, clk);
  dff _27510_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _02690_, clk);
  dff _27511_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _02562_, clk);
  dff _27512_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _02525_, clk);
  dff _27513_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _02694_, clk);
  dff _27514_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _02565_, clk);
  dff _27515_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _02692_, clk);
  dff _27516_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _02559_, clk);
  dff _27517_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _01488_, clk);
  dff _27518_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _02555_, clk);
  dff _27519_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _02522_, clk);
  dff _27520_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _02700_, clk);
  dff _27521_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _02557_, clk);
  dff _27522_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _02698_, clk);
  dff _27523_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _02553_, clk);
  dff _27524_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _02520_, clk);
  dff _27525_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _02921_, clk);
  dff _27526_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _02696_, clk);
  dff _27527_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _02666_, clk);
  dff _27528_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _02656_, clk);
  dff _27529_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _02655_, clk);
  dff _27530_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _02549_, clk);
  dff _27531_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _02518_, clk);
  dff _27532_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _02704_, clk);
  dff _27533_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _03593_, clk);
  dff _27534_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _02702_, clk);
  dff _27535_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _02671_, clk);
  dff _27536_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _02668_, clk);
  dff _27537_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _02709_, clk);
  dff _27538_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _02547_, clk);
  dff _27539_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _02707_, clk);
  dff _27540_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _02677_, clk);
  dff _27541_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _03596_, clk);
  dff _27542_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _09234_, clk);
  dff _27543_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _01741_, clk);
  dff _27544_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _09629_, clk);
  dff _27545_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _09639_, clk);
  dff _27546_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _09636_, clk);
  dff _27547_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _09633_, clk);
  dff _27548_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _03196_, clk);
  dff _27549_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _12852_, clk);
  dff _27550_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _12846_, clk);
  dff _27551_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _12842_, clk);
  dff _27552_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _12840_, clk);
  dff _27553_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _02602_, clk);
  dff _27554_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _12781_, clk);
  dff _27555_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _12774_, clk);
  dff _27556_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _02472_, clk);
  dff _27557_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _13155_, clk);
  dff _27558_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _00411_, clk);
  dff _27559_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _00422_, clk);
  dff _27560_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _12133_, clk);
  dff _27561_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _12136_, clk);
  dff _27562_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _12116_, clk);
  dff _27563_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _12113_, clk);
  dff _27564_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _12110_, clk);
  dff _27565_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _12122_, clk);
  dff _27566_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _12085_, clk);
  dff _27567_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _00415_, clk);
  dff _27568_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _12152_, clk);
  dff _27569_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _12155_, clk);
  dff _27570_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _12170_, clk);
  dff _27571_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _12161_, clk);
  dff _27572_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _12167_, clk);
  dff _27573_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _12164_, clk);
  dff _27574_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _12238_, clk);
  dff _27575_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _00419_, clk);
  dff _27576_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _00417_, clk);
  dff _27577_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _00383_, clk);
  dff _27578_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _12174_, clk);
  dff _27579_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _12191_, clk);
  dff _27580_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _12199_, clk);
  dff _27581_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _12196_, clk);
  dff _27582_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _12251_, clk);
  dff _27583_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _12244_, clk);
  dff _27584_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _12247_, clk);
  dff _27585_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _00387_, clk);
  dff _27586_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _12348_, clk);
  dff _27587_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _12317_, clk);
  dff _27588_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _12320_, clk);
  dff _27589_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _12331_, clk);
  dff _27590_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _12335_, clk);
  dff _27591_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _12296_, clk);
  dff _27592_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _12293_, clk);
  dff _27593_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _00385_, clk);
  dff _27594_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _00399_, clk);
  dff _27595_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _12359_, clk);
  dff _27596_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _12375_, clk);
  dff _27597_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _12366_, clk);
  dff _27598_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _12372_, clk);
  dff _27599_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _12391_, clk);
  dff _27600_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _12383_, clk);
  dff _27601_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _12388_, clk);
  dff _27602_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _00395_, clk);
  dff _27603_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01940_, clk);
  dff _27604_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01937_, clk);
  dff _27605_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01934_, clk);
  dff _27606_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01931_, clk);
  dff _27607_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _05216_, clk);
  dff _27608_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _12309_, clk);
  dff _27609_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _12306_, clk);
  dff _27610_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _12302_, clk);
  dff _27611_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _12299_, clk);
  dff _27612_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _07864_, clk);
  dff _27613_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _12342_, clk);
  dff _27614_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01860_, clk);
  dff _27615_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _12271_, clk);
  dff _27616_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _12267_, clk);
  dff _27617_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _07878_, clk);
  dff _27618_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _11138_, clk);
  dff _27619_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _12206_, clk);
  dff _27620_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _07900_, clk);
  dff _27621_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _12218_, clk);
  dff _27622_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01920_, clk);
  dff _27623_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01917_, clk);
  dff _27624_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _01752_, clk);
  dff _27625_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _09843_, clk);
  dff _27626_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _10730_, clk);
  dff _27627_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _10755_, clk);
  dff _27628_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _10746_, clk);
  dff _27629_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _10739_, clk);
  dff _27630_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _10736_, clk);
  dff _27631_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01914_, clk);
  dff _27632_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _10660_, clk);
  dff _27633_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _10649_, clk);
  dff _27634_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _10645_, clk);
  dff _27635_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _12226_, clk);
  dff _27636_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _10684_, clk);
  dff _27637_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _10709_, clk);
  dff _27638_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _10705_, clk);
  dff _27639_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01911_, clk);
  dff _27640_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01908_, clk);
  dff _27641_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _10524_, clk);
  dff _27642_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _12261_, clk);
  dff _27643_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _10600_, clk);
  dff _27644_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _10597_, clk);
  dff _27645_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _10587_, clk);
  dff _27646_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _10585_, clk);
  dff _27647_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _10582_, clk);
  dff _27648_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01851_, clk);
  dff _27649_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _03173_, clk);
  dff _27650_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _03170_, clk);
  dff _27651_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _03167_, clk);
  dff _27652_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _03165_, clk);
  dff _27653_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _03153_, clk);
  dff _27654_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _03151_, clk);
  dff _27655_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _03149_, clk);
  dff _27656_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _03147_, clk);
  dff _27657_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _03145_, clk);
  dff _27658_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _03143_, clk);
  dff _27659_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _03135_, clk);
  dff _27660_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _03191_, clk);
  dff _27661_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _09231_, clk);
  dff _27662_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _10104_, clk);
  dff _27663_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _01600_, clk);
  dff _27664_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _03686_, clk);
  dff _27665_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _03659_, clk);
  dff _27666_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _03599_, clk);
  dff _27667_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _03114_, clk);
  dff _27668_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _03571_, clk);
  dff _27669_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _03994_, clk);
  dff _27670_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _07758_, clk);
  dff _27671_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01619_, clk);
  dff _27672_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _03532_, clk);
  dff _27673_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _03112_, clk);
  dff _27674_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _02503_, clk);
  dff _27675_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01513_, clk);
  dff _27676_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01500_, clk);
  dff _27677_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01498_, clk);
  dff _27678_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01447_, clk);
  dff _27679_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _08247_, clk);
  dff _27680_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _03193_, clk);
  dff _27681_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _03186_, clk);
  dff _27682_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _03155_, clk);
  dff _27683_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _03085_, clk);
  dff _27684_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _03059_, clk);
  dff _27685_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _07189_, clk);
  dff _27686_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _07175_, clk);
  dff _27687_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _08250_, clk);
  dff _27688_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _02897_, clk);
  dff _27689_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _10942_, clk);
  dff _27690_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _07036_, clk);
  dff _27691_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _10974_, clk);
  dff _27692_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _10966_, clk);
  dff _27693_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _11006_, clk);
  dff _27694_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _10985_, clk);
  dff _27695_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _11161_, clk);
  dff _27696_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _11073_, clk);
  dff _27697_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _12398_, clk);
  dff _27698_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _11983_, clk);
  dff _27699_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _02878_, clk);
  dff _27700_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _00031_, clk);
  dff _27701_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _12951_, clk);
  dff _27702_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _00263_, clk);
  dff _27703_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _00128_, clk);
  dff _27704_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _06965_, clk);
  dff _27705_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _00472_, clk);
  dff _27706_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _00451_, clk);
  dff _27707_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _02688_, clk);
  dff _27708_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01043_, clk);
  dff _27709_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _00929_, clk);
  dff _27710_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _06961_, clk);
  dff _27711_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01468_, clk);
  dff _27712_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01453_, clk);
  dff _27713_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _07022_, clk);
  dff _27714_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _07047_, clk);
  dff _27715_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _02626_, clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [0], ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [1], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [2], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [3], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [4], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [5], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [6], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [7], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [8], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [9], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [10], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [11], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [12], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [13], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [14], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [15], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [16], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [0], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [1], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [2], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [3], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [4], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [5], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [6], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [7], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [0], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [1], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [2], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [3], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [4], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [5], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [6], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [7], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.mulOv , ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [0], ABINPUT000000[1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [1], ABINPUT000000[2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [2], ABINPUT000000[3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [3], ABINPUT000000[4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [4], ABINPUT000000[5]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [5], ABINPUT000000[6]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [6], ABINPUT000000[7]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [7], ABINPUT000000[8]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [0], ABINPUT000000[9]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [1], ABINPUT000000[10]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], ABINPUT000000[11]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], ABINPUT000000[12]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], ABINPUT000000[13]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], ABINPUT000000[14]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], ABINPUT000000[15]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], ABINPUT000000[16]);
  buf(\oc8051_top_1.oc8051_alu1.divOv , ABINPUT000000[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [0], ABINPUT000000[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [1], ABINPUT000000[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [2], ABINPUT000000[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [3], ABINPUT000000[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [4], ABINPUT000000[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [5], ABINPUT000000[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [6], ABINPUT000000[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [7], ABINPUT000000[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [8], ABINPUT000000[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [9], ABINPUT000000[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [10], ABINPUT000000[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [11], ABINPUT000000[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [12], ABINPUT000000[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [13], ABINPUT000000[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [14], ABINPUT000000[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [15], ABINPUT000000[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [16], ABINPUT000000[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.ABINPUT000 [0], ABINPUT000[0]);
  buf(\oc8051_top_1.ABINPUT000 [1], ABINPUT000[1]);
  buf(\oc8051_top_1.ABINPUT000 [2], ABINPUT000[2]);
  buf(\oc8051_top_1.ABINPUT000 [3], ABINPUT000[3]);
  buf(\oc8051_top_1.ABINPUT000 [4], ABINPUT000[4]);
  buf(\oc8051_top_1.ABINPUT000 [5], ABINPUT000[5]);
  buf(\oc8051_top_1.ABINPUT000 [6], ABINPUT000[6]);
  buf(\oc8051_top_1.ABINPUT000 [7], ABINPUT000[7]);
  buf(\oc8051_top_1.ABINPUT000 [8], ABINPUT000[8]);
  buf(\oc8051_top_1.ABINPUT000 [9], ABINPUT000[9]);
  buf(\oc8051_top_1.ABINPUT000 [10], ABINPUT000[10]);
  buf(\oc8051_top_1.ABINPUT000 [11], ABINPUT000[11]);
  buf(\oc8051_top_1.ABINPUT000 [12], ABINPUT000[12]);
  buf(\oc8051_top_1.ABINPUT000 [13], ABINPUT000[13]);
  buf(\oc8051_top_1.ABINPUT000 [14], ABINPUT000[14]);
  buf(\oc8051_top_1.ABINPUT000 [15], ABINPUT000[15]);
  buf(\oc8051_top_1.ABINPUT000 [16], ABINPUT000[16]);
  buf(\oc8051_top_1.ABINPUT000000 [0], ABINPUT000000[0]);
  buf(\oc8051_top_1.ABINPUT000000 [1], ABINPUT000000[1]);
  buf(\oc8051_top_1.ABINPUT000000 [2], ABINPUT000000[2]);
  buf(\oc8051_top_1.ABINPUT000000 [3], ABINPUT000000[3]);
  buf(\oc8051_top_1.ABINPUT000000 [4], ABINPUT000000[4]);
  buf(\oc8051_top_1.ABINPUT000000 [5], ABINPUT000000[5]);
  buf(\oc8051_top_1.ABINPUT000000 [6], ABINPUT000000[6]);
  buf(\oc8051_top_1.ABINPUT000000 [7], ABINPUT000000[7]);
  buf(\oc8051_top_1.ABINPUT000000 [8], ABINPUT000000[8]);
  buf(\oc8051_top_1.ABINPUT000000 [9], ABINPUT000000[9]);
  buf(\oc8051_top_1.ABINPUT000000 [10], ABINPUT000000[10]);
  buf(\oc8051_top_1.ABINPUT000000 [11], ABINPUT000000[11]);
  buf(\oc8051_top_1.ABINPUT000000 [12], ABINPUT000000[12]);
  buf(\oc8051_top_1.ABINPUT000000 [13], ABINPUT000000[13]);
  buf(\oc8051_top_1.ABINPUT000000 [14], ABINPUT000000[14]);
  buf(\oc8051_top_1.ABINPUT000000 [15], ABINPUT000000[15]);
  buf(\oc8051_top_1.ABINPUT000000 [16], ABINPUT000000[16]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.decoder_new_valid_pc , pc_log_change);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log_change , pc_log_change);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
