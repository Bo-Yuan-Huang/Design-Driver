
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_pc, ABINPUT, ABINPUT000, ABINPUT001, ABINPUT002, ABINPUT003, ABINPUT004, ABINPUT005, ABINPUT006, ABINPUT007, ABINPUT008, ABINPUT009);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire [7:0] _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire [7:0] _30753_;
  wire [7:0] _30754_;
  wire [7:0] _30755_;
  wire [7:0] _30756_;
  wire [7:0] _30757_;
  wire [7:0] _30758_;
  wire [7:0] _30759_;
  wire [7:0] _30760_;
  wire [7:0] _30761_;
  wire [7:0] _30762_;
  input [34:0] ABINPUT;
  input [7:0] ABINPUT000;
  input [7:0] ABINPUT001;
  input [7:0] ABINPUT002;
  input [7:0] ABINPUT003;
  input [7:0] ABINPUT004;
  input [7:0] ABINPUT005;
  input [7:0] ABINPUT006;
  input [7:0] ABINPUT007;
  input [7:0] ABINPUT008;
  input [127:0] ABINPUT009;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IP_gm;
  wire [127:0] IRAM_gm;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PSW_gm;
  wire [7:0] PSW_gm_next;
  wire [7:0] SBUF_gm;
  wire [7:0] SCON_gm;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TH0_gm;
  wire [7:0] TH1_gm;
  wire [7:0] TL0_gm;
  wire [7:0] TL1_gm;
  wire [7:0] TMOD_gm;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire eq_state;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT000 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT001 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT002 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT003 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT004 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT005 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT006 ;
  wire [7:0] \oc8051_golden_model_1.ABINPUT007 ;
  wire [127:0] \oc8051_golden_model_1.ABINPUT008 ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_next ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.B_next ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPH_next ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.DPL_next ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [127:0] \oc8051_golden_model_1.IRAM_full ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P0_next ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P1_next ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P2_next ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [7:0] \oc8051_golden_model_1.P3_next ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_fa ;
  wire [7:0] \oc8051_golden_model_1.PSW_fb ;
  wire [7:0] \oc8051_golden_model_1.PSW_fc ;
  wire [7:0] \oc8051_golden_model_1.PSW_fd ;
  wire [7:0] \oc8051_golden_model_1.PSW_fe ;
  wire [7:0] \oc8051_golden_model_1.PSW_ff ;
  wire [7:0] \oc8051_golden_model_1.PSW_next ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0573 ;
  wire [7:0] \oc8051_golden_model_1.n0606 ;
  wire [15:0] \oc8051_golden_model_1.n0713 ;
  wire [15:0] \oc8051_golden_model_1.n0745 ;
  wire [15:0] \oc8051_golden_model_1.n1004 ;
  wire [6:0] \oc8051_golden_model_1.n1008 ;
  wire \oc8051_golden_model_1.n1009 ;
  wire \oc8051_golden_model_1.n1010 ;
  wire \oc8051_golden_model_1.n1011 ;
  wire \oc8051_golden_model_1.n1012 ;
  wire \oc8051_golden_model_1.n1013 ;
  wire \oc8051_golden_model_1.n1014 ;
  wire \oc8051_golden_model_1.n1015 ;
  wire \oc8051_golden_model_1.n1016 ;
  wire \oc8051_golden_model_1.n1023 ;
  wire [7:0] \oc8051_golden_model_1.n1024 ;
  wire [7:0] \oc8051_golden_model_1.n1031 ;
  wire \oc8051_golden_model_1.n1032 ;
  wire \oc8051_golden_model_1.n1033 ;
  wire \oc8051_golden_model_1.n1034 ;
  wire \oc8051_golden_model_1.n1035 ;
  wire \oc8051_golden_model_1.n1036 ;
  wire \oc8051_golden_model_1.n1037 ;
  wire \oc8051_golden_model_1.n1038 ;
  wire \oc8051_golden_model_1.n1039 ;
  wire [7:0] \oc8051_golden_model_1.n1047 ;
  wire [7:0] \oc8051_golden_model_1.n1064 ;
  wire [3:0] \oc8051_golden_model_1.n1157 ;
  wire [3:0] \oc8051_golden_model_1.n1159 ;
  wire [3:0] \oc8051_golden_model_1.n1161 ;
  wire [3:0] \oc8051_golden_model_1.n1162 ;
  wire [3:0] \oc8051_golden_model_1.n1163 ;
  wire [3:0] \oc8051_golden_model_1.n1164 ;
  wire [3:0] \oc8051_golden_model_1.n1165 ;
  wire [3:0] \oc8051_golden_model_1.n1166 ;
  wire [3:0] \oc8051_golden_model_1.n1167 ;
  wire \oc8051_golden_model_1.n1259 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1261 ;
  wire [7:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [2:0] \oc8051_golden_model_1.n1264 ;
  wire \oc8051_golden_model_1.n1265 ;
  wire [1:0] \oc8051_golden_model_1.n1266 ;
  wire [7:0] \oc8051_golden_model_1.n1267 ;
  wire [6:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1269 ;
  wire \oc8051_golden_model_1.n1270 ;
  wire \oc8051_golden_model_1.n1271 ;
  wire \oc8051_golden_model_1.n1272 ;
  wire \oc8051_golden_model_1.n1273 ;
  wire \oc8051_golden_model_1.n1274 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire \oc8051_golden_model_1.n1276 ;
  wire [7:0] \oc8051_golden_model_1.n1284 ;
  wire [7:0] \oc8051_golden_model_1.n1301 ;
  wire [15:0] \oc8051_golden_model_1.n1343 ;
  wire [7:0] \oc8051_golden_model_1.n1345 ;
  wire \oc8051_golden_model_1.n1346 ;
  wire \oc8051_golden_model_1.n1347 ;
  wire \oc8051_golden_model_1.n1348 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire \oc8051_golden_model_1.n1350 ;
  wire \oc8051_golden_model_1.n1351 ;
  wire \oc8051_golden_model_1.n1352 ;
  wire \oc8051_golden_model_1.n1353 ;
  wire [7:0] \oc8051_golden_model_1.n1361 ;
  wire [8:0] \oc8051_golden_model_1.n1363 ;
  wire [3:0] \oc8051_golden_model_1.n1369 ;
  wire [4:0] \oc8051_golden_model_1.n1370 ;
  wire [8:0] \oc8051_golden_model_1.n1376 ;
  wire [7:0] \oc8051_golden_model_1.n1385 ;
  wire [6:0] \oc8051_golden_model_1.n1386 ;
  wire [7:0] \oc8051_golden_model_1.n1402 ;
  wire [7:0] \oc8051_golden_model_1.n1440 ;
  wire [6:0] \oc8051_golden_model_1.n1441 ;
  wire [7:0] \oc8051_golden_model_1.n1457 ;
  wire [8:0] \oc8051_golden_model_1.n1459 ;
  wire [3:0] \oc8051_golden_model_1.n1463 ;
  wire [4:0] \oc8051_golden_model_1.n1464 ;
  wire [4:0] \oc8051_golden_model_1.n1466 ;
  wire \oc8051_golden_model_1.n1467 ;
  wire [8:0] \oc8051_golden_model_1.n1468 ;
  wire [7:0] \oc8051_golden_model_1.n1476 ;
  wire [6:0] \oc8051_golden_model_1.n1477 ;
  wire \oc8051_golden_model_1.n1492 ;
  wire [7:0] \oc8051_golden_model_1.n1493 ;
  wire [7:0] \oc8051_golden_model_1.n1505 ;
  wire [6:0] \oc8051_golden_model_1.n1506 ;
  wire [7:0] \oc8051_golden_model_1.n1507 ;
  wire [8:0] \oc8051_golden_model_1.n1509 ;
  wire [8:0] \oc8051_golden_model_1.n1511 ;
  wire \oc8051_golden_model_1.n1512 ;
  wire [4:0] \oc8051_golden_model_1.n1513 ;
  wire [4:0] \oc8051_golden_model_1.n1515 ;
  wire \oc8051_golden_model_1.n1516 ;
  wire [8:0] \oc8051_golden_model_1.n1517 ;
  wire \oc8051_golden_model_1.n1524 ;
  wire [7:0] \oc8051_golden_model_1.n1525 ;
  wire [6:0] \oc8051_golden_model_1.n1526 ;
  wire \oc8051_golden_model_1.n1541 ;
  wire [7:0] \oc8051_golden_model_1.n1542 ;
  wire [4:0] \oc8051_golden_model_1.n1544 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [6:0] \oc8051_golden_model_1.n1547 ;
  wire [7:0] \oc8051_golden_model_1.n1548 ;
  wire [8:0] \oc8051_golden_model_1.n1550 ;
  wire \oc8051_golden_model_1.n1551 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire [7:0] \oc8051_golden_model_1.n1559 ;
  wire [6:0] \oc8051_golden_model_1.n1560 ;
  wire [7:0] \oc8051_golden_model_1.n1561 ;
  wire [7:0] \oc8051_golden_model_1.n1562 ;
  wire [6:0] \oc8051_golden_model_1.n1563 ;
  wire [7:0] \oc8051_golden_model_1.n1564 ;
  wire [8:0] \oc8051_golden_model_1.n1567 ;
  wire [8:0] \oc8051_golden_model_1.n1568 ;
  wire [7:0] \oc8051_golden_model_1.n1569 ;
  wire [7:0] \oc8051_golden_model_1.n1570 ;
  wire [6:0] \oc8051_golden_model_1.n1571 ;
  wire \oc8051_golden_model_1.n1572 ;
  wire \oc8051_golden_model_1.n1573 ;
  wire \oc8051_golden_model_1.n1574 ;
  wire \oc8051_golden_model_1.n1575 ;
  wire \oc8051_golden_model_1.n1576 ;
  wire \oc8051_golden_model_1.n1577 ;
  wire \oc8051_golden_model_1.n1578 ;
  wire \oc8051_golden_model_1.n1579 ;
  wire [7:0] \oc8051_golden_model_1.n1587 ;
  wire [7:0] \oc8051_golden_model_1.n1588 ;
  wire [8:0] \oc8051_golden_model_1.n1591 ;
  wire [4:0] \oc8051_golden_model_1.n1595 ;
  wire [7:0] \oc8051_golden_model_1.n1606 ;
  wire [6:0] \oc8051_golden_model_1.n1607 ;
  wire [7:0] \oc8051_golden_model_1.n1623 ;
  wire [7:0] \oc8051_golden_model_1.n1639 ;
  wire [6:0] \oc8051_golden_model_1.n1640 ;
  wire [7:0] \oc8051_golden_model_1.n1656 ;
  wire [8:0] \oc8051_golden_model_1.n1660 ;
  wire \oc8051_golden_model_1.n1661 ;
  wire [4:0] \oc8051_golden_model_1.n1663 ;
  wire \oc8051_golden_model_1.n1664 ;
  wire \oc8051_golden_model_1.n1671 ;
  wire [7:0] \oc8051_golden_model_1.n1672 ;
  wire [6:0] \oc8051_golden_model_1.n1673 ;
  wire \oc8051_golden_model_1.n1688 ;
  wire [7:0] \oc8051_golden_model_1.n1689 ;
  wire [8:0] \oc8051_golden_model_1.n1693 ;
  wire \oc8051_golden_model_1.n1694 ;
  wire [4:0] \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1697 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire [6:0] \oc8051_golden_model_1.n1706 ;
  wire \oc8051_golden_model_1.n1721 ;
  wire [7:0] \oc8051_golden_model_1.n1722 ;
  wire [7:0] \oc8051_golden_model_1.n1749 ;
  wire \oc8051_golden_model_1.n1804 ;
  wire [7:0] \oc8051_golden_model_1.n1805 ;
  wire \oc8051_golden_model_1.n1821 ;
  wire [7:0] \oc8051_golden_model_1.n1822 ;
  wire \oc8051_golden_model_1.n1838 ;
  wire [7:0] \oc8051_golden_model_1.n1839 ;
  wire \oc8051_golden_model_1.n1855 ;
  wire [7:0] \oc8051_golden_model_1.n1856 ;
  wire [7:0] \oc8051_golden_model_1.n1881 ;
  wire [7:0] \oc8051_golden_model_1.n1937 ;
  wire [7:0] \oc8051_golden_model_1.n1954 ;
  wire \oc8051_golden_model_1.n1970 ;
  wire [7:0] \oc8051_golden_model_1.n1971 ;
  wire \oc8051_golden_model_1.n1987 ;
  wire [7:0] \oc8051_golden_model_1.n1988 ;
  wire [7:0] \oc8051_golden_model_1.n2086 ;
  wire [7:0] \oc8051_golden_model_1.n2103 ;
  wire \oc8051_golden_model_1.n2119 ;
  wire [7:0] \oc8051_golden_model_1.n2120 ;
  wire \oc8051_golden_model_1.n2136 ;
  wire [7:0] \oc8051_golden_model_1.n2137 ;
  wire [6:0] \oc8051_golden_model_1.n2142 ;
  wire [7:0] \oc8051_golden_model_1.n2143 ;
  wire [6:0] \oc8051_golden_model_1.n2144 ;
  wire [7:0] \oc8051_golden_model_1.n2145 ;
  wire \oc8051_golden_model_1.n2160 ;
  wire [7:0] \oc8051_golden_model_1.n2161 ;
  wire \oc8051_golden_model_1.n2200 ;
  wire [7:0] \oc8051_golden_model_1.n2201 ;
  wire [6:0] \oc8051_golden_model_1.n2202 ;
  wire [7:0] \oc8051_golden_model_1.n2203 ;
  wire [3:0] \oc8051_golden_model_1.n2210 ;
  wire \oc8051_golden_model_1.n2211 ;
  wire [7:0] \oc8051_golden_model_1.n2212 ;
  wire [6:0] \oc8051_golden_model_1.n2213 ;
  wire \oc8051_golden_model_1.n2228 ;
  wire [7:0] \oc8051_golden_model_1.n2229 ;
  wire [7:0] \oc8051_golden_model_1.n2441 ;
  wire [7:0] \oc8051_golden_model_1.n2453 ;
  wire [6:0] \oc8051_golden_model_1.n2454 ;
  wire \oc8051_golden_model_1.n2469 ;
  wire [7:0] \oc8051_golden_model_1.n2470 ;
  wire \oc8051_golden_model_1.n2474 ;
  wire \oc8051_golden_model_1.n2476 ;
  wire \oc8051_golden_model_1.n2482 ;
  wire [7:0] \oc8051_golden_model_1.n2483 ;
  wire [6:0] \oc8051_golden_model_1.n2484 ;
  wire \oc8051_golden_model_1.n2499 ;
  wire [7:0] \oc8051_golden_model_1.n2500 ;
  wire \oc8051_golden_model_1.n2504 ;
  wire \oc8051_golden_model_1.n2506 ;
  wire \oc8051_golden_model_1.n2512 ;
  wire [7:0] \oc8051_golden_model_1.n2513 ;
  wire [6:0] \oc8051_golden_model_1.n2514 ;
  wire \oc8051_golden_model_1.n2529 ;
  wire [7:0] \oc8051_golden_model_1.n2530 ;
  wire \oc8051_golden_model_1.n2534 ;
  wire \oc8051_golden_model_1.n2536 ;
  wire \oc8051_golden_model_1.n2542 ;
  wire [7:0] \oc8051_golden_model_1.n2543 ;
  wire [6:0] \oc8051_golden_model_1.n2544 ;
  wire \oc8051_golden_model_1.n2559 ;
  wire [7:0] \oc8051_golden_model_1.n2560 ;
  wire [7:0] \oc8051_golden_model_1.n2563 ;
  wire [6:0] \oc8051_golden_model_1.n2564 ;
  wire [7:0] \oc8051_golden_model_1.n2565 ;
  wire [7:0] \oc8051_golden_model_1.n2566 ;
  wire [6:0] \oc8051_golden_model_1.n2567 ;
  wire [7:0] \oc8051_golden_model_1.n2568 ;
  wire [15:0] \oc8051_golden_model_1.n2572 ;
  wire \oc8051_golden_model_1.n2578 ;
  wire [7:0] \oc8051_golden_model_1.n2579 ;
  wire [6:0] \oc8051_golden_model_1.n2580 ;
  wire \oc8051_golden_model_1.n2595 ;
  wire [7:0] \oc8051_golden_model_1.n2596 ;
  wire \oc8051_golden_model_1.n2599 ;
  wire [7:0] \oc8051_golden_model_1.n2600 ;
  wire [6:0] \oc8051_golden_model_1.n2601 ;
  wire [7:0] \oc8051_golden_model_1.n2602 ;
  wire \oc8051_golden_model_1.n2634 ;
  wire [7:0] \oc8051_golden_model_1.n2635 ;
  wire [6:0] \oc8051_golden_model_1.n2636 ;
  wire [7:0] \oc8051_golden_model_1.n2637 ;
  wire \oc8051_golden_model_1.n2642 ;
  wire [7:0] \oc8051_golden_model_1.n2643 ;
  wire [6:0] \oc8051_golden_model_1.n2644 ;
  wire [7:0] \oc8051_golden_model_1.n2645 ;
  wire \oc8051_golden_model_1.n2650 ;
  wire [7:0] \oc8051_golden_model_1.n2651 ;
  wire [6:0] \oc8051_golden_model_1.n2652 ;
  wire [7:0] \oc8051_golden_model_1.n2653 ;
  wire \oc8051_golden_model_1.n2658 ;
  wire [7:0] \oc8051_golden_model_1.n2659 ;
  wire [6:0] \oc8051_golden_model_1.n2660 ;
  wire [7:0] \oc8051_golden_model_1.n2661 ;
  wire \oc8051_golden_model_1.n2666 ;
  wire [7:0] \oc8051_golden_model_1.n2667 ;
  wire [6:0] \oc8051_golden_model_1.n2668 ;
  wire [7:0] \oc8051_golden_model_1.n2669 ;
  wire [7:0] \oc8051_golden_model_1.n2694 ;
  wire [6:0] \oc8051_golden_model_1.n2695 ;
  wire [7:0] \oc8051_golden_model_1.n2696 ;
  wire [3:0] \oc8051_golden_model_1.n2697 ;
  wire [7:0] \oc8051_golden_model_1.n2698 ;
  wire \oc8051_golden_model_1.n2699 ;
  wire \oc8051_golden_model_1.n2700 ;
  wire \oc8051_golden_model_1.n2701 ;
  wire \oc8051_golden_model_1.n2702 ;
  wire \oc8051_golden_model_1.n2703 ;
  wire \oc8051_golden_model_1.n2704 ;
  wire \oc8051_golden_model_1.n2705 ;
  wire \oc8051_golden_model_1.n2706 ;
  wire \oc8051_golden_model_1.n2713 ;
  wire [7:0] \oc8051_golden_model_1.n2714 ;
  wire \oc8051_golden_model_1.n2752 ;
  wire \oc8051_golden_model_1.n2753 ;
  wire \oc8051_golden_model_1.n2754 ;
  wire \oc8051_golden_model_1.n2755 ;
  wire \oc8051_golden_model_1.n2756 ;
  wire \oc8051_golden_model_1.n2757 ;
  wire \oc8051_golden_model_1.n2758 ;
  wire \oc8051_golden_model_1.n2759 ;
  wire \oc8051_golden_model_1.n2766 ;
  wire [7:0] \oc8051_golden_model_1.n2767 ;
  wire \oc8051_golden_model_1.n2768 ;
  wire \oc8051_golden_model_1.n2769 ;
  wire \oc8051_golden_model_1.n2770 ;
  wire \oc8051_golden_model_1.n2771 ;
  wire \oc8051_golden_model_1.n2772 ;
  wire \oc8051_golden_model_1.n2773 ;
  wire \oc8051_golden_model_1.n2774 ;
  wire \oc8051_golden_model_1.n2775 ;
  wire \oc8051_golden_model_1.n2782 ;
  wire [7:0] \oc8051_golden_model_1.n2783 ;
  wire [7:0] \oc8051_golden_model_1.n2815 ;
  wire [6:0] \oc8051_golden_model_1.n2816 ;
  wire [7:0] \oc8051_golden_model_1.n2817 ;
  wire \oc8051_golden_model_1.n2836 ;
  wire [7:0] \oc8051_golden_model_1.n2837 ;
  wire [6:0] \oc8051_golden_model_1.n2838 ;
  wire [7:0] \oc8051_golden_model_1.n2854 ;
  wire [7:0] \oc8051_golden_model_1.n2858 ;
  wire [3:0] \oc8051_golden_model_1.n2859 ;
  wire [7:0] \oc8051_golden_model_1.n2860 ;
  wire \oc8051_golden_model_1.n2861 ;
  wire \oc8051_golden_model_1.n2862 ;
  wire \oc8051_golden_model_1.n2863 ;
  wire \oc8051_golden_model_1.n2864 ;
  wire \oc8051_golden_model_1.n2865 ;
  wire \oc8051_golden_model_1.n2866 ;
  wire \oc8051_golden_model_1.n2867 ;
  wire \oc8051_golden_model_1.n2868 ;
  wire [7:0] \oc8051_golden_model_1.n2876 ;
  wire \oc8051_golden_model_1.n2894 ;
  wire [7:0] \oc8051_golden_model_1.n2895 ;
  wire [7:0] \oc8051_golden_model_1.n2896 ;
  wire \oc8051_golden_model_1.n2912 ;
  wire [7:0] \oc8051_golden_model_1.n2913 ;
  wire \oc8051_golden_model_1.rst ;
  wire [34:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.des1 ;
  wire [7:0] \oc8051_top_1.des2 ;
  wire \oc8051_top_1.desAc ;
  wire \oc8051_top_1.desCy ;
  wire \oc8051_top_1.desOv ;
  wire [7:0] \oc8051_top_1.des_acc ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire [7:0] \oc8051_top_1.ie ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.des ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.data_in ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.alu ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des1 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des2 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des_acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.wr_dat ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_data_in ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat2 ;
  wire \oc8051_top_1.oc8051_sfr1.desAc ;
  wire \oc8051_top_1.oc8051_sfr1.desOv ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.des_acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire [7:0] \oc8051_top_1.sub_result ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire [7:0] \oc8051_top_1.wr_dat ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire p1_valid_r;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_pc;
  wire property_valid_psw_1_r;
  wire property_valid_sp_1_r;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  wire regs_always_zero;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_27053_, rst);
  not (_16883_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_16893_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_16904_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _16893_);
  and (_16915_, _16904_, _16883_);
  and (_16926_, \oc8051_top_1.oc8051_decoder1.wr , _16893_);
  not (_16937_, _16926_);
  nor (_16948_, _16937_, _16915_);
  and (_16959_, _16948_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_16970_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _16893_);
  and (_16980_, _16970_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_16991_, _16980_, _16883_);
  not (_17002_, _16991_);
  not (_17013_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and (_17024_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_17035_, _17024_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_17046_, _17035_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_17057_, _17046_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_17067_, _17057_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_17078_, _17067_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_17089_, _17078_, _17013_);
  and (_17100_, _17078_, _17013_);
  nor (_17111_, _17100_, _17089_);
  nor (_17122_, _17111_, _17002_);
  not (_17133_, _17122_);
  nor (_17144_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_17154_, _17144_, _16904_);
  and (_17165_, _17154_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not (_17176_, _17165_);
  and (_17187_, _16980_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_17198_, _17187_);
  not (_17209_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_17220_, _16970_, _17209_);
  and (_17231_, _17220_, _16883_);
  and (_17241_, _17231_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and (_17252_, _17220_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_17263_, _17252_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_17274_, _17263_, _17241_);
  and (_17285_, _17274_, _17198_);
  and (_17296_, _17285_, _17176_);
  and (_17307_, _17296_, _17133_);
  not (_17318_, _17307_);
  not (_17328_, _17067_);
  nor (_17339_, _17057_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_17350_, _17339_, _17002_);
  and (_17361_, _17350_, _17328_);
  not (_17372_, _17361_);
  and (_17383_, _17252_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_17394_, _17383_, _17187_);
  and (_17405_, _17154_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_17415_, _17231_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_17426_, _17415_, _17405_);
  and (_17437_, _17426_, _17394_);
  and (_17448_, _17437_, _17372_);
  not (_17469_, _17078_);
  nor (_17470_, _17067_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_17481_, _17470_, _17002_);
  and (_17492_, _17481_, _17469_);
  not (_17502_, _17492_);
  and (_17513_, _17231_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_17524_, _17513_, _17187_);
  and (_17535_, _17154_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_17546_, _17252_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_17557_, _17546_, _17535_);
  and (_17568_, _17557_, _17524_);
  and (_17579_, _17568_, _17502_);
  nor (_17589_, _17579_, _17448_);
  and (_17600_, _17252_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_17611_, _17231_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_17622_, _17611_, _17600_);
  nor (_17633_, _17035_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_17644_, _17633_, _17046_);
  and (_17655_, _17644_, _16991_);
  not (_17666_, _17655_);
  nor (_17676_, _17144_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_17687_, _17676_, _16904_);
  and (_17698_, _17687_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_17709_, _17154_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_17720_, _17709_, _17698_);
  and (_17731_, _17720_, _17666_);
  and (_17742_, _17731_, _17622_);
  not (_17753_, _17742_);
  not (_17763_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_17774_, _17046_, _17763_);
  nor (_17785_, _17046_, _17763_);
  nor (_17796_, _17785_, _17774_);
  nor (_17807_, _17796_, _17002_);
  not (_17818_, _17807_);
  and (_17829_, _17252_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_17840_, _17829_, _17187_);
  and (_17850_, _17687_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_17861_, _17154_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_17872_, _17861_, _17850_);
  and (_17893_, _17231_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  not (_17894_, _17893_);
  and (_17905_, _17894_, _17872_);
  and (_17916_, _17905_, _17840_);
  and (_17937_, _17916_, _17818_);
  nor (_17938_, _17937_, _17753_);
  and (_17949_, _17938_, _17589_);
  and (_17960_, _17949_, _17318_);
  nor (_17971_, _17024_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_17982_, _17971_, _17035_);
  and (_17993_, _17982_, _16991_);
  and (_18004_, _17154_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_18015_, _18004_, _17993_);
  and (_18026_, _17252_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_18037_, _17231_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_18048_, _17687_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_18059_, _18048_, _18037_);
  nor (_18070_, _18059_, _18026_);
  and (_18081_, _18070_, _18015_);
  not (_18092_, _18081_);
  and (_18103_, _17231_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_18114_, _17154_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_18124_, _18114_, _18103_);
  and (_18135_, _17252_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not (_18146_, _18135_);
  not (_18157_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_18168_, _16991_, _18157_);
  and (_18179_, _17687_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_18190_, _18179_, _18168_);
  and (_18201_, _18190_, _18146_);
  and (_18212_, _18201_, _18124_);
  and (_18223_, _17252_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor (_18234_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_18245_, _18234_, _17024_);
  and (_18256_, _18245_, _16991_);
  nor (_18267_, _18256_, _18223_);
  and (_18278_, _17154_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and (_18289_, _17687_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_18300_, _17231_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or (_18311_, _18300_, _18289_);
  nor (_18322_, _18311_, _18278_);
  and (_18333_, _18322_, _18267_);
  nor (_18344_, _18333_, _18212_);
  and (_18355_, _18344_, _18092_);
  and (_18366_, _18355_, _17960_);
  or (_18377_, _18366_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  not (_18388_, ABINPUT[0]);
  nand (_18399_, _18366_, _18388_);
  and (_18410_, _18399_, _18377_);
  and (_18421_, _18410_, _16959_);
  not (_18432_, _16948_);
  and (_18443_, _18432_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  not (_18454_, ABINPUT[26]);
  and (_18465_, _18333_, _18212_);
  and (_18476_, _18465_, _18081_);
  and (_18487_, _18476_, _17960_);
  nand (_18498_, _18487_, _18454_);
  not (_18509_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_18520_, _16948_, _18509_);
  or (_18531_, _18487_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_18541_, _18531_, _18520_);
  and (_18552_, _18541_, _18498_);
  or (_18563_, _18552_, _18443_);
  or (_18574_, _18563_, _18421_);
  and (_05301_, _18574_, _27053_);
  not (_18595_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor (_18606_, _18487_, _18595_);
  and (_18617_, _18476_, ABINPUT[0]);
  and (_18628_, _18617_, _17960_);
  or (_18639_, _18628_, _18606_);
  and (_18650_, _18639_, _16959_);
  nor (_18661_, _16948_, _18595_);
  and (_18672_, _18487_, ABINPUT[19]);
  or (_18683_, _18672_, _18606_);
  and (_18694_, _18683_, _18520_);
  or (_18705_, _18694_, _18661_);
  or (_18716_, _18705_, _18650_);
  and (_24640_, _18716_, _27053_);
  not (_18737_, _18212_);
  and (_18748_, _18333_, _18737_);
  and (_18759_, _18748_, _18081_);
  nand (_18770_, _18759_, _17960_);
  and (_18781_, _18770_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_18792_, _18759_, ABINPUT[0]);
  and (_18803_, _18792_, _17960_);
  or (_18814_, _18803_, _18781_);
  and (_18835_, _18814_, _16959_);
  and (_18836_, _18432_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  not (_18847_, ABINPUT[20]);
  nand (_18858_, _18487_, _18847_);
  or (_18869_, _18487_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_18880_, _18869_, _18520_);
  and (_18891_, _18880_, _18858_);
  or (_18902_, _18891_, _18836_);
  or (_18913_, _18902_, _18835_);
  and (_24650_, _18913_, _27053_);
  nor (_18933_, _18333_, _18737_);
  and (_18944_, _18933_, _18081_);
  nand (_18955_, _18944_, _17960_);
  and (_18966_, _18955_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_18977_, _18944_, ABINPUT[0]);
  and (_18988_, _18977_, _17960_);
  or (_18999_, _18988_, _18966_);
  and (_19010_, _18999_, _16959_);
  not (_19021_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nor (_19032_, _16948_, _19021_);
  and (_19043_, _18487_, ABINPUT[21]);
  nor (_19054_, _18487_, _19021_);
  or (_19065_, _19054_, _19043_);
  and (_19076_, _19065_, _18520_);
  or (_19087_, _19076_, _19032_);
  or (_19098_, _19087_, _19010_);
  and (_24660_, _19098_, _27053_);
  and (_19119_, _18344_, _18081_);
  nand (_19130_, _19119_, _17960_);
  and (_19141_, _19130_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_19152_, _19119_, ABINPUT[0]);
  and (_19163_, _19152_, _17960_);
  or (_19174_, _19163_, _19141_);
  and (_19185_, _19174_, _16959_);
  and (_19196_, _18432_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not (_19207_, ABINPUT[22]);
  nand (_19218_, _18487_, _19207_);
  or (_19229_, _18487_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_19240_, _19229_, _18520_);
  and (_19251_, _19240_, _19218_);
  or (_19262_, _19251_, _19196_);
  or (_19273_, _19262_, _19185_);
  and (_24671_, _19273_, _27053_);
  and (_19293_, _18465_, _18092_);
  nand (_19304_, _19293_, _17960_);
  and (_19315_, _19304_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_19337_, _19293_, ABINPUT[0]);
  and (_19338_, _19337_, _17960_);
  or (_19360_, _19338_, _19315_);
  and (_19361_, _19360_, _16959_);
  not (_19383_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor (_19384_, _16948_, _19383_);
  and (_19406_, _18487_, ABINPUT[23]);
  nor (_19407_, _18487_, _19383_);
  or (_19418_, _19407_, _19406_);
  and (_19429_, _19418_, _18520_);
  or (_19440_, _19429_, _19384_);
  or (_19451_, _19440_, _19361_);
  and (_24681_, _19451_, _27053_);
  and (_19472_, _18748_, _18092_);
  nand (_19483_, _19472_, _17960_);
  and (_19494_, _19483_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_19505_, _19472_, ABINPUT[0]);
  and (_19516_, _19505_, _17960_);
  or (_19527_, _19516_, _19494_);
  and (_19538_, _19527_, _16959_);
  and (_19549_, _18432_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_19560_, ABINPUT[24]);
  nand (_19571_, _18487_, _19560_);
  or (_19582_, _18487_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_19593_, _19582_, _18520_);
  and (_19604_, _19593_, _19571_);
  or (_19615_, _19604_, _19549_);
  or (_19626_, _19615_, _19538_);
  and (_24692_, _19626_, _27053_);
  and (_19646_, _18933_, _18092_);
  nand (_19657_, _19646_, _17960_);
  and (_19668_, _19657_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_19679_, _19646_, ABINPUT[0]);
  and (_19690_, _19679_, _17960_);
  or (_19701_, _19690_, _19668_);
  and (_19712_, _19701_, _16959_);
  not (_19723_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor (_19734_, _16948_, _19723_);
  and (_19745_, _18487_, ABINPUT[25]);
  nor (_19756_, _18487_, _19723_);
  or (_19767_, _19756_, _19745_);
  and (_19778_, _19767_, _18520_);
  or (_19789_, _19778_, _19734_);
  or (_19800_, _19789_, _19712_);
  and (_24702_, _19800_, _27053_);
  and (_19821_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_19832_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_19843_, _19832_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_19854_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_19865_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_19876_, _19865_, _19854_);
  and (_19887_, _19832_, _16893_);
  and (_19898_, _19887_, _19876_);
  and (_19909_, _19876_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_19920_, _19909_, _19898_);
  and (_19931_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_19942_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_19953_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_19964_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_19975_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_19986_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_19997_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_20007_, _19997_, _19986_);
  and (_20018_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not (_20029_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_20040_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _20029_);
  and (_20051_, _20040_, _19986_);
  and (_20062_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_20073_, _20062_, _20018_);
  nor (_20084_, _19997_, _19986_);
  and (_20095_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_20106_, _19997_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_20117_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_20128_, _20117_, _20095_);
  and (_20139_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_20150_, _20139_, _19986_);
  and (_20161_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  not (_20172_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_20183_, _20172_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_20194_, _20183_, _19986_);
  and (_20205_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_20216_, _20205_, _20161_);
  and (_20227_, _20216_, _20128_);
  and (_20238_, _20227_, _20073_);
  nor (_20249_, _20238_, _19975_);
  and (_20260_, _20249_, _19964_);
  or (_20271_, _20260_, _19953_);
  and (_20282_, _20271_, _19942_);
  nor (_20293_, _20282_, _19931_);
  and (_20304_, _20293_, _19898_);
  nor (_20315_, _20304_, _19920_);
  not (_20326_, _20315_);
  and (_20337_, _19876_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_20348_, _20337_, _19898_);
  not (_20359_, _19898_);
  and (_20369_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_20380_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_20391_, _20380_, _20369_);
  and (_20402_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  not (_20413_, _20402_);
  and (_20424_, _20413_, _20391_);
  and (_20435_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_20446_, _20435_, _19975_);
  and (_20457_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_20468_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_20479_, _20468_, _20457_);
  and (_20490_, _20479_, _20446_);
  and (_20501_, _20490_, _20424_);
  and (_20512_, _20501_, _19964_);
  nor (_20523_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _19964_);
  or (_20534_, _20523_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_20545_, _20534_, _20512_);
  and (_20556_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_20567_, _20556_, _20545_);
  nor (_20578_, _20567_, _20359_);
  nor (_20589_, _20578_, _20348_);
  not (_20600_, _20589_);
  and (_20611_, _19876_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_20622_, _20611_, _19898_);
  and (_20633_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_20644_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_20655_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_20666_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_20677_, _20666_, _20655_);
  and (_20688_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_20699_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_20710_, _20699_, _20688_);
  and (_20721_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_20731_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_20742_, _20731_, _20721_);
  and (_20753_, _20742_, _20710_);
  and (_20764_, _20753_, _20677_);
  nor (_20775_, _20764_, _19975_);
  and (_20786_, _20775_, _19964_);
  or (_20797_, _20786_, _20644_);
  and (_20808_, _20797_, _19942_);
  nor (_20819_, _20808_, _20633_);
  and (_20830_, _20819_, _19898_);
  nor (_20841_, _20830_, _20622_);
  and (_20852_, _19876_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_20863_, _20852_, _19898_);
  and (_20874_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_20885_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_20896_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_20907_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_20918_, _20907_, _20896_);
  and (_20929_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_20940_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_20951_, _20940_, _20929_);
  and (_20962_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_20973_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_20984_, _20973_, _20962_);
  and (_20995_, _20984_, _20951_);
  and (_21006_, _20995_, _20918_);
  nor (_21017_, _21006_, _19975_);
  and (_21028_, _21017_, _19964_);
  or (_21039_, _21028_, _20885_);
  and (_21050_, _21039_, _19942_);
  nor (_21061_, _21050_, _20874_);
  and (_21071_, _21061_, _19898_);
  nor (_21082_, _21071_, _20863_);
  or (_21093_, _21082_, _20841_);
  nor (_21104_, _21093_, _20600_);
  and (_21115_, _21104_, _20326_);
  and (_21126_, _19876_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_21137_, _21126_, _19898_);
  and (_21148_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_21159_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_21170_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_21181_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_21192_, _21181_, _21170_);
  and (_21203_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_21214_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_21225_, _21214_, _21203_);
  and (_21236_, _21225_, _21192_);
  and (_21247_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_21258_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_21269_, _21258_, _21247_);
  and (_21280_, _21269_, _21236_);
  nor (_21291_, _21280_, _19975_);
  and (_21302_, _21291_, _19964_);
  or (_21313_, _21302_, _21159_);
  and (_21324_, _21313_, _19942_);
  nor (_21335_, _21324_, _21148_);
  and (_21346_, _21335_, _19898_);
  nor (_21357_, _21346_, _21137_);
  and (_21368_, _19876_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_21379_, _21368_, _19898_);
  and (_21390_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_21400_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_21411_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_21422_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_21433_, _21422_, _21411_);
  and (_21444_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_21455_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_21466_, _21455_, _21444_);
  and (_21477_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and (_21488_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_21499_, _21488_, _21477_);
  and (_21510_, _21499_, _21466_);
  and (_21521_, _21510_, _21433_);
  nor (_21532_, _21521_, _19975_);
  and (_21543_, _21532_, _19964_);
  or (_21554_, _21543_, _21400_);
  and (_21565_, _21554_, _19942_);
  nor (_21576_, _21565_, _21390_);
  and (_21587_, _21576_, _19898_);
  nor (_21598_, _21587_, _21379_);
  not (_21609_, _21598_);
  nor (_21620_, _21609_, _21357_);
  and (_21631_, _19876_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_21642_, _21631_, _19898_);
  and (_21653_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_21664_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_21675_, _21664_, _21653_);
  and (_21686_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_21697_, _21686_, _19975_);
  and (_21708_, _21697_, _21675_);
  and (_21718_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  not (_21729_, _21718_);
  and (_21740_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_21751_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_21762_, _21751_, _21740_);
  and (_21773_, _21762_, _21729_);
  and (_21784_, _21773_, _21708_);
  and (_21795_, _21784_, _19964_);
  nor (_21806_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _19964_);
  nor (_21817_, _21806_, _21795_);
  nor (_21828_, _21817_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_21839_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _19942_);
  nor (_21850_, _21839_, _21828_);
  nor (_21861_, _21850_, _20359_);
  nor (_21872_, _21861_, _21642_);
  and (_21883_, _19876_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_21894_, _21883_, _19898_);
  and (_21905_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_21916_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_21927_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_21938_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_21949_, _21938_, _21927_);
  and (_21960_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_21971_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_21982_, _21971_, _21960_);
  and (_21993_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_22004_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_22015_, _22004_, _21993_);
  and (_22025_, _22015_, _21982_);
  and (_22036_, _22025_, _21949_);
  nor (_22047_, _22036_, _19975_);
  and (_22058_, _22047_, _19964_);
  or (_22069_, _22058_, _21916_);
  and (_22080_, _22069_, _19942_);
  nor (_22091_, _22080_, _21905_);
  and (_22102_, _22091_, _19898_);
  nor (_22113_, _22102_, _21894_);
  and (_22124_, _22113_, _21872_);
  and (_22135_, _22124_, _21620_);
  and (_22146_, _22135_, _21115_);
  not (_22157_, _21872_);
  not (_22168_, _22113_);
  and (_22179_, _22168_, _21357_);
  and (_22190_, _22179_, _21598_);
  and (_22201_, _22190_, _22157_);
  and (_22212_, _22201_, _21115_);
  nor (_22223_, _22212_, _22146_);
  not (_22234_, _22223_);
  not (_22245_, _21082_);
  and (_22256_, _22245_, _20841_);
  and (_22267_, _22256_, _20600_);
  nor (_22278_, _21598_, _21357_);
  and (_22289_, _22278_, _22168_);
  and (_22300_, _22289_, _21872_);
  and (_22311_, _22300_, _22267_);
  and (_22322_, _22311_, _20315_);
  nor (_22333_, _22322_, _22234_);
  and (_22343_, _22179_, _21609_);
  and (_22354_, _22343_, _22157_);
  and (_22365_, _22267_, _20315_);
  and (_22376_, _22365_, _22354_);
  and (_22387_, _22113_, _21620_);
  or (_22398_, _20589_, _20315_);
  nor (_22409_, _22398_, _21093_);
  and (_22420_, _22409_, _22387_);
  nor (_22431_, _22420_, _22376_);
  and (_22442_, _22190_, _21872_);
  and (_22453_, _22442_, _22365_);
  and (_22464_, _22113_, _21357_);
  and (_22475_, _22464_, _21609_);
  and (_22486_, _22475_, _21872_);
  and (_22497_, _22486_, _21115_);
  and (_22508_, _22354_, _21104_);
  nor (_22519_, _22508_, _22497_);
  not (_22530_, _22519_);
  nor (_22541_, _22530_, _22453_);
  and (_22552_, _22541_, _22431_);
  and (_22563_, _22552_, _22333_);
  not (_22574_, _22563_);
  and (_22585_, _22168_, _21620_);
  and (_22596_, _22585_, _22157_);
  and (_22607_, _22596_, _21115_);
  and (_22618_, _22343_, _21872_);
  and (_22629_, _22618_, _21104_);
  nor (_22639_, _22629_, _22607_);
  not (_22650_, _22639_);
  not (_22661_, _22365_);
  and (_22672_, _22278_, _22113_);
  nor (_22683_, _22672_, _22618_);
  nor (_22694_, _22683_, _22661_);
  not (_22705_, _22694_);
  and (_22716_, _22585_, _21872_);
  and (_22727_, _22716_, _21115_);
  and (_22738_, _22596_, _22365_);
  nor (_22749_, _22738_, _22727_);
  nand (_22760_, _22749_, _22705_);
  or (_22771_, _22760_, _22650_);
  and (_22782_, _22672_, _21115_);
  and (_22793_, _22157_, _21082_);
  and (_22804_, _22793_, _22387_);
  nor (_22815_, _22804_, _22782_);
  and (_22826_, _22409_, _22190_);
  and (_22837_, _22475_, _22157_);
  and (_22848_, _22837_, _21104_);
  nor (_22859_, _22848_, _22826_);
  nand (_22870_, _22859_, _22815_);
  and (_22881_, _22442_, _21115_);
  and (_22892_, _22113_, _22157_);
  and (_22903_, _22892_, _21620_);
  and (_22914_, _22903_, _21115_);
  nor (_22925_, _22914_, _22881_);
  and (_22936_, _22672_, _22409_);
  and (_22946_, _22936_, _22157_);
  and (_22954_, _22278_, _22124_);
  or (_22961_, _22954_, _22300_);
  and (_22969_, _22961_, _22409_);
  nor (_22977_, _22969_, _22946_);
  nand (_22984_, _22977_, _22925_);
  or (_22992_, _22984_, _22870_);
  and (_23000_, _22837_, _22365_);
  and (_23007_, _22267_, _22201_);
  and (_23010_, _23007_, _20315_);
  or (_23011_, _23010_, _23000_);
  and (_23012_, _21598_, _21357_);
  and (_23019_, _22892_, _23012_);
  and (_23030_, _23019_, _22365_);
  and (_23041_, _22256_, _20589_);
  and (_23052_, _23041_, _22157_);
  and (_23063_, _23052_, _22387_);
  or (_23074_, _23063_, _23030_);
  and (_23085_, _22289_, _22157_);
  and (_23096_, _23085_, _22365_);
  and (_23107_, _21620_, _21872_);
  and (_23118_, _23107_, _22365_);
  or (_23129_, _23118_, _23096_);
  or (_23140_, _23129_, _23074_);
  or (_23151_, _23140_, _23011_);
  or (_23162_, _23151_, _22992_);
  or (_23173_, _23162_, _22771_);
  nor (_23184_, _23173_, _22574_);
  nor (_23195_, _23184_, _19843_);
  not (_23206_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_23216_, \oc8051_top_1.oc8051_decoder1.state [1], _16893_);
  and (_23227_, _23216_, _23206_);
  and (_23237_, _22409_, _22300_);
  or (_23248_, _23237_, _22946_);
  and (_23259_, _23248_, _23227_);
  and (_23270_, _21609_, _21357_);
  and (_23280_, _22409_, _23270_);
  and (_23291_, _23280_, _23227_);
  and (_23302_, _22782_, _23216_);
  and (_23313_, _23302_, \oc8051_top_1.oc8051_decoder1.state [0]);
  or (_23324_, _23313_, _23291_);
  or (_23335_, _23324_, _23259_);
  nor (_23345_, _23335_, _23195_);
  nor (_23356_, _23345_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_23367_, _23356_, _19821_);
  not (_23378_, _23367_);
  and (_23389_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_23400_, _20841_, _20589_);
  and (_23411_, _21872_, _22245_);
  and (_23422_, _23411_, _23400_);
  and (_23433_, _23422_, _22343_);
  and (_23444_, _23041_, _22672_);
  or (_23455_, _23444_, _23433_);
  not (_23466_, _23455_);
  and (_23477_, _22442_, _22409_);
  and (_23488_, _23041_, _22596_);
  nor (_23499_, _23488_, _23477_);
  and (_23510_, _23041_, _22289_);
  and (_23521_, _23041_, _22135_);
  nor (_23532_, _23521_, _23510_);
  not (_23543_, _23532_);
  and (_23554_, _23041_, _22837_);
  nor (_23565_, _23554_, _23543_);
  and (_23576_, _23565_, _23499_);
  and (_23587_, _23576_, _23466_);
  and (_23598_, _21104_, _20315_);
  and (_23609_, _22903_, _23598_);
  and (_23620_, _22716_, _23598_);
  and (_23631_, _23598_, _22486_);
  nor (_23642_, _23631_, _23620_);
  not (_23653_, _23642_);
  nor (_23664_, _23653_, _23609_);
  and (_23675_, _23041_, _22190_);
  and (_23686_, _23041_, _22716_);
  nor (_23697_, _23686_, _23675_);
  and (_23708_, _22464_, _21598_);
  or (_23719_, _23708_, _22343_);
  and (_23730_, _23719_, _23052_);
  nor (_23741_, _23730_, _22782_);
  and (_23752_, _23741_, _23697_);
  and (_23763_, _23752_, _23664_);
  and (_23774_, _23763_, _23587_);
  nor (_23785_, _23774_, _19843_);
  and (_23796_, _23227_, _22475_);
  and (_23807_, _23796_, _22409_);
  or (_23818_, _23807_, _23313_);
  nor (_23829_, _23818_, _23785_);
  nor (_23840_, _23829_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_23851_, _23840_, _23389_);
  and (_23862_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_23873_, _22267_, _20326_);
  and (_23884_, _23873_, _22596_);
  and (_23895_, _23873_, _22903_);
  nor (_23906_, _23895_, _23884_);
  and (_23917_, _23906_, _23664_);
  nor (_23928_, _23917_, _19843_);
  or (_23939_, _23906_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_23950_, _23939_, _19832_);
  nor (_23961_, _23950_, _23291_);
  not (_23972_, _23961_);
  nor (_23983_, _23972_, _23928_);
  nor (_23994_, _23983_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_24005_, _23994_, _23862_);
  nand (_24016_, _24005_, _27053_);
  nor (_03222_, _24016_, _23851_);
  and (_25177_, _03222_, _23378_);
  not (_24047_, _18520_);
  not (_24058_, _17579_);
  nor (_24069_, _24058_, _17307_);
  and (_24080_, _17937_, _17448_);
  and (_24091_, _24080_, _24069_);
  and (_24102_, _24091_, _17742_);
  nand (_24113_, _24102_, _18759_);
  nor (_24124_, _24113_, _24047_);
  and (_24135_, _24124_, ABINPUT[10]);
  nor (_24146_, _24124_, _17013_);
  nor (_24157_, _24146_, _24135_);
  not (_24168_, _24157_);
  not (_24179_, _24124_);
  and (_24190_, _24179_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_24201_, _24124_, ABINPUT[9]);
  nor (_24212_, _24201_, _24190_);
  and (_24223_, _24179_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_24234_, _24124_, ABINPUT[8]);
  nor (_24245_, _24234_, _24223_);
  nor (_24256_, _24124_, _17763_);
  and (_24261_, _24124_, ABINPUT[7]);
  nor (_24262_, _24261_, _24256_);
  and (_24263_, _24179_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_24264_, _24124_, ABINPUT[6]);
  nor (_24265_, _24264_, _24263_);
  and (_24266_, _24179_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_24267_, _24124_, ABINPUT[5]);
  nor (_24268_, _24267_, _24266_);
  and (_24269_, _24179_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_24270_, _24124_, ABINPUT[4]);
  nor (_24271_, _24270_, _24269_);
  nor (_24272_, _24124_, _18157_);
  and (_24273_, _24124_, ABINPUT[3]);
  nor (_24274_, _24273_, _24272_);
  and (_24275_, _24274_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_24276_, _24275_, _24271_);
  and (_24277_, _24276_, _24268_);
  and (_24278_, _24277_, _24265_);
  and (_24279_, _24278_, _24262_);
  and (_24280_, _24279_, _24245_);
  and (_24281_, _24280_, _24212_);
  and (_24282_, _24281_, _24168_);
  nor (_24283_, _24281_, _24168_);
  nor (_24284_, _24283_, _24282_);
  and (_24285_, _24284_, _17002_);
  nor (_24286_, _24285_, _17122_);
  nor (_24287_, _24286_, _24124_);
  nor (_24288_, _24287_, _24135_);
  nor (_25196_, _24288_, rst);
  not (_24289_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_24290_, _24274_, _24289_);
  nor (_24291_, _24274_, _24289_);
  nor (_24292_, _24291_, _24290_);
  and (_24293_, _24292_, _17002_);
  nor (_24294_, _24293_, _18168_);
  nor (_24295_, _24294_, _24124_);
  nor (_24296_, _24295_, _24273_);
  nand (_26240_, _24296_, _27053_);
  nor (_24297_, _24275_, _24271_);
  nor (_24298_, _24297_, _24276_);
  nor (_24299_, _24298_, _16991_);
  nor (_24300_, _24299_, _18256_);
  nor (_24301_, _24300_, _24124_);
  nor (_24302_, _24301_, _24270_);
  nand (_26249_, _24302_, _27053_);
  nor (_24303_, _24276_, _24268_);
  nor (_24304_, _24303_, _24277_);
  nor (_24305_, _24304_, _16991_);
  nor (_24306_, _24305_, _17993_);
  nor (_24307_, _24306_, _24124_);
  nor (_24308_, _24307_, _24267_);
  nand (_26257_, _24308_, _27053_);
  nor (_24309_, _24277_, _24265_);
  nor (_24310_, _24309_, _24278_);
  nor (_24311_, _24310_, _16991_);
  nor (_24312_, _24311_, _17655_);
  nor (_24313_, _24312_, _24124_);
  nor (_24314_, _24313_, _24264_);
  nor (_26266_, _24314_, rst);
  nor (_24315_, _24278_, _24262_);
  nor (_24316_, _24315_, _24279_);
  nor (_24317_, _24316_, _16991_);
  nor (_24318_, _24317_, _17807_);
  nor (_24319_, _24318_, _24124_);
  nor (_24320_, _24319_, _24261_);
  nor (_26274_, _24320_, rst);
  nor (_24321_, _24279_, _24245_);
  nor (_24322_, _24321_, _24280_);
  nor (_24323_, _24322_, _16991_);
  nor (_24324_, _24323_, _17361_);
  nor (_24325_, _24324_, _24124_);
  nor (_24326_, _24325_, _24234_);
  nor (_26283_, _24326_, rst);
  nor (_24327_, _24280_, _24212_);
  nor (_24328_, _24327_, _24281_);
  nor (_24329_, _24328_, _16991_);
  nor (_24330_, _24329_, _17492_);
  nor (_24331_, _24330_, _24124_);
  nor (_24332_, _24331_, _24201_);
  nor (_26291_, _24332_, rst);
  and (_24333_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _16893_);
  and (_24334_, _24333_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_24335_, _18520_, _17742_);
  and (_24336_, _24091_, _19119_);
  and (_24337_, _24336_, _24335_);
  or (_24338_, _24337_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nand (_24339_, _24337_, _18454_);
  and (_24340_, _24339_, _24338_);
  or (_24341_, _24340_, _24334_);
  not (_24342_, ABINPUT[18]);
  nand (_24343_, _24334_, _24342_);
  and (_24344_, _24343_, _27053_);
  and (_28181_, _24344_, _24341_);
  and (_24345_, _18944_, _17742_);
  nand (_24346_, _24345_, _24091_);
  nor (_24347_, _24346_, _24047_);
  nor (_24348_, _24347_, _24334_);
  and (_24349_, _24348_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nor (_24350_, _24348_, _18454_);
  or (_24351_, _24350_, _24349_);
  and (_28202_, _24351_, _27053_);
  and (_24352_, _19119_, _17742_);
  nand (_24353_, _24352_, _24091_);
  nor (_24354_, _24353_, _24047_);
  or (_24355_, _24354_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_24356_, ABINPUT[19]);
  nand (_24357_, _24354_, _24356_);
  and (_24358_, _24357_, _24355_);
  or (_24359_, _24358_, _24334_);
  not (_24360_, ABINPUT[11]);
  nand (_24361_, _24334_, _24360_);
  and (_24362_, _24361_, _27053_);
  and (_29419_, _24362_, _24359_);
  or (_24363_, _24337_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nand (_24364_, _24337_, _18847_);
  and (_24365_, _24364_, _24363_);
  or (_24366_, _24365_, _24334_);
  not (_24367_, ABINPUT[12]);
  nand (_24368_, _24334_, _24367_);
  and (_24369_, _24368_, _27053_);
  and (_29430_, _24369_, _24366_);
  or (_24370_, _24337_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_24371_, ABINPUT[21]);
  nand (_24372_, _24337_, _24371_);
  and (_24373_, _24372_, _24370_);
  or (_24374_, _24373_, _24334_);
  not (_24375_, ABINPUT[13]);
  nand (_24376_, _24334_, _24375_);
  and (_24377_, _24376_, _27053_);
  and (_29441_, _24377_, _24374_);
  or (_24378_, _24337_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nand (_24379_, _24337_, _19207_);
  and (_24380_, _24379_, _24378_);
  or (_24381_, _24380_, _24334_);
  not (_24382_, ABINPUT[14]);
  nand (_24383_, _24334_, _24382_);
  and (_24384_, _24383_, _27053_);
  and (_29452_, _24384_, _24381_);
  or (_24385_, _24354_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_24386_, ABINPUT[23]);
  nand (_24387_, _24354_, _24386_);
  and (_24388_, _24387_, _24385_);
  or (_24389_, _24388_, _24334_);
  not (_24390_, ABINPUT[15]);
  nand (_24391_, _24334_, _24390_);
  and (_24392_, _24391_, _27053_);
  and (_29463_, _24392_, _24389_);
  or (_24393_, _24354_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand (_24394_, _24354_, _19560_);
  and (_24395_, _24394_, _24393_);
  or (_24396_, _24395_, _24334_);
  not (_24397_, ABINPUT[16]);
  nand (_24398_, _24334_, _24397_);
  and (_24399_, _24398_, _27053_);
  and (_29474_, _24399_, _24396_);
  or (_24400_, _24337_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_24401_, ABINPUT[25]);
  nand (_24402_, _24337_, _24401_);
  and (_24403_, _24402_, _24400_);
  or (_24404_, _24403_, _24334_);
  not (_24405_, ABINPUT[17]);
  nand (_24406_, _24334_, _24405_);
  and (_24407_, _24406_, _27053_);
  and (_29485_, _24407_, _24404_);
  and (_24408_, _24348_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nor (_24409_, _24348_, _24356_);
  or (_24410_, _24409_, _24408_);
  and (_29496_, _24410_, _27053_);
  and (_24411_, _24348_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nor (_24412_, _24348_, _18847_);
  or (_24413_, _24412_, _24411_);
  and (_29507_, _24413_, _27053_);
  and (_24414_, _24348_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nor (_24415_, _24348_, _24371_);
  or (_24416_, _24415_, _24414_);
  and (_29518_, _24416_, _27053_);
  and (_24417_, _24348_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nor (_24418_, _24348_, _19207_);
  or (_24419_, _24418_, _24417_);
  and (_29529_, _24419_, _27053_);
  and (_24420_, _24348_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nor (_24421_, _24348_, _24386_);
  or (_24422_, _24421_, _24420_);
  and (_29540_, _24422_, _27053_);
  and (_24423_, _24348_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nor (_24424_, _24348_, _19560_);
  or (_24425_, _24424_, _24423_);
  and (_29551_, _24425_, _27053_);
  and (_24426_, _24348_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nor (_24427_, _24348_, _24401_);
  or (_24428_, _24427_, _24426_);
  and (_29562_, _24428_, _27053_);
  and (_24429_, _17938_, _17448_);
  and (_24430_, _24429_, _24058_);
  not (_24431_, _16959_);
  nor (_24432_, _24431_, _17307_);
  and (_24433_, _24432_, _24430_);
  and (_24434_, _18355_, ABINPUT[0]);
  not (_24435_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_24436_, _18355_, _24435_);
  nor (_24437_, _24436_, _24434_);
  nand (_24438_, _24437_, _24433_);
  nor (_24439_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nor (_24440_, _24439_, _18388_);
  and (_24441_, _24439_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_24442_, _24441_, _24440_);
  or (_24443_, _24442_, _24433_);
  and (_24444_, _24443_, _24438_);
  and (_24445_, _18520_, _18476_);
  and (_24446_, _24445_, _17318_);
  and (_24447_, _24446_, _24430_);
  not (_24448_, _24447_);
  and (_24449_, _24448_, _24444_);
  and (_24450_, _24447_, ABINPUT[10]);
  or (_24451_, _24450_, _24449_);
  and (_01583_, _24451_, _27053_);
  nand (_24452_, _24433_, _18759_);
  and (_24453_, _24452_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_24454_, _24433_, _18792_);
  or (_24455_, _24454_, _24447_);
  or (_24456_, _24455_, _24453_);
  not (_24457_, ABINPUT[4]);
  nand (_24458_, _24447_, _24457_);
  and (_24459_, _24458_, _24456_);
  and (_06362_, _24459_, _27053_);
  not (_24460_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_24461_, _18944_, _24460_);
  nor (_24462_, _24461_, _18977_);
  nand (_24463_, _24462_, _24433_);
  and (_24464_, ABINPUT[2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nor (_24465_, \oc8051_top_1.oc8051_decoder1.psw_set [1], _24460_);
  or (_24466_, _24465_, _24464_);
  or (_24467_, _24466_, _24433_);
  and (_24468_, _24467_, _24463_);
  and (_24469_, _24468_, _24448_);
  and (_24470_, _24447_, ABINPUT[5]);
  or (_24471_, _24470_, _24469_);
  and (_06373_, _24471_, _27053_);
  nor (_24472_, _17579_, _17307_);
  and (_24473_, _24445_, _24429_);
  and (_24474_, _24473_, _24472_);
  not (_24475_, _24474_);
  nand (_24476_, _24433_, _19119_);
  and (_24477_, _24476_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_24478_, _24433_, _19152_);
  or (_24479_, _24478_, _24477_);
  and (_24480_, _24479_, _24475_);
  and (_24481_, _18476_, _17742_);
  not (_24482_, _24481_);
  not (_24483_, _17937_);
  and (_24484_, _24483_, _17448_);
  nand (_24485_, _24484_, _24472_);
  nor (_24486_, _24485_, _24482_);
  and (_24487_, _24486_, _18520_);
  and (_24488_, _24487_, ABINPUT[6]);
  or (_24489_, _24488_, _24480_);
  and (_06384_, _24489_, _27053_);
  nand (_24490_, _24433_, _19293_);
  and (_24491_, _24490_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_24492_, _24433_, _19337_);
  or (_24493_, _24492_, _24491_);
  and (_24494_, _24493_, _24475_);
  and (_24495_, _24487_, ABINPUT[7]);
  or (_24496_, _24495_, _24494_);
  and (_06394_, _24496_, _27053_);
  nand (_24497_, _24433_, _19472_);
  and (_24498_, _24497_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_24499_, _24433_, _19505_);
  or (_24500_, _24499_, _24447_);
  or (_24501_, _24500_, _24498_);
  not (_24502_, ABINPUT[8]);
  nand (_24503_, _24447_, _24502_);
  and (_24504_, _24503_, _24501_);
  and (_06405_, _24504_, _27053_);
  not (_24505_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_24506_, _19646_, _24505_);
  nor (_24507_, _24506_, _19679_);
  nand (_24508_, _24507_, _24433_);
  and (_24509_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_24510_, _24509_, ABINPUT[1]);
  nor (_24511_, _24509_, _24505_);
  or (_24512_, _24511_, _24510_);
  or (_24513_, _24512_, _24433_);
  and (_24514_, _24513_, _24508_);
  and (_24515_, _24514_, _24448_);
  and (_24516_, _24447_, ABINPUT[9]);
  or (_24517_, _24516_, _24515_);
  and (_06416_, _24517_, _27053_);
  not (_24518_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_24519_, _24333_, _24518_);
  and (_24520_, _24519_, ABINPUT[18]);
  nor (_24521_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_24522_, _24521_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not (_24523_, _17448_);
  and (_24524_, _17937_, _24523_);
  nand (_24525_, _24524_, _24472_);
  nor (_24526_, _24525_, _24482_);
  and (_24527_, _24526_, _18520_);
  nor (_24528_, _24527_, _24522_);
  not (_24529_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_24530_, _17937_, _17742_);
  and (_24531_, _24530_, _17589_);
  and (_24532_, _24531_, _24432_);
  and (_24533_, _24532_, _18355_);
  nor (_24534_, _24533_, _24529_);
  and (_24535_, _24532_, _24434_);
  nor (_24536_, _24535_, _24534_);
  and (_24537_, _24536_, _24528_);
  nor (_24538_, _24528_, ABINPUT[26]);
  or (_24539_, _24538_, _24537_);
  nor (_24540_, _24539_, _24519_);
  nor (_24541_, _24540_, _24520_);
  nor (_07125_, _24541_, rst);
  and (_24542_, _24519_, ABINPUT[11]);
  not (_24543_, _24519_);
  nor (_24544_, _24528_, _24356_);
  and (_24545_, _24530_, _17318_);
  and (_24546_, _16959_, _17589_);
  and (_24547_, _24546_, _24545_);
  or (_24548_, _24519_, _18476_);
  nand (_24549_, _24548_, _24547_);
  and (_24550_, _24549_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_24551_, _24547_, _18617_);
  or (_24552_, _24551_, _24550_);
  and (_24553_, _24552_, _24528_);
  or (_24554_, _24553_, _24544_);
  and (_24555_, _24554_, _24543_);
  nor (_24556_, _24555_, _24542_);
  nor (_08829_, _24556_, rst);
  and (_24557_, _24528_, _24543_);
  not (_24558_, _24557_);
  nand (_24559_, _24547_, _18759_);
  and (_24560_, _24559_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_24561_, _24532_, _18792_);
  nor (_24562_, _24561_, _24560_);
  nor (_24563_, _24562_, _24558_);
  not (_24564_, _24563_);
  and (_24565_, _24519_, ABINPUT[12]);
  or (_24566_, _24519_, _18847_);
  nor (_24567_, _24566_, _24528_);
  nor (_24568_, _24567_, _24565_);
  and (_24569_, _24568_, _24564_);
  nor (_08840_, _24569_, rst);
  and (_24570_, _24519_, ABINPUT[13]);
  not (_24571_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_24572_, _24532_, _18944_);
  nor (_24573_, _24572_, _24571_);
  and (_24574_, _24532_, _18977_);
  nor (_24575_, _24574_, _24573_);
  nor (_24576_, _24575_, _24558_);
  nor (_24577_, _24528_, _24371_);
  or (_24578_, _24577_, _24576_);
  and (_24579_, _24578_, _24543_);
  nor (_24580_, _24579_, _24570_);
  nor (_08851_, _24580_, rst);
  and (_24581_, _24519_, ABINPUT[14]);
  nor (_24582_, _24528_, _19207_);
  not (_24583_, _24528_);
  nand (_24584_, _24547_, _19119_);
  and (_24585_, _24584_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_24586_, _24547_, _19152_);
  nor (_24587_, _24586_, _24585_);
  nor (_24588_, _24587_, _24583_);
  nor (_24589_, _24588_, _24582_);
  nor (_24590_, _24589_, _24519_);
  nor (_24591_, _24590_, _24581_);
  nor (_08862_, _24591_, rst);
  not (_24592_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_24593_, _24532_, _19293_);
  nor (_24594_, _24593_, _24592_);
  and (_24595_, _24532_, _19337_);
  nor (_24596_, _24595_, _24594_);
  nor (_24597_, _24596_, _24558_);
  not (_24598_, _24597_);
  and (_24599_, _24519_, ABINPUT[15]);
  or (_24600_, _24519_, _24386_);
  nor (_24601_, _24600_, _24528_);
  nor (_24602_, _24601_, _24599_);
  and (_24603_, _24602_, _24598_);
  nor (_08873_, _24603_, rst);
  and (_24604_, _24519_, ABINPUT[16]);
  nor (_24605_, _24528_, _19560_);
  nand (_24606_, _24547_, _19472_);
  and (_24607_, _24606_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_24608_, _24532_, _19505_);
  nor (_24609_, _24608_, _24607_);
  nor (_24610_, _24609_, _24583_);
  nor (_24611_, _24610_, _24605_);
  nor (_24612_, _24611_, _24519_);
  nor (_24613_, _24612_, _24604_);
  nor (_08884_, _24613_, rst);
  not (_24614_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_24615_, _24532_, _19646_);
  nor (_24616_, _24615_, _24614_);
  and (_24617_, _24532_, _19679_);
  nor (_24618_, _24617_, _24616_);
  nor (_24619_, _24618_, _24558_);
  not (_24620_, _24619_);
  and (_24621_, _24519_, ABINPUT[17]);
  or (_24622_, _24519_, _24401_);
  nor (_24623_, _24622_, _24528_);
  nor (_24624_, _24623_, _24621_);
  and (_24625_, _24624_, _24620_);
  nor (_08895_, _24625_, rst);
  and (_24626_, _24102_, _18355_);
  or (_24627_, _24626_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nand (_24628_, _24626_, _18388_);
  and (_24629_, _24628_, _16959_);
  and (_24630_, _24629_, _24627_);
  not (_24631_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_24632_, _24091_, _24481_);
  nor (_24633_, _24632_, _24631_);
  and (_24634_, _24632_, ABINPUT[10]);
  or (_24635_, _24634_, _24633_);
  and (_24636_, _24635_, _18520_);
  nor (_24637_, _16948_, _24631_);
  or (_24638_, _24637_, rst);
  or (_24639_, _24638_, _24636_);
  or (_19326_, _24639_, _24630_);
  and (_24641_, _24429_, _24069_);
  and (_24642_, _24641_, _18476_);
  and (_24643_, _24642_, ABINPUT[10]);
  not (_24644_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_24645_, _24642_, _24644_);
  or (_24646_, _24645_, _24643_);
  and (_24647_, _24646_, _18520_);
  nor (_24648_, _18355_, _24644_);
  or (_24649_, _24648_, _24434_);
  and (_24651_, _24649_, _24641_);
  nor (_24652_, _24641_, _24644_);
  or (_24653_, _24652_, _24651_);
  and (_24654_, _24653_, _16959_);
  nor (_24655_, _16948_, _24644_);
  or (_24656_, _24655_, rst);
  or (_24657_, _24656_, _24654_);
  or (_19349_, _24657_, _24647_);
  and (_24658_, _24524_, _24069_);
  and (_24659_, _24658_, _24481_);
  and (_24661_, _24659_, ABINPUT[10]);
  not (_24662_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_24663_, _24659_, _24662_);
  or (_24664_, _24663_, _24661_);
  and (_24665_, _24664_, _18520_);
  and (_24666_, _17579_, _24523_);
  and (_24667_, _24666_, _24545_);
  nor (_24668_, _18355_, _24662_);
  or (_24669_, _24668_, _24434_);
  and (_24670_, _24669_, _24667_);
  nor (_24672_, _24667_, _24662_);
  or (_24673_, _24672_, _24670_);
  and (_24674_, _24673_, _16959_);
  nor (_24675_, _16948_, _24662_);
  or (_24676_, _24675_, rst);
  or (_24677_, _24676_, _24674_);
  or (_19372_, _24677_, _24665_);
  not (_24678_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_24679_, _17937_, _17448_);
  and (_24680_, _24069_, _24679_);
  and (_24682_, _24680_, _24481_);
  nor (_24683_, _24682_, _24678_);
  and (_24684_, _24682_, ABINPUT[10]);
  or (_24685_, _24684_, _24683_);
  and (_24686_, _24685_, _18520_);
  and (_24687_, _24666_, _17318_);
  and (_24688_, _24687_, _17938_);
  nor (_24689_, _24688_, _24678_);
  nor (_24690_, _18355_, _24678_);
  or (_24691_, _24690_, _24434_);
  and (_24693_, _24691_, _24688_);
  or (_24694_, _24693_, _24689_);
  and (_24695_, _24694_, _16959_);
  nor (_24696_, _16948_, _24678_);
  or (_24697_, _24696_, rst);
  or (_24698_, _24697_, _24695_);
  or (_19395_, _24698_, _24686_);
  not (_24699_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_24700_, _24632_, _24699_);
  and (_24701_, _24102_, _18617_);
  or (_24703_, _24701_, _24700_);
  and (_24704_, _24703_, _16959_);
  and (_24705_, _24632_, ABINPUT[3]);
  or (_24706_, _24705_, _24700_);
  and (_24707_, _24706_, _18520_);
  nor (_24708_, _16948_, _24699_);
  or (_24709_, _24708_, rst);
  or (_24710_, _24709_, _24707_);
  or (_26462_, _24710_, _24704_);
  and (_24711_, _24113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_24712_, _24102_, _18792_);
  or (_24713_, _24712_, _24711_);
  and (_24714_, _24713_, _16959_);
  not (_24715_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_24716_, _24632_, _24715_);
  and (_24717_, _24632_, ABINPUT[4]);
  or (_24718_, _24717_, _24716_);
  and (_24719_, _24718_, _18520_);
  nor (_24720_, _16948_, _24715_);
  or (_24721_, _24720_, _24719_);
  or (_24722_, _24721_, _24714_);
  or (_26464_, _24722_, rst);
  not (_24723_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_24724_, _24632_, _24723_);
  and (_24725_, _24632_, ABINPUT[5]);
  or (_24726_, _24725_, _24724_);
  and (_24727_, _24726_, _18520_);
  and (_24728_, _24346_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_24729_, _24102_, _18977_);
  or (_24730_, _24729_, _24728_);
  and (_24731_, _24730_, _16959_);
  nor (_24732_, _16948_, _24723_);
  or (_24733_, _24732_, rst);
  or (_24734_, _24733_, _24731_);
  or (_26466_, _24734_, _24727_);
  not (_24735_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_24736_, _24632_, _24735_);
  and (_24737_, _24632_, ABINPUT[6]);
  or (_24738_, _24737_, _24736_);
  and (_24739_, _24738_, _18520_);
  and (_24740_, _24353_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_24741_, _24102_, _19152_);
  or (_24742_, _24741_, _24740_);
  and (_24743_, _24742_, _16959_);
  nor (_24744_, _16948_, _24735_);
  or (_24745_, _24744_, rst);
  or (_24746_, _24745_, _24743_);
  or (_26468_, _24746_, _24739_);
  and (_24747_, _24102_, _19293_);
  or (_24748_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand (_24749_, _24747_, _18388_);
  and (_24750_, _24749_, _16959_);
  and (_24751_, _24750_, _24748_);
  not (_24752_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_24753_, _24632_, _24752_);
  and (_24754_, _24632_, ABINPUT[7]);
  or (_24755_, _24754_, _24753_);
  and (_24756_, _24755_, _18520_);
  nor (_24757_, _16948_, _24752_);
  or (_24758_, _24757_, rst);
  or (_24759_, _24758_, _24756_);
  or (_26469_, _24759_, _24751_);
  nand (_24760_, _24102_, _19472_);
  and (_24761_, _24760_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_24762_, _24102_, _19505_);
  or (_24763_, _24762_, _24761_);
  and (_24764_, _24763_, _16959_);
  not (_24765_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_24766_, _24632_, _24765_);
  and (_24767_, _24632_, ABINPUT[8]);
  or (_24768_, _24767_, _24766_);
  and (_24769_, _24768_, _18520_);
  nor (_24770_, _16948_, _24765_);
  or (_24771_, _24770_, rst);
  or (_24772_, _24771_, _24769_);
  or (_26471_, _24772_, _24764_);
  nand (_24773_, _24102_, _19646_);
  and (_24774_, _24773_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_24775_, _24102_, _19679_);
  or (_24776_, _24775_, _24774_);
  and (_24777_, _24776_, _16959_);
  not (_24778_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_24779_, _24632_, _24778_);
  and (_24780_, _24632_, ABINPUT[9]);
  or (_24781_, _24780_, _24779_);
  and (_24782_, _24781_, _18520_);
  nor (_24783_, _16948_, _24778_);
  or (_24784_, _24783_, rst);
  or (_24785_, _24784_, _24782_);
  or (_26473_, _24785_, _24777_);
  not (_24786_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_24787_, _24642_, _24786_);
  and (_24788_, _24642_, ABINPUT[3]);
  or (_24789_, _24788_, _24787_);
  and (_24790_, _24789_, _18520_);
  or (_24791_, _24787_, _18617_);
  or (_24792_, _24641_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_24793_, _24792_, _16959_);
  and (_24794_, _24793_, _24791_);
  nor (_24795_, _16948_, _24786_);
  or (_24796_, _24795_, rst);
  or (_24797_, _24796_, _24794_);
  or (_26474_, _24797_, _24790_);
  and (_24798_, _24642_, ABINPUT[4]);
  not (_24799_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_24800_, _24642_, _24799_);
  or (_24801_, _24800_, _24798_);
  and (_24802_, _24801_, _18520_);
  nor (_24803_, _18759_, _24799_);
  or (_24804_, _24803_, _18792_);
  and (_24805_, _24804_, _24641_);
  nor (_24806_, _24641_, _24799_);
  or (_24807_, _24806_, _24805_);
  and (_24808_, _24807_, _16959_);
  nor (_24809_, _16948_, _24799_);
  or (_24810_, _24809_, rst);
  or (_24811_, _24810_, _24808_);
  or (_26476_, _24811_, _24802_);
  and (_24812_, _24642_, ABINPUT[5]);
  not (_24813_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_24814_, _24642_, _24813_);
  or (_24815_, _24814_, _24812_);
  and (_24816_, _24815_, _18520_);
  nor (_24817_, _18944_, _24813_);
  or (_24818_, _24817_, _18977_);
  and (_24819_, _24818_, _24641_);
  nor (_24820_, _24641_, _24813_);
  or (_24821_, _24820_, _24819_);
  and (_24822_, _24821_, _16959_);
  nor (_24823_, _16948_, _24813_);
  or (_24824_, _24823_, rst);
  or (_24825_, _24824_, _24822_);
  or (_26478_, _24825_, _24816_);
  and (_24826_, _24642_, ABINPUT[6]);
  not (_24827_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_24828_, _24642_, _24827_);
  or (_24829_, _24828_, _24826_);
  and (_24830_, _24829_, _18520_);
  nor (_24831_, _19119_, _24827_);
  or (_24832_, _24831_, _19152_);
  and (_24833_, _24832_, _24641_);
  nor (_24834_, _24641_, _24827_);
  or (_24835_, _24834_, _24833_);
  and (_24836_, _24835_, _16959_);
  nor (_24837_, _16948_, _24827_);
  or (_24838_, _24837_, rst);
  or (_24839_, _24838_, _24836_);
  or (_26480_, _24839_, _24830_);
  and (_24840_, _24642_, ABINPUT[7]);
  not (_24841_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nor (_24842_, _24642_, _24841_);
  or (_24843_, _24842_, _24840_);
  and (_24844_, _24843_, _18520_);
  nor (_24845_, _19293_, _24841_);
  or (_24846_, _24845_, _19337_);
  and (_24847_, _24846_, _24641_);
  nor (_24848_, _24641_, _24841_);
  or (_24849_, _24848_, _24847_);
  and (_24850_, _24849_, _16959_);
  nor (_24851_, _16948_, _24841_);
  or (_24852_, _24851_, rst);
  or (_24853_, _24852_, _24850_);
  or (_26482_, _24853_, _24844_);
  and (_24854_, _24642_, ABINPUT[8]);
  not (_24855_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_24856_, _24642_, _24855_);
  or (_24857_, _24856_, _24854_);
  and (_24858_, _24857_, _18520_);
  nor (_24859_, _19472_, _24855_);
  or (_24860_, _24859_, _19505_);
  and (_24861_, _24860_, _24641_);
  nor (_24862_, _24641_, _24855_);
  or (_24863_, _24862_, _24861_);
  and (_24864_, _24863_, _16959_);
  nor (_24865_, _16948_, _24855_);
  or (_24866_, _24865_, rst);
  or (_24867_, _24866_, _24864_);
  or (_26483_, _24867_, _24858_);
  and (_24868_, _24642_, ABINPUT[9]);
  not (_24869_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_24870_, _24642_, _24869_);
  or (_24871_, _24870_, _24868_);
  and (_24872_, _24871_, _18520_);
  nor (_24873_, _19646_, _24869_);
  or (_24874_, _24873_, _19679_);
  and (_24875_, _24874_, _24641_);
  nor (_24876_, _24641_, _24869_);
  or (_24877_, _24876_, _24875_);
  and (_24878_, _24877_, _16959_);
  nor (_24879_, _16948_, _24869_);
  or (_24880_, _24879_, rst);
  or (_24881_, _24880_, _24878_);
  or (_26485_, _24881_, _24872_);
  and (_24882_, _24659_, ABINPUT[3]);
  not (_24883_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_24884_, _24659_, _24883_);
  or (_24885_, _24884_, _24882_);
  and (_24886_, _24885_, _18520_);
  nor (_24887_, _18476_, _24883_);
  or (_24888_, _24887_, _18617_);
  and (_24889_, _24888_, _24667_);
  nor (_24890_, _24667_, _24883_);
  or (_24891_, _24890_, _24889_);
  and (_24892_, _24891_, _16959_);
  nor (_24893_, _16948_, _24883_);
  or (_24894_, _24893_, rst);
  or (_24895_, _24894_, _24892_);
  or (_26487_, _24895_, _24886_);
  and (_24896_, _24659_, ABINPUT[4]);
  not (_24897_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_24898_, _24659_, _24897_);
  or (_24899_, _24898_, _24896_);
  and (_24900_, _24899_, _18520_);
  nor (_24901_, _18759_, _24897_);
  or (_24902_, _24901_, _18792_);
  and (_24903_, _24902_, _24667_);
  nor (_24904_, _24667_, _24897_);
  or (_24905_, _24904_, _24903_);
  and (_24906_, _24905_, _16959_);
  nor (_24907_, _16948_, _24897_);
  or (_24908_, _24907_, rst);
  or (_24909_, _24908_, _24906_);
  or (_26489_, _24909_, _24900_);
  and (_24910_, _24659_, ABINPUT[5]);
  not (_24911_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_24912_, _24659_, _24911_);
  or (_24913_, _24912_, _24910_);
  and (_24914_, _24913_, _18520_);
  nor (_24915_, _18944_, _24911_);
  or (_24916_, _24915_, _18977_);
  and (_24917_, _24916_, _24667_);
  nor (_24918_, _24667_, _24911_);
  or (_24919_, _24918_, _24917_);
  and (_24920_, _24919_, _16959_);
  nor (_24921_, _16948_, _24911_);
  or (_24922_, _24921_, rst);
  or (_24923_, _24922_, _24920_);
  or (_26490_, _24923_, _24914_);
  and (_24924_, _24659_, ABINPUT[6]);
  not (_24925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor (_24926_, _24659_, _24925_);
  or (_24927_, _24926_, _24924_);
  and (_24928_, _24927_, _18520_);
  nor (_24929_, _19119_, _24925_);
  or (_24930_, _24929_, _19152_);
  and (_24931_, _24930_, _24667_);
  nor (_24932_, _24667_, _24925_);
  or (_24933_, _24932_, _24931_);
  and (_24934_, _24933_, _16959_);
  nor (_24935_, _16948_, _24925_);
  or (_24936_, _24935_, rst);
  or (_24937_, _24936_, _24934_);
  or (_26492_, _24937_, _24928_);
  not (_24938_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor (_24939_, _19293_, _24938_);
  or (_24940_, _24939_, _19337_);
  and (_24941_, _24940_, _24667_);
  nor (_24942_, _24667_, _24938_);
  or (_24943_, _24942_, _24941_);
  and (_24944_, _24943_, _16959_);
  and (_24945_, _24659_, ABINPUT[7]);
  nor (_24946_, _24659_, _24938_);
  or (_24947_, _24946_, _24945_);
  and (_24948_, _24947_, _18520_);
  nor (_24949_, _16948_, _24938_);
  or (_24950_, _24949_, rst);
  or (_24951_, _24950_, _24948_);
  or (_26494_, _24951_, _24944_);
  not (_24952_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor (_24953_, _19472_, _24952_);
  or (_24954_, _24953_, _19505_);
  and (_24955_, _24954_, _24667_);
  nor (_24956_, _24667_, _24952_);
  or (_24957_, _24956_, _24955_);
  and (_24958_, _24957_, _16959_);
  and (_24959_, _24659_, ABINPUT[8]);
  nor (_24960_, _24659_, _24952_);
  or (_24961_, _24960_, _24959_);
  and (_24962_, _24961_, _18520_);
  nor (_24963_, _16948_, _24952_);
  or (_24964_, _24963_, rst);
  or (_24965_, _24964_, _24962_);
  or (_26496_, _24965_, _24958_);
  not (_24966_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_24967_, _19646_, _24966_);
  or (_24968_, _24967_, _19679_);
  and (_24969_, _24968_, _24667_);
  nor (_24970_, _24667_, _24966_);
  or (_24971_, _24970_, _24969_);
  and (_24972_, _24971_, _16959_);
  and (_24973_, _24659_, ABINPUT[9]);
  nor (_24974_, _24659_, _24966_);
  or (_24975_, _24974_, _24973_);
  and (_24976_, _24975_, _18520_);
  nor (_24977_, _16948_, _24966_);
  or (_24978_, _24977_, rst);
  or (_24979_, _24978_, _24976_);
  or (_26497_, _24979_, _24972_);
  and (_24980_, _24682_, ABINPUT[3]);
  not (_24981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_24982_, _24682_, _24981_);
  or (_24983_, _24982_, _24980_);
  and (_24984_, _24983_, _18520_);
  nor (_24985_, _24688_, _24981_);
  nor (_24986_, _18476_, _24981_);
  or (_24987_, _24986_, _18617_);
  and (_24988_, _24987_, _24688_);
  or (_24989_, _24988_, _24985_);
  and (_24990_, _24989_, _16959_);
  nor (_24991_, _16948_, _24981_);
  or (_24992_, _24991_, rst);
  or (_24993_, _24992_, _24990_);
  or (_26499_, _24993_, _24984_);
  not (_24994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_24995_, _24682_, _24994_);
  and (_24996_, _24682_, ABINPUT[4]);
  or (_24997_, _24996_, _24995_);
  and (_24998_, _24997_, _18520_);
  nor (_24999_, _24688_, _24994_);
  nor (_25000_, _18759_, _24994_);
  or (_25001_, _25000_, _18792_);
  and (_25002_, _25001_, _24688_);
  or (_25003_, _25002_, _24999_);
  and (_25004_, _25003_, _16959_);
  nor (_25005_, _16948_, _24994_);
  or (_25006_, _25005_, rst);
  or (_25007_, _25006_, _25004_);
  or (_26501_, _25007_, _24998_);
  not (_25008_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_25009_, _24682_, _25008_);
  and (_25010_, _24682_, ABINPUT[5]);
  or (_25011_, _25010_, _25009_);
  and (_25012_, _25011_, _18520_);
  nor (_25013_, _24688_, _25008_);
  nor (_25014_, _18944_, _25008_);
  or (_25015_, _25014_, _18977_);
  and (_25016_, _25015_, _24688_);
  or (_25017_, _25016_, _25013_);
  and (_25018_, _25017_, _16959_);
  nor (_25019_, _16948_, _25008_);
  or (_25020_, _25019_, rst);
  or (_25021_, _25020_, _25018_);
  or (_26503_, _25021_, _25012_);
  not (_25022_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_25023_, _24682_, _25022_);
  and (_25024_, _24682_, ABINPUT[6]);
  or (_25025_, _25024_, _25023_);
  and (_25026_, _25025_, _18520_);
  nor (_25027_, _24688_, _25022_);
  nor (_25028_, _19119_, _25022_);
  or (_25029_, _25028_, _19152_);
  and (_25030_, _25029_, _24688_);
  or (_25031_, _25030_, _25027_);
  and (_25032_, _25031_, _16959_);
  nor (_25033_, _16948_, _25022_);
  or (_25034_, _25033_, rst);
  or (_25035_, _25034_, _25032_);
  or (_26504_, _25035_, _25026_);
  not (_25036_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor (_25037_, _24682_, _25036_);
  and (_25038_, _24682_, ABINPUT[7]);
  or (_25039_, _25038_, _25037_);
  and (_25040_, _25039_, _18520_);
  nor (_25041_, _24688_, _25036_);
  nor (_25042_, _19293_, _25036_);
  or (_25043_, _25042_, _19337_);
  and (_25044_, _25043_, _24688_);
  or (_25045_, _25044_, _25041_);
  and (_25046_, _25045_, _16959_);
  nor (_25047_, _16948_, _25036_);
  or (_25048_, _25047_, rst);
  or (_25049_, _25048_, _25046_);
  or (_26506_, _25049_, _25040_);
  not (_25050_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor (_25051_, _24682_, _25050_);
  and (_25052_, _24682_, ABINPUT[8]);
  or (_25053_, _25052_, _25051_);
  and (_25054_, _25053_, _18520_);
  nor (_25055_, _24688_, _25050_);
  nor (_25056_, _19472_, _25050_);
  or (_25057_, _25056_, _19505_);
  and (_25058_, _25057_, _24688_);
  or (_25059_, _25058_, _25055_);
  and (_25060_, _25059_, _16959_);
  nor (_25061_, _16948_, _25050_);
  or (_25062_, _25061_, rst);
  or (_25063_, _25062_, _25060_);
  or (_26508_, _25063_, _25054_);
  not (_25064_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_25065_, _24682_, _25064_);
  and (_25066_, _24682_, ABINPUT[9]);
  or (_25067_, _25066_, _25065_);
  and (_25068_, _25067_, _18520_);
  nor (_25069_, _24688_, _25064_);
  nor (_25070_, _19646_, _25064_);
  or (_25071_, _25070_, _19679_);
  and (_25072_, _25071_, _24688_);
  or (_25073_, _25072_, _25069_);
  and (_25074_, _25073_, _16959_);
  nor (_25075_, _16948_, _25064_);
  or (_25076_, _25075_, rst);
  or (_25077_, _25076_, _25074_);
  or (_26510_, _25077_, _25068_);
  and (_25078_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_25079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _27053_);
  and (_27056_, _25079_, _25078_);
  and (_25080_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_25081_, _25080_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_25082_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_25083_, _25082_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor (_25084_, _25083_, _25081_);
  not (_25085_, _25084_);
  and (_25086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_25087_, _25086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_25088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_25089_, _25088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_25090_, _25089_, _25087_);
  nor (_25091_, _25090_, _25085_);
  not (_25092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_25093_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_25094_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_25095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_25096_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _25095_);
  or (_25097_, _25096_, _25094_);
  nor (_25098_, _25097_, _25093_);
  nor (_25099_, _25098_, _25092_);
  nor (_25100_, _25099_, _25091_);
  not (_25101_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_25102_, _25080_, _25101_);
  not (_25103_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_25104_, _25082_, _25103_);
  nor (_25105_, _25104_, _25102_);
  not (_25106_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_25107_, _25086_, _25106_);
  not (_25108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_25109_, _25088_, _25108_);
  nor (_25110_, _25109_, _25107_);
  and (_25111_, _25110_, _25105_);
  nor (_25112_, _25111_, _25093_);
  and (_25113_, _25112_, _25092_);
  nor (_25114_, _25113_, _25100_);
  and (_25115_, _25114_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_25116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _25095_);
  and (_25117_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _25095_);
  nor (_25118_, _25117_, _25116_);
  not (_25119_, _25118_);
  and (_25120_, _25119_, _25100_);
  or (_25121_, _25120_, _25078_);
  or (_25122_, _25121_, _25115_);
  not (_25123_, _25078_);
  or (_25124_, _25118_, _25123_);
  and (_25125_, _25124_, _27053_);
  and (_27058_, _25125_, _25122_);
  nand (_25126_, _25091_, _25092_);
  or (_25127_, _25126_, _25112_);
  nand (_25128_, _25116_, _25078_);
  and (_25129_, _25128_, _27053_);
  and (_27061_, _25129_, _25127_);
  and (_25130_, _25114_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  not (_25131_, _25089_);
  and (_25132_, _25131_, _25084_);
  and (_25133_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25134_, _25133_, _25132_);
  and (_25135_, _25087_, _25095_);
  or (_25136_, _25085_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_25137_, _25136_, _25135_);
  and (_25138_, _25137_, _25134_);
  and (_25139_, _25138_, _25100_);
  or (_25140_, _25139_, _25130_);
  and (_25141_, _25113_, _25091_);
  and (_25142_, _25107_, _25095_);
  or (_25143_, _25142_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  not (_25144_, _25105_);
  and (_25145_, _25109_, _25095_);
  nor (_25146_, _25145_, _25144_);
  and (_25147_, _25146_, _25143_);
  and (_25148_, _25133_, _25144_);
  or (_25149_, _25148_, _25147_);
  and (_25150_, _25149_, _25141_);
  or (_25151_, _25150_, _25078_);
  or (_25152_, _25151_, _25140_);
  or (_25153_, _25123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_25154_, _25153_, _27053_);
  and (_27064_, _25154_, _25152_);
  and (_25155_, _25114_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_25156_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _25095_);
  or (_25157_, _25156_, _25132_);
  and (_25158_, _25087_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25159_, _25085_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_25160_, _25159_, _25158_);
  and (_25161_, _25160_, _25157_);
  and (_25162_, _25161_, _25100_);
  or (_25163_, _25162_, _25155_);
  and (_25164_, _25107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25165_, _25164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_25166_, _25109_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_25167_, _25166_, _25144_);
  and (_25168_, _25167_, _25165_);
  and (_25169_, _25156_, _25144_);
  or (_25170_, _25169_, _25168_);
  and (_25171_, _25170_, _25141_);
  or (_25172_, _25171_, _25078_);
  or (_25173_, _25172_, _25163_);
  or (_25174_, _25123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_25175_, _25174_, _27053_);
  and (_27066_, _25175_, _25173_);
  nor (_25176_, _25078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_25178_, _25176_, _25100_);
  nand (_25179_, _25113_, _25095_);
  and (_25180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _27053_);
  nand (_25181_, _25180_, _25179_);
  nor (_27068_, _25181_, _25178_);
  nor (_25182_, _25078_, _25095_);
  and (_25183_, _25182_, _25100_);
  nand (_25184_, _25113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_25185_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _27053_);
  nand (_25186_, _25185_, _25184_);
  nor (_27070_, _25186_, _25183_);
  nor (_25187_, _24431_, _17742_);
  and (_25188_, _25187_, _24091_);
  and (_25189_, _25188_, _19119_);
  nand (_25190_, _25189_, _18388_);
  and (_25191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_25192_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _25095_);
  and (_25193_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_25194_, _25193_, _25192_);
  nor (_25195_, _25194_, _25092_);
  nand (_25197_, _25195_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and (_25198_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _25095_);
  and (_25199_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_25200_, _25199_, _25198_);
  nor (_25201_, _25200_, _25092_);
  nor (_25202_, _25156_, _25133_);
  nand (_25203_, _25202_, _25201_);
  or (_25204_, _25203_, _25197_);
  and (_25205_, _25204_, _25191_);
  or (_25206_, _25205_, _25189_);
  and (_25207_, _25206_, _25190_);
  and (_25208_, _24445_, _17753_);
  and (_25209_, _25208_, _24091_);
  or (_25210_, _25209_, _25207_);
  not (_25211_, ABINPUT[6]);
  nand (_25212_, _25209_, _25211_);
  and (_25213_, _25212_, _27053_);
  and (_27105_, _25213_, _25210_);
  and (_25214_, _25188_, _18759_);
  nand (_25215_, _25214_, _18388_);
  not (_25216_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_25217_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _25216_);
  nor (_25218_, _25202_, _25092_);
  or (_25219_, _25218_, _25201_);
  or (_25220_, _25219_, _25197_);
  and (_25221_, _25220_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_25222_, _25221_, _25217_);
  or (_25223_, _25222_, _25214_);
  and (_25224_, _25223_, _25215_);
  or (_25225_, _25224_, _25209_);
  nand (_25226_, _25209_, _24457_);
  and (_25227_, _25226_, _27053_);
  and (_27107_, _25227_, _25225_);
  not (_25228_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_25229_, _25195_, _25228_);
  or (_25230_, _25229_, _25203_);
  nand (_25231_, _25230_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_25232_, _25188_, _19472_);
  nor (_25233_, _25232_, _25231_);
  and (_25234_, _25232_, ABINPUT[0]);
  or (_25235_, _25234_, _25209_);
  or (_25236_, _25235_, _25233_);
  nand (_25237_, _25209_, _24502_);
  and (_25238_, _25237_, _27053_);
  and (_27109_, _25238_, _25236_);
  nand (_25239_, _25218_, _25200_);
  or (_25240_, _25239_, _25229_);
  nand (_25241_, _25240_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_25242_, _25188_, _18355_);
  nor (_25243_, _25242_, _25241_);
  and (_25244_, _25242_, ABINPUT[0]);
  or (_25245_, _25244_, _25209_);
  or (_25246_, _25245_, _25243_);
  not (_25247_, ABINPUT[10]);
  nand (_25248_, _25209_, _25247_);
  and (_25249_, _25248_, _27053_);
  and (_27111_, _25249_, _25246_);
  nand (_25250_, _25188_, _19646_);
  and (_25251_, _25250_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_25252_, _25188_, _19679_);
  or (_25253_, _25252_, _25209_);
  or (_25254_, _25253_, _25251_);
  not (_25255_, ABINPUT[9]);
  nand (_25256_, _25209_, _25255_);
  and (_25257_, _25256_, _27053_);
  and (_27113_, _25257_, _25254_);
  and (_25258_, _25208_, _24658_);
  and (_25259_, _25187_, _24658_);
  and (_25260_, _25259_, _18355_);
  nand (_25261_, _25260_, _18388_);
  or (_25262_, _25260_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_25263_, _25262_, _25261_);
  or (_25264_, _25263_, _25258_);
  nand (_25265_, _25258_, _25247_);
  and (_25266_, _25265_, _27053_);
  and (_27115_, _25266_, _25264_);
  and (_25267_, _25187_, _24483_);
  and (_25268_, _25267_, _24687_);
  and (_25269_, _25268_, _18355_);
  nand (_25270_, _25269_, _18388_);
  or (_25271_, _25269_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_25272_, _25271_, _25270_);
  and (_25273_, _25208_, _24680_);
  or (_25274_, _25273_, _25272_);
  nand (_25275_, _25273_, _25247_);
  and (_25276_, _25275_, _27053_);
  and (_27117_, _25276_, _25274_);
  nor (_25277_, _25114_, _25078_);
  and (_25278_, _25078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_25279_, _25278_, _25277_);
  and (_27993_, _25279_, _27053_);
  and (_25280_, _25078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_25281_, _25280_, _25277_);
  and (_27995_, _25281_, _27053_);
  and (_25282_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _27053_);
  and (_27997_, _25282_, _25078_);
  not (_25283_, _25104_);
  nor (_25284_, _25107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_25285_, _25284_, _25109_);
  or (_25286_, _25285_, _25102_);
  and (_25287_, _25286_, _25283_);
  and (_25288_, _25287_, _25141_);
  not (_25289_, _25083_);
  or (_25290_, _25087_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_25291_, _25290_, _25131_);
  or (_25292_, _25291_, _25081_);
  and (_25293_, _25292_, _25289_);
  and (_25294_, _25293_, _25100_);
  or (_25295_, _25294_, _25078_);
  or (_25296_, _25295_, _25288_);
  or (_25297_, _25123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_25298_, _25297_, _27053_);
  and (_27999_, _25298_, _25296_);
  not (_25299_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nand (_25300_, _25110_, _25299_);
  and (_25301_, _25300_, _25105_);
  and (_25302_, _25301_, _25141_);
  or (_25303_, _25090_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_25304_, _25303_, _25084_);
  and (_25305_, _25304_, _25100_);
  or (_25306_, _25305_, _25078_);
  or (_25307_, _25306_, _25302_);
  nand (_25308_, _25078_, _25299_);
  and (_25309_, _25308_, _27053_);
  and (_28001_, _25309_, _25307_);
  and (_25310_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _27053_);
  and (_28003_, _25310_, _25078_);
  and (_25311_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _27053_);
  and (_28005_, _25311_, _25078_);
  nand (_25312_, _25176_, _25114_);
  nor (_25313_, _25100_, _25078_);
  or (_25314_, _25313_, _25095_);
  and (_25315_, _25314_, _27053_);
  and (_28007_, _25315_, _25312_);
  not (_25316_, _25277_);
  and (_25317_, _25316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_25318_, _25135_);
  and (_25319_, _25318_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_25320_, _25089_, _25095_);
  or (_25321_, _25320_, _25081_);
  or (_25322_, _25321_, _25319_);
  not (_25323_, _25081_);
  or (_25324_, _25193_, _25323_);
  and (_25325_, _25324_, _25322_);
  or (_25326_, _25325_, _25083_);
  or (_25327_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _25095_);
  or (_25328_, _25327_, _25289_);
  and (_25329_, _25328_, _25100_);
  and (_25330_, _25329_, _25326_);
  not (_25331_, _25142_);
  and (_25332_, _25331_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_25333_, _25145_, _25102_);
  or (_25334_, _25333_, _25332_);
  not (_25335_, _25102_);
  or (_25336_, _25193_, _25335_);
  and (_25337_, _25336_, _25283_);
  and (_25338_, _25337_, _25334_);
  and (_25339_, _25327_, _25104_);
  or (_25340_, _25339_, _25338_);
  and (_25341_, _25340_, _25141_);
  or (_25342_, _25341_, _25330_);
  and (_25343_, _25342_, _25123_);
  or (_25344_, _25343_, _25317_);
  and (_28009_, _25344_, _27053_);
  and (_25345_, _25318_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_25346_, _25345_, _25321_);
  or (_25357_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _25095_);
  or (_25359_, _25357_, _25323_);
  and (_25360_, _25359_, _25346_);
  or (_25361_, _25360_, _25083_);
  or (_25362_, _25199_, _25289_);
  and (_25363_, _25362_, _25100_);
  and (_25364_, _25363_, _25361_);
  and (_25365_, _25114_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_25366_, _25365_, _25364_);
  and (_25367_, _25366_, _25123_);
  and (_25368_, _25078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_25369_, _25331_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_25370_, _25369_, _25333_);
  or (_25371_, _25357_, _25335_);
  and (_25372_, _25371_, _25283_);
  and (_25373_, _25372_, _25370_);
  and (_25374_, _25199_, _25104_);
  or (_25375_, _25374_, _25373_);
  and (_25376_, _25375_, _25141_);
  or (_25377_, _25376_, _25368_);
  or (_25378_, _25377_, _25367_);
  and (_28011_, _25378_, _27053_);
  and (_25379_, _25316_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  not (_25380_, _25158_);
  and (_25381_, _25380_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_25382_, _25089_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25383_, _25382_, _25081_);
  or (_25384_, _25383_, _25381_);
  or (_25385_, _25192_, _25323_);
  and (_25386_, _25385_, _25384_);
  or (_25387_, _25386_, _25083_);
  or (_25388_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25389_, _25388_, _25289_);
  and (_25390_, _25389_, _25100_);
  and (_25391_, _25390_, _25387_);
  not (_25392_, _25164_);
  and (_25393_, _25392_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_25394_, _25166_, _25102_);
  or (_25395_, _25394_, _25393_);
  or (_25396_, _25192_, _25335_);
  and (_25397_, _25396_, _25283_);
  and (_25398_, _25397_, _25395_);
  and (_25399_, _25388_, _25104_);
  or (_25400_, _25399_, _25398_);
  and (_25401_, _25400_, _25141_);
  or (_25402_, _25401_, _25391_);
  and (_25403_, _25402_, _25123_);
  or (_25404_, _25403_, _25379_);
  and (_28013_, _25404_, _27053_);
  and (_25405_, _25380_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_25406_, _25405_, _25383_);
  or (_25407_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_25408_, _25407_, _25323_);
  and (_25409_, _25408_, _25406_);
  or (_25410_, _25409_, _25083_);
  or (_25411_, _25198_, _25289_);
  and (_25412_, _25411_, _25100_);
  and (_25413_, _25412_, _25410_);
  and (_25414_, _25114_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_25415_, _25414_, _25413_);
  and (_25416_, _25415_, _25123_);
  and (_25417_, _25078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_25418_, _25392_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_25419_, _25418_, _25394_);
  or (_25420_, _25407_, _25335_);
  and (_25421_, _25420_, _25419_);
  or (_25422_, _25421_, _25104_);
  or (_25423_, _25198_, _25283_);
  and (_25424_, _25423_, _25422_);
  and (_25425_, _25424_, _25141_);
  or (_25426_, _25425_, _25417_);
  or (_25427_, _25426_, _25416_);
  and (_28015_, _25427_, _27053_);
  and (_25428_, _25179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or (_25429_, _25428_, _25178_);
  and (_28017_, _25429_, _27053_);
  and (_25430_, _25184_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or (_25431_, _25430_, _25183_);
  and (_28019_, _25431_, _27053_);
  nand (_25432_, _25188_, _18476_);
  and (_25433_, _25432_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_25434_, _25188_, _18617_);
  or (_25435_, _25434_, _25209_);
  or (_25436_, _25435_, _25433_);
  not (_25437_, ABINPUT[3]);
  nand (_25438_, _25209_, _25437_);
  and (_25439_, _25438_, _27053_);
  and (_28021_, _25439_, _25436_);
  nand (_25440_, _25188_, _18944_);
  nand (_25441_, _25440_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nor (_25442_, _25440_, _18388_);
  nor (_25443_, _25442_, _25209_);
  nand (_25444_, _25443_, _25441_);
  not (_25445_, ABINPUT[5]);
  nand (_25446_, _25209_, _25445_);
  and (_25447_, _25446_, _27053_);
  and (_28023_, _25447_, _25444_);
  nand (_25448_, _25188_, _19293_);
  and (_25449_, _25448_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_25450_, _25188_, _19337_);
  or (_25451_, _25450_, _25209_);
  or (_25452_, _25451_, _25449_);
  not (_25453_, ABINPUT[7]);
  nand (_25454_, _25209_, _25453_);
  and (_25455_, _25454_, _27053_);
  and (_28025_, _25455_, _25452_);
  nand (_25456_, _25259_, _18476_);
  and (_25457_, _25456_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_25458_, _25259_, _18617_);
  or (_25459_, _25458_, _25258_);
  or (_25460_, _25459_, _25457_);
  nand (_25461_, _25258_, _25437_);
  and (_25462_, _25461_, _27053_);
  and (_28027_, _25462_, _25460_);
  nand (_25463_, _25259_, _18759_);
  and (_25464_, _25463_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_25465_, _25259_, _18792_);
  or (_25466_, _25465_, _25258_);
  or (_25467_, _25466_, _25464_);
  nand (_25468_, _25258_, _24457_);
  and (_25469_, _25468_, _27053_);
  and (_28029_, _25469_, _25467_);
  nand (_25470_, _25259_, _18944_);
  and (_25471_, _25470_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_25472_, _25259_, _18977_);
  or (_25473_, _25472_, _25258_);
  or (_25474_, _25473_, _25471_);
  nand (_25475_, _25258_, _25445_);
  and (_25476_, _25475_, _27053_);
  and (_28031_, _25476_, _25474_);
  nand (_25477_, _25259_, _19119_);
  and (_25478_, _25477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_25479_, _25259_, _19152_);
  or (_25480_, _25479_, _25258_);
  or (_25481_, _25480_, _25478_);
  nand (_25482_, _25258_, _25211_);
  and (_25483_, _25482_, _27053_);
  and (_28033_, _25483_, _25481_);
  nand (_25484_, _25259_, _19293_);
  and (_25485_, _25484_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_25486_, _25259_, _19337_);
  or (_25487_, _25486_, _25258_);
  or (_25488_, _25487_, _25485_);
  nand (_25489_, _25258_, _25453_);
  and (_25490_, _25489_, _27053_);
  and (_28035_, _25490_, _25488_);
  nand (_25491_, _25259_, _19472_);
  and (_25492_, _25491_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_25493_, _25259_, _19505_);
  or (_25494_, _25493_, _25258_);
  or (_25495_, _25494_, _25492_);
  nand (_25496_, _25258_, _24502_);
  and (_25497_, _25496_, _27053_);
  and (_28037_, _25497_, _25495_);
  nand (_25498_, _25259_, _19646_);
  and (_25499_, _25498_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_25500_, _25259_, _19679_);
  or (_25501_, _25500_, _25258_);
  or (_25502_, _25501_, _25499_);
  nand (_25503_, _25258_, _25255_);
  and (_25504_, _25503_, _27053_);
  and (_28039_, _25504_, _25502_);
  and (_25505_, _25187_, _24679_);
  and (_25506_, _25505_, _24069_);
  nand (_25507_, _25506_, _18476_);
  and (_25508_, _25507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_25509_, _25268_, _18617_);
  or (_25510_, _25509_, _25273_);
  or (_25511_, _25510_, _25508_);
  nand (_25512_, _25273_, _25437_);
  and (_25513_, _25512_, _27053_);
  and (_28041_, _25513_, _25511_);
  nand (_25514_, _25506_, _18759_);
  and (_25515_, _25514_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_25516_, _25268_, _18792_);
  or (_25517_, _25516_, _25273_);
  or (_25518_, _25517_, _25515_);
  nand (_25519_, _25273_, _24457_);
  and (_25520_, _25519_, _27053_);
  and (_28043_, _25520_, _25518_);
  and (_25521_, _25268_, _18944_);
  or (_25522_, _25521_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nand (_25523_, _25521_, _18388_);
  and (_25524_, _25523_, _25522_);
  or (_25525_, _25524_, _25273_);
  nand (_25526_, _25273_, _25445_);
  and (_25527_, _25526_, _27053_);
  and (_28045_, _25527_, _25525_);
  nand (_25528_, _25506_, _19119_);
  and (_25529_, _25528_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_25530_, _25268_, _19152_);
  or (_25531_, _25530_, _25273_);
  or (_25532_, _25531_, _25529_);
  nand (_25533_, _25273_, _25211_);
  and (_25534_, _25533_, _27053_);
  and (_28047_, _25534_, _25532_);
  nand (_25535_, _25506_, _19293_);
  and (_25536_, _25535_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_25537_, _25268_, _19337_);
  or (_25538_, _25537_, _25273_);
  or (_25539_, _25538_, _25536_);
  nand (_25540_, _25273_, _25453_);
  and (_25541_, _25540_, _27053_);
  and (_28049_, _25541_, _25539_);
  nand (_25542_, _25506_, _19472_);
  and (_25543_, _25542_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_25544_, _25268_, _19505_);
  or (_25545_, _25544_, _25273_);
  or (_25546_, _25545_, _25543_);
  nand (_25547_, _25273_, _24502_);
  and (_25548_, _25547_, _27053_);
  and (_28051_, _25548_, _25546_);
  nand (_25549_, _25506_, _19646_);
  and (_25550_, _25549_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_25551_, _25268_, _19679_);
  or (_25552_, _25551_, _25273_);
  or (_25553_, _25552_, _25550_);
  nand (_25554_, _25273_, _25255_);
  and (_25555_, _25554_, _27053_);
  and (_28053_, _25555_, _25553_);
  and (_25556_, _16926_, _17285_);
  not (_25557_, _25556_);
  not (_25558_, _24005_);
  and (_25559_, _24005_, _23851_);
  and (_25560_, _25559_, _23378_);
  not (_25561_, _19887_);
  and (_25562_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_25563_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_25564_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_25565_, _25564_, _25563_);
  and (_25566_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_25567_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_25568_, _25567_, _25566_);
  and (_25569_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_25570_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_25571_, _25570_, _25569_);
  and (_25572_, _25571_, _25568_);
  and (_25573_, _25572_, _25565_);
  nor (_25574_, _19975_, _25561_);
  not (_25575_, _25574_);
  nor (_25576_, _25575_, _25573_);
  nor (_25577_, _25576_, _25562_);
  not (_25578_, _25577_);
  and (_25579_, _25578_, _25560_);
  nor (_25580_, _25579_, _25558_);
  nor (_25581_, _23851_, _23378_);
  and (_25582_, _25581_, _24005_);
  not (_25583_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_25584_, _24474_, _25583_);
  nor (_25585_, _25584_, _24488_);
  nor (_25586_, _25585_, _17753_);
  and (_25587_, _25585_, _17753_);
  nor (_25588_, _25587_, _25586_);
  nor (_25589_, _18092_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_25590_, _25589_, _18333_);
  and (_25591_, _25590_, _25556_);
  and (_25592_, _20315_, _18212_);
  nor (_25593_, _20315_, _18212_);
  nor (_25594_, _25593_, _25592_);
  and (_25595_, _25594_, _25591_);
  and (_25596_, _25595_, _25588_);
  nor (_25597_, _25585_, _20315_);
  and (_25598_, _25597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_25599_, _25585_, _20315_);
  and (_25600_, _25599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor (_25601_, _25600_, _25598_);
  nor (_25602_, _25585_, _20326_);
  and (_25603_, _25602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_25604_, _25585_, _20326_);
  and (_25605_, _25604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_25606_, _25605_, _25603_);
  and (_25607_, _25606_, _25601_);
  nor (_25608_, _25607_, _25596_);
  and (_25609_, _25596_, ABINPUT[10]);
  nor (_25610_, _25609_, _25608_);
  not (_25611_, _25610_);
  and (_25612_, _25611_, _25582_);
  nor (_25613_, _23851_, _23367_);
  and (_25614_, _25613_, _24005_);
  not (_25615_, _24288_);
  and (_25616_, _25615_, _25614_);
  nor (_25617_, _25616_, _25612_);
  and (_25618_, _25617_, _25580_);
  and (_25619_, _22892_, _22278_);
  and (_25620_, _25619_, _22409_);
  nor (_25621_, _25620_, _22727_);
  and (_25622_, _25621_, _22925_);
  and (_25623_, _22954_, _22409_);
  nor (_25624_, _23237_, _25623_);
  and (_25625_, _25624_, _22223_);
  and (_25626_, _22903_, _22409_);
  nor (_25627_, _25626_, _22497_);
  and (_25628_, _22409_, _22135_);
  nor (_25629_, _25628_, _22607_);
  and (_25630_, _25629_, _25627_);
  and (_25631_, _25630_, _25625_);
  and (_25632_, _25631_, _25622_);
  nor (_25633_, _25632_, _19843_);
  not (_25634_, _23227_);
  nor (_25635_, _25634_, _25624_);
  nor (_25636_, _25635_, _25633_);
  not (_25637_, _25636_);
  and (_25638_, _25637_, _25618_);
  and (_25639_, _25599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_25640_, _25597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_25641_, _25640_, _25639_);
  and (_25642_, _25602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_25643_, _25604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_25644_, _25643_, _25642_);
  and (_25645_, _25644_, _25641_);
  nor (_25646_, _25645_, _25596_);
  and (_25647_, _25596_, ABINPUT[6]);
  nor (_25648_, _25647_, _25646_);
  not (_25649_, _25648_);
  and (_25650_, _25649_, _25582_);
  not (_25651_, _25650_);
  not (_25652_, _24314_);
  and (_25653_, _25652_, _25614_);
  not (_25654_, _25653_);
  not (_25655_, _25585_);
  and (_25656_, _25559_, _23367_);
  and (_25657_, _25656_, _25655_);
  and (_25658_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_25659_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_25660_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_25661_, _25660_, _25659_);
  and (_25662_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_25663_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_25664_, _25663_, _25662_);
  and (_25665_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_25666_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_25667_, _25666_, _25665_);
  and (_25668_, _25667_, _25664_);
  and (_25669_, _25668_, _25661_);
  nor (_25670_, _25669_, _25575_);
  nor (_25671_, _25670_, _25658_);
  not (_25672_, _25671_);
  and (_25673_, _25672_, _25560_);
  nor (_25674_, _25673_, _25657_);
  and (_25675_, _25674_, _25654_);
  and (_25676_, _25675_, _25651_);
  not (_25677_, _25676_);
  and (_25678_, _25677_, _25638_);
  and (_25679_, _25597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_25680_, _25599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_25681_, _25680_, _25679_);
  and (_25682_, _25602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_25683_, _25604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_25684_, _25683_, _25682_);
  and (_25685_, _25684_, _25681_);
  nor (_25686_, _25685_, _25596_);
  and (_25687_, _25596_, ABINPUT[3]);
  nor (_25688_, _25687_, _25686_);
  not (_25689_, _25688_);
  and (_25690_, _25689_, _25582_);
  not (_25691_, _25690_);
  not (_25692_, _24296_);
  and (_25693_, _25692_, _25614_);
  not (_25694_, _25693_);
  and (_25695_, _25656_, _20315_);
  and (_25696_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_25697_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_25698_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_25699_, _25698_, _25697_);
  and (_25700_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_25701_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_25702_, _25701_, _25700_);
  and (_25703_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_25704_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_25705_, _25704_, _25703_);
  and (_25706_, _25705_, _25702_);
  and (_25707_, _25706_, _25699_);
  nor (_25708_, _25707_, _25575_);
  nor (_25709_, _25708_, _25696_);
  not (_25710_, _25709_);
  and (_25711_, _25710_, _25560_);
  nor (_25712_, _25711_, _25695_);
  and (_25713_, _25712_, _25694_);
  and (_25714_, _25713_, _25691_);
  nor (_25715_, _25714_, _25637_);
  nor (_25716_, _25715_, _25678_);
  and (_25717_, _17307_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_25718_, _25717_, _17753_);
  nor (_25719_, _18212_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_25720_, _25719_, _25718_);
  not (_25721_, _25720_);
  and (_25722_, _25721_, _25716_);
  nor (_25723_, _25722_, _25557_);
  and (_25724_, _25597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_25725_, _25599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_25726_, _25725_, _25724_);
  and (_25727_, _25602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_25728_, _25604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_25729_, _25728_, _25727_);
  and (_25730_, _25729_, _25726_);
  nor (_25731_, _25730_, _25596_);
  and (_25732_, _25596_, ABINPUT[8]);
  nor (_25733_, _25732_, _25731_);
  not (_25734_, _25733_);
  and (_25735_, _25734_, _25582_);
  not (_25736_, _25735_);
  and (_25737_, _24326_, _24005_);
  not (_25738_, _25737_);
  and (_25739_, _25738_, _25613_);
  not (_25740_, _25739_);
  and (_25741_, _25558_, _23851_);
  and (_25742_, _25741_, _23367_);
  and (_25743_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_25744_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_25745_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_25746_, _25745_, _25744_);
  and (_25747_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_25748_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_25749_, _25748_, _25747_);
  and (_25750_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_25751_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_25752_, _25751_, _25750_);
  and (_25753_, _25752_, _25749_);
  and (_25754_, _25753_, _25746_);
  nor (_25755_, _25754_, _25575_);
  nor (_25756_, _25755_, _25743_);
  not (_25757_, _25756_);
  and (_25758_, _25757_, _25560_);
  nor (_25759_, _25758_, _25742_);
  and (_25760_, _25759_, _25740_);
  and (_25761_, _25760_, _25736_);
  not (_25762_, _25761_);
  and (_25763_, _25762_, _25638_);
  not (_25764_, _24308_);
  and (_25765_, _25764_, _25614_);
  not (_25766_, _25765_);
  and (_25767_, _25656_, _20841_);
  and (_25768_, _25597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_25769_, _25599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_25770_, _25769_, _25768_);
  and (_25771_, _25602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_25772_, _25604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_25773_, _25772_, _25771_);
  and (_25774_, _25773_, _25770_);
  nor (_25775_, _25774_, _25596_);
  and (_25776_, _25596_, ABINPUT[5]);
  nor (_25777_, _25776_, _25775_);
  not (_25778_, _25777_);
  and (_25779_, _25778_, _25582_);
  and (_25780_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_25781_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_25782_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_25783_, _25782_, _25781_);
  and (_25784_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_25785_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_25786_, _25785_, _25784_);
  and (_25787_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_25788_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_25789_, _25788_, _25787_);
  and (_25790_, _25789_, _25786_);
  and (_25791_, _25790_, _25783_);
  nor (_25792_, _25791_, _25575_);
  nor (_25793_, _25792_, _25780_);
  not (_25794_, _25793_);
  and (_25795_, _25794_, _25560_);
  or (_25796_, _25795_, _25779_);
  nor (_25797_, _25796_, _25767_);
  and (_25798_, _25797_, _25766_);
  nor (_25799_, _25798_, _25637_);
  nor (_25800_, _25799_, _25763_);
  and (_25801_, _25717_, _24523_);
  nor (_25802_, _18081_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_25803_, _25802_, _25801_);
  not (_25804_, _25803_);
  and (_25805_, _25804_, _25800_);
  nor (_25806_, _25721_, _25716_);
  nor (_25807_, _25806_, _25805_);
  and (_25808_, _25807_, _25723_);
  not (_25809_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_25810_, _24474_, _25809_);
  nor (_25811_, _25810_, _24495_);
  not (_25812_, _25811_);
  and (_25813_, _25812_, _25656_);
  not (_25814_, _25813_);
  and (_25815_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_25816_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_25817_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_25818_, _25817_, _25816_);
  and (_25819_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_25820_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_25821_, _25820_, _25819_);
  and (_25822_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_25823_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_25824_, _25823_, _25822_);
  and (_25825_, _25824_, _25821_);
  and (_25826_, _25825_, _25818_);
  nor (_25827_, _25826_, _25575_);
  nor (_25828_, _25827_, _25815_);
  not (_25829_, _25828_);
  and (_25830_, _25829_, _25560_);
  nor (_25831_, _25830_, _25741_);
  and (_25832_, _25831_, _25814_);
  not (_25833_, _24320_);
  and (_25834_, _25833_, _25614_);
  and (_25835_, _25602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  not (_25836_, _25835_);
  and (_25837_, _25599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_25838_, _25597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_25839_, _25838_, _25837_);
  and (_25840_, _25839_, _25836_);
  and (_25841_, _25604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_25842_, _25841_, _25596_);
  and (_25843_, _25842_, _25840_);
  and (_25844_, _25596_, _25453_);
  or (_25845_, _25844_, _25843_);
  not (_25846_, _25845_);
  and (_25847_, _25846_, _25582_);
  nor (_25848_, _25847_, _25834_);
  and (_25849_, _25848_, _25832_);
  not (_25850_, _25849_);
  and (_25851_, _25850_, _25638_);
  and (_25852_, _25656_, _20589_);
  and (_25853_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_25854_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_25855_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_25856_, _25855_, _25854_);
  and (_25857_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_25858_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_25859_, _25858_, _25857_);
  and (_25860_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_25861_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_25862_, _25861_, _25860_);
  and (_25863_, _25862_, _25859_);
  and (_25864_, _25863_, _25856_);
  nor (_25865_, _25864_, _25575_);
  nor (_25866_, _25865_, _25853_);
  not (_25867_, _25866_);
  and (_25868_, _25867_, _25560_);
  nor (_25869_, _25868_, _25852_);
  and (_25870_, _25599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_25871_, _25597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_25872_, _25871_, _25870_);
  and (_25873_, _25602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_25874_, _25604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_25875_, _25874_, _25873_);
  and (_25876_, _25875_, _25872_);
  nor (_25877_, _25876_, _25596_);
  and (_25878_, _25596_, ABINPUT[4]);
  nor (_25879_, _25878_, _25877_);
  not (_25880_, _25879_);
  and (_25881_, _25880_, _25582_);
  not (_25882_, _25881_);
  and (_25883_, _25581_, _25558_);
  not (_25884_, _24302_);
  and (_25885_, _25884_, _25614_);
  nor (_25886_, _25885_, _25883_);
  and (_25887_, _25886_, _25882_);
  and (_25888_, _25887_, _25869_);
  nor (_25889_, _25888_, _25637_);
  nor (_25890_, _25889_, _25851_);
  and (_25891_, _25717_, _24483_);
  nor (_25892_, _18333_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_25893_, _25892_, _25891_);
  nand (_25894_, _25893_, _25890_);
  or (_25895_, _25893_, _25890_);
  and (_25896_, _25895_, _25894_);
  not (_25897_, _25896_);
  nor (_25898_, _25804_, _25800_);
  not (_25899_, _25898_);
  nor (_25900_, _25677_, _25638_);
  and (_25901_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_25902_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_25903_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_25904_, _25903_, _25902_);
  and (_25905_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_25906_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_25907_, _25906_, _25905_);
  and (_25908_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_25909_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_25910_, _25909_, _25908_);
  and (_25911_, _25910_, _25907_);
  and (_25912_, _25911_, _25904_);
  nor (_25913_, _25912_, _25575_);
  nor (_25914_, _25913_, _25901_);
  not (_25915_, _25914_);
  and (_25916_, _25915_, _25560_);
  nor (_25917_, _25581_, _24005_);
  nor (_25918_, _25917_, _25916_);
  and (_25919_, _25602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  not (_25920_, _25919_);
  and (_25921_, _25599_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_25922_, _25597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_25923_, _25922_, _25921_);
  and (_25924_, _25923_, _25920_);
  and (_25925_, _25604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_25926_, _25925_, _25596_);
  and (_25927_, _25926_, _25924_);
  and (_25928_, _25596_, _25255_);
  or (_25929_, _25928_, _25927_);
  not (_25930_, _25929_);
  and (_25931_, _25930_, _25582_);
  not (_25932_, _24332_);
  and (_25933_, _25932_, _25614_);
  nor (_25934_, _25933_, _25931_);
  and (_25935_, _25934_, _25918_);
  and (_25936_, _25935_, _25638_);
  nor (_25937_, _25936_, _25900_);
  nor (_25938_, _25717_, _17753_);
  and (_25939_, _25717_, _17579_);
  nor (_25940_, _25939_, _25938_);
  not (_25941_, _25940_);
  and (_25942_, _25941_, _25937_);
  nor (_25943_, _25941_, _25937_);
  nor (_25944_, _25943_, _25942_);
  and (_25945_, _25944_, _25899_);
  and (_25946_, _25945_, _25897_);
  and (_25947_, _25946_, _25808_);
  not (_25948_, _25800_);
  or (_25949_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  not (_25950_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nand (_25951_, _25716_, _25950_);
  and (_25952_, _25951_, _25890_);
  and (_25953_, _25952_, _25949_);
  not (_25954_, _25890_);
  not (_25955_, _25716_);
  and (_25956_, _25955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_25957_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_25958_, _25957_, _25956_);
  and (_25959_, _25958_, _25954_);
  or (_25960_, _25959_, _25953_);
  or (_25961_, _25960_, _25948_);
  not (_25962_, _25937_);
  and (_25963_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not (_25964_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor (_25965_, _25716_, _25964_);
  or (_25966_, _25965_, _25963_);
  and (_25967_, _25966_, _25890_);
  not (_25968_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_25969_, _25716_, _25968_);
  and (_25970_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_25971_, _25970_, _25969_);
  and (_25972_, _25971_, _25954_);
  or (_25973_, _25972_, _25967_);
  or (_25974_, _25973_, _25800_);
  and (_25975_, _25974_, _25962_);
  and (_25976_, _25975_, _25961_);
  not (_25977_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_25978_, _25716_, _25977_);
  or (_25979_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_25980_, _25979_, _25978_);
  and (_25981_, _25980_, _25890_);
  or (_25982_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_25983_, _25955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and (_25984_, _25983_, _25982_);
  and (_25985_, _25984_, _25954_);
  or (_25986_, _25985_, _25981_);
  or (_25987_, _25986_, _25948_);
  not (_25988_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_25989_, _25716_, _25988_);
  or (_25990_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_25991_, _25990_, _25989_);
  and (_25992_, _25991_, _25890_);
  or (_25993_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_25994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_25995_, _25716_, _25994_);
  and (_25996_, _25995_, _25993_);
  and (_25997_, _25996_, _25954_);
  or (_25998_, _25997_, _25992_);
  or (_25999_, _25998_, _25800_);
  and (_26000_, _25999_, _25937_);
  and (_26001_, _26000_, _25987_);
  or (_26002_, _26001_, _25976_);
  or (_26003_, _26002_, _25947_);
  not (_26004_, _25947_);
  or (_26005_, _26004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_26006_, _26005_, _27053_);
  and (_28138_, _26006_, _26003_);
  nor (_26007_, _25720_, _25557_);
  nor (_26008_, _25893_, _25557_);
  and (_26009_, _26008_, _26007_);
  and (_26010_, _25940_, _25556_);
  nor (_26011_, _25803_, _25557_);
  and (_26012_, _26011_, _26010_);
  and (_26013_, _26012_, _26009_);
  or (_26014_, _26013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_26015_, _26013_);
  and (_26016_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26017_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26018_, _26017_, _26016_);
  and (_26019_, _26018_, ABINPUT[0]);
  not (_26020_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_26021_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_26022_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_26023_, _26022_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_26024_, _26023_, _26021_);
  and (_26025_, _26016_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_26026_, _26025_);
  and (_26027_, _26026_, _26024_);
  or (_26028_, _26027_, _26020_);
  or (_26029_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , ABINPUT[10]);
  and (_26030_, _26029_, _26028_);
  or (_26031_, _26030_, _26019_);
  and (_26032_, _26031_, _25556_);
  or (_26033_, _26032_, _26015_);
  and (_28150_, _26033_, _26014_);
  not (_26034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_26035_, _26011_, _26010_);
  nor (_26036_, _26008_, _26007_);
  and (_26037_, _26036_, _25556_);
  and (_26038_, _26037_, _26035_);
  nor (_26039_, _26038_, _26034_);
  not (_26040_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_26041_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _26040_);
  nor (_26042_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26043_, _26042_, _26041_);
  and (_26044_, _26043_, ABINPUT[0]);
  and (_26045_, _26020_, ABINPUT[3]);
  or (_26046_, _26045_, _26044_);
  and (_26047_, _26042_, _26040_);
  nor (_26048_, _26047_, _26020_);
  nor (_26049_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_26050_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _26022_);
  nor (_26051_, _26050_, _26049_);
  and (_26052_, _26051_, _26048_);
  or (_26053_, _26052_, _26046_);
  and (_26054_, _26053_, _25556_);
  and (_26055_, _26054_, _26038_);
  or (_28438_, _26055_, _26039_);
  not (_26056_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_26057_, _26038_, _26056_);
  nor (_26058_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_26059_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _26022_);
  nor (_26060_, _26059_, _26058_);
  not (_26061_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  nor (_26062_, _26061_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26063_, _26062_, _26040_);
  nor (_26064_, _26063_, _26020_);
  and (_26065_, _26064_, _26060_);
  and (_26066_, _26062_, _26041_);
  and (_26067_, _26066_, ABINPUT[0]);
  and (_26068_, _26020_, ABINPUT[4]);
  or (_26069_, _26068_, _26067_);
  or (_26070_, _26069_, _26065_);
  and (_26071_, _26070_, _25556_);
  and (_26072_, _26071_, _26038_);
  or (_28444_, _26072_, _26057_);
  not (_26073_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_26074_, _26038_, _26073_);
  nor (_26075_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  nor (_26076_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _26022_);
  nor (_26077_, _26076_, _26075_);
  and (_26078_, _26061_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_26079_, _26078_, _26040_);
  nor (_26080_, _26079_, _26020_);
  and (_26081_, _26080_, _26077_);
  and (_26082_, _26041_, _26078_);
  and (_26083_, _26082_, ABINPUT[0]);
  and (_26084_, _26020_, ABINPUT[5]);
  or (_26085_, _26084_, _26083_);
  or (_26086_, _26085_, _26081_);
  and (_26087_, _26086_, _25556_);
  and (_26088_, _26087_, _26038_);
  or (_28450_, _26088_, _26074_);
  not (_26089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_26090_, _26038_, _26089_);
  and (_26091_, _26041_, _26016_);
  and (_26092_, _26091_, ABINPUT[0]);
  nor (_26093_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_26094_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _26022_);
  nor (_26095_, _26094_, _26093_);
  and (_26096_, _26016_, _26040_);
  not (_26097_, _26096_);
  and (_26098_, _26097_, _26095_);
  or (_26099_, _26098_, _26020_);
  or (_26100_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , ABINPUT[6]);
  and (_26101_, _26100_, _26099_);
  or (_26102_, _26101_, _26092_);
  and (_26103_, _26102_, _25556_);
  and (_26104_, _26103_, _26038_);
  or (_28456_, _26104_, _26090_);
  not (_26105_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_26106_, _26038_, _26105_);
  nor (_26107_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_26108_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _26022_);
  nor (_26109_, _26108_, _26107_);
  and (_26110_, _26042_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_26111_, _26110_, _26020_);
  and (_26112_, _26111_, _26109_);
  and (_26113_, _26042_, _26017_);
  and (_26114_, _26113_, ABINPUT[0]);
  and (_26115_, _26020_, ABINPUT[7]);
  or (_26116_, _26115_, _26114_);
  or (_26117_, _26116_, _26112_);
  and (_26118_, _26117_, _25556_);
  and (_26119_, _26118_, _26038_);
  or (_28462_, _26119_, _26106_);
  not (_26120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_26121_, _26038_, _26120_);
  nor (_26122_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_26123_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _26022_);
  nor (_26124_, _26123_, _26122_);
  and (_26125_, _26062_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_26126_, _26125_, _26020_);
  and (_26127_, _26126_, _26124_);
  and (_26128_, _26062_, _26017_);
  and (_26129_, _26128_, ABINPUT[0]);
  and (_26130_, _26020_, ABINPUT[8]);
  or (_26131_, _26130_, _26129_);
  or (_26132_, _26131_, _26127_);
  and (_26133_, _26132_, _25556_);
  and (_26134_, _26133_, _26038_);
  or (_28467_, _26134_, _26121_);
  not (_26135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_26136_, _26038_, _26135_);
  nor (_26137_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_26138_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _26022_);
  nor (_26139_, _26138_, _26137_);
  and (_26140_, _26078_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_26141_, _26140_, _26020_);
  and (_26142_, _26141_, _26139_);
  and (_26143_, _26078_, _26017_);
  and (_26144_, _26143_, ABINPUT[0]);
  and (_26145_, _26020_, ABINPUT[9]);
  or (_26146_, _26145_, _26144_);
  or (_26147_, _26146_, _26142_);
  and (_26148_, _26147_, _25556_);
  and (_26149_, _26148_, _26038_);
  or (_28473_, _26149_, _26136_);
  nor (_26150_, _26038_, _25950_);
  and (_26151_, _26038_, _26032_);
  or (_28476_, _26151_, _26150_);
  not (_26152_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_26153_, _26007_, _25893_);
  and (_26154_, _26153_, _26035_);
  nor (_26155_, _26154_, _26152_);
  and (_26156_, _26154_, _26054_);
  or (_28484_, _26156_, _26155_);
  or (_26157_, _26154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  not (_26158_, _26154_);
  or (_26159_, _26158_, _26071_);
  and (_28488_, _26159_, _26157_);
  not (_26160_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_26161_, _26154_, _26160_);
  and (_26162_, _26154_, _26087_);
  or (_28492_, _26162_, _26161_);
  not (_26163_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_26164_, _26154_, _26163_);
  and (_26165_, _26154_, _26103_);
  or (_28496_, _26165_, _26164_);
  not (_26166_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_26167_, _26154_, _26166_);
  and (_26168_, _26154_, _26118_);
  or (_28500_, _26168_, _26167_);
  not (_26169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_26170_, _26154_, _26169_);
  and (_26171_, _26154_, _26133_);
  or (_28504_, _26171_, _26170_);
  not (_26172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_26173_, _26154_, _26172_);
  and (_26174_, _26154_, _26148_);
  or (_28507_, _26174_, _26173_);
  or (_26175_, _26154_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_26176_, _26158_, _26032_);
  and (_28510_, _26176_, _26175_);
  not (_26177_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_26178_, _26008_, _25720_);
  and (_26179_, _26178_, _26035_);
  nor (_26180_, _26179_, _26177_);
  and (_26181_, _26179_, _26054_);
  or (_28518_, _26181_, _26180_);
  or (_26182_, _26179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  not (_26183_, _26179_);
  or (_26184_, _26183_, _26071_);
  and (_28522_, _26184_, _26182_);
  not (_26185_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_26186_, _26179_, _26185_);
  and (_26187_, _26179_, _26087_);
  or (_28526_, _26187_, _26186_);
  or (_26188_, _26179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_26189_, _26183_, _26103_);
  and (_28530_, _26189_, _26188_);
  not (_26190_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_26191_, _26179_, _26190_);
  and (_26192_, _26179_, _26118_);
  or (_28534_, _26192_, _26191_);
  and (_26193_, _26183_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_26194_, _26179_, _26133_);
  or (_28538_, _26194_, _26193_);
  not (_26195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_26196_, _26179_, _26195_);
  and (_26197_, _26179_, _26148_);
  or (_28542_, _26197_, _26196_);
  or (_26198_, _26179_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_26199_, _26183_, _26032_);
  and (_28545_, _26199_, _26198_);
  not (_26200_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_26201_, _26035_, _26009_);
  nor (_26202_, _26201_, _26200_);
  and (_26203_, _26201_, _26054_);
  or (_28551_, _26203_, _26202_);
  or (_26204_, _26201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  not (_26205_, _26201_);
  or (_26206_, _26205_, _26071_);
  and (_28554_, _26206_, _26204_);
  not (_26207_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_26208_, _26201_, _26207_);
  and (_26209_, _26201_, _26087_);
  or (_28558_, _26209_, _26208_);
  or (_26210_, _26201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_26211_, _26205_, _26103_);
  and (_28562_, _26211_, _26210_);
  not (_26212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_26213_, _26201_, _26212_);
  and (_26214_, _26201_, _26118_);
  or (_28566_, _26214_, _26213_);
  or (_26215_, _26201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_26216_, _26205_, _26133_);
  and (_28570_, _26216_, _26215_);
  not (_26217_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_26218_, _26201_, _26217_);
  and (_26219_, _26201_, _26148_);
  or (_28574_, _26219_, _26218_);
  or (_26220_, _26201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_26221_, _26205_, _26032_);
  and (_28577_, _26221_, _26220_);
  not (_26222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_26223_, _26011_, _25941_);
  and (_26224_, _26223_, _26036_);
  nor (_26225_, _26224_, _26222_);
  and (_26226_, _26224_, _26054_);
  or (_28585_, _26226_, _26225_);
  not (_26227_, _26224_);
  and (_26228_, _26227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  and (_26229_, _26224_, _26071_);
  or (_28589_, _26229_, _26228_);
  not (_26230_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_26231_, _26224_, _26230_);
  and (_26232_, _26224_, _26087_);
  or (_28593_, _26232_, _26231_);
  or (_26233_, _26224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_26234_, _26227_, _26103_);
  and (_28597_, _26234_, _26233_);
  not (_26235_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_26236_, _26224_, _26235_);
  and (_26237_, _26224_, _26118_);
  or (_28600_, _26237_, _26236_);
  or (_26238_, _26224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_26239_, _26227_, _26133_);
  and (_28604_, _26239_, _26238_);
  not (_26241_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_26242_, _26224_, _26241_);
  and (_26243_, _26224_, _26148_);
  or (_28608_, _26243_, _26242_);
  or (_26244_, _26224_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_26245_, _26227_, _26032_);
  and (_28611_, _26245_, _26244_);
  not (_26246_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_26247_, _26223_, _26153_);
  nor (_26248_, _26247_, _26246_);
  and (_26250_, _26247_, _26054_);
  or (_28616_, _26250_, _26248_);
  not (_26251_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_26252_, _26247_, _26251_);
  and (_26253_, _26247_, _26071_);
  or (_28620_, _26253_, _26252_);
  not (_26254_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_26255_, _26247_, _26254_);
  and (_26256_, _26247_, _26087_);
  or (_28624_, _26256_, _26255_);
  not (_26258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_26259_, _26247_, _26258_);
  and (_26260_, _26247_, _26103_);
  or (_28628_, _26260_, _26259_);
  not (_26261_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_26262_, _26247_, _26261_);
  and (_26263_, _26247_, _26118_);
  or (_28632_, _26263_, _26262_);
  or (_26264_, _26247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  not (_26265_, _26247_);
  or (_26267_, _26265_, _26133_);
  and (_28636_, _26267_, _26264_);
  not (_26268_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_26269_, _26247_, _26268_);
  and (_26270_, _26247_, _26148_);
  or (_28640_, _26270_, _26269_);
  nor (_26271_, _26247_, _25964_);
  and (_26272_, _26247_, _26032_);
  or (_28643_, _26272_, _26271_);
  not (_26273_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_26275_, _26223_, _26178_);
  nor (_26276_, _26275_, _26273_);
  and (_26277_, _26275_, _26054_);
  or (_28647_, _26277_, _26276_);
  not (_26278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_26279_, _26275_, _26278_);
  and (_26280_, _26275_, _26071_);
  or (_28651_, _26280_, _26279_);
  not (_26281_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_26282_, _26275_, _26281_);
  and (_26284_, _26275_, _26087_);
  or (_28655_, _26284_, _26282_);
  or (_26285_, _26275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  not (_26286_, _26275_);
  or (_26287_, _26286_, _26103_);
  and (_28659_, _26287_, _26285_);
  not (_26288_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_26289_, _26275_, _26288_);
  and (_26290_, _26275_, _26118_);
  or (_28663_, _26290_, _26289_);
  or (_26292_, _26275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_26293_, _26286_, _26133_);
  and (_28667_, _26293_, _26292_);
  not (_26294_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_26295_, _26275_, _26294_);
  and (_26296_, _26275_, _26148_);
  or (_28671_, _26296_, _26295_);
  or (_26297_, _26275_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_26298_, _26286_, _26032_);
  and (_28674_, _26298_, _26297_);
  not (_26299_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_26300_, _26223_, _26009_);
  nor (_26301_, _26300_, _26299_);
  and (_26302_, _26300_, _26054_);
  or (_28679_, _26302_, _26301_);
  or (_26303_, _26300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  not (_26304_, _26300_);
  or (_26305_, _26304_, _26071_);
  and (_28683_, _26305_, _26303_);
  not (_26306_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_26307_, _26300_, _26306_);
  and (_26308_, _26300_, _26087_);
  or (_28687_, _26308_, _26307_);
  not (_26309_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_26310_, _26300_, _26309_);
  and (_26311_, _26300_, _26103_);
  or (_28690_, _26311_, _26310_);
  not (_26312_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_26313_, _26300_, _26312_);
  and (_26314_, _26300_, _26118_);
  or (_28694_, _26314_, _26313_);
  not (_26315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_26316_, _26300_, _26315_);
  and (_26317_, _26300_, _26133_);
  or (_28698_, _26317_, _26316_);
  not (_26318_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_26319_, _26300_, _26318_);
  and (_26320_, _26300_, _26148_);
  or (_28702_, _26320_, _26319_);
  nor (_26321_, _26300_, _25968_);
  and (_26322_, _26300_, _26032_);
  or (_28705_, _26322_, _26321_);
  not (_26323_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_26324_, _26010_, _25803_);
  and (_26325_, _26324_, _26036_);
  nor (_26326_, _26325_, _26323_);
  and (_26327_, _26325_, _26054_);
  or (_28713_, _26327_, _26326_);
  not (_26328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_26329_, _26325_, _26328_);
  and (_26330_, _26325_, _26071_);
  or (_28717_, _26330_, _26329_);
  not (_26331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_26332_, _26325_, _26331_);
  and (_26333_, _26325_, _26087_);
  or (_28721_, _26333_, _26332_);
  or (_26334_, _26325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  not (_26335_, _26325_);
  or (_26336_, _26335_, _26103_);
  and (_28725_, _26336_, _26334_);
  not (_26337_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_26338_, _26325_, _26337_);
  and (_26339_, _26325_, _26118_);
  or (_28729_, _26339_, _26338_);
  not (_26340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_26341_, _26325_, _26340_);
  and (_26342_, _26325_, _26133_);
  or (_28733_, _26342_, _26341_);
  not (_26343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_26344_, _26325_, _26343_);
  and (_26345_, _26325_, _26148_);
  or (_28736_, _26345_, _26344_);
  nor (_26346_, _26325_, _25977_);
  and (_26347_, _26325_, _26032_);
  or (_28739_, _26347_, _26346_);
  not (_26348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_26349_, _26324_, _26153_);
  nor (_26350_, _26349_, _26348_);
  and (_26351_, _26349_, _26054_);
  or (_28743_, _26351_, _26350_);
  or (_26352_, _26349_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  not (_26353_, _26349_);
  or (_26354_, _26353_, _26071_);
  and (_28744_, _26354_, _26352_);
  not (_26355_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_26356_, _26349_, _26355_);
  and (_26357_, _26349_, _26087_);
  or (_28746_, _26357_, _26356_);
  not (_26358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_26359_, _26349_, _26358_);
  and (_26360_, _26349_, _26103_);
  or (_28750_, _26360_, _26359_);
  not (_26361_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_26362_, _26349_, _26361_);
  and (_26363_, _26349_, _26118_);
  or (_28754_, _26363_, _26362_);
  and (_26364_, _26353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_26365_, _26349_, _26133_);
  or (_28758_, _26365_, _26364_);
  not (_26366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_26367_, _26349_, _26366_);
  and (_26368_, _26349_, _26148_);
  or (_28762_, _26368_, _26367_);
  and (_26369_, _26353_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_26370_, _26349_, _26032_);
  or (_28772_, _26370_, _26369_);
  not (_26371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_26372_, _26324_, _26178_);
  nor (_26373_, _26372_, _26371_);
  and (_26374_, _26372_, _26054_);
  or (_28791_, _26374_, _26373_);
  or (_26375_, _26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  not (_26376_, _26372_);
  or (_26377_, _26376_, _26071_);
  and (_28807_, _26377_, _26375_);
  not (_26378_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_26379_, _26372_, _26378_);
  and (_26380_, _26372_, _26087_);
  or (_28820_, _26380_, _26379_);
  or (_26381_, _26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_26382_, _26376_, _26103_);
  and (_28838_, _26382_, _26381_);
  not (_26383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_26384_, _26372_, _26383_);
  and (_26385_, _26372_, _26118_);
  or (_28849_, _26385_, _26384_);
  not (_26386_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_26387_, _26372_, _26386_);
  and (_26388_, _26372_, _26133_);
  or (_28866_, _26388_, _26387_);
  not (_26393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_26396_, _26372_, _26393_);
  and (_26401_, _26372_, _26148_);
  or (_28885_, _26401_, _26396_);
  or (_26405_, _26372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_26408_, _26376_, _26032_);
  and (_28895_, _26408_, _26405_);
  not (_26413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_26416_, _26324_, _26009_);
  nor (_26421_, _26416_, _26413_);
  and (_26423_, _26416_, _26054_);
  or (_28921_, _26423_, _26421_);
  or (_26424_, _26416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  not (_26425_, _26416_);
  or (_26426_, _26425_, _26071_);
  and (_28939_, _26426_, _26424_);
  not (_26427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_26428_, _26416_, _26427_);
  and (_26429_, _26416_, _26087_);
  or (_28957_, _26429_, _26428_);
  not (_26430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_26431_, _26416_, _26430_);
  and (_26432_, _26416_, _26103_);
  or (_28978_, _26432_, _26431_);
  not (_26433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_26434_, _26416_, _26433_);
  and (_26435_, _26416_, _26118_);
  or (_28998_, _26435_, _26434_);
  and (_26436_, _26425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_26437_, _26416_, _26133_);
  or (_29012_, _26437_, _26436_);
  not (_26438_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_26439_, _26416_, _26438_);
  and (_26440_, _26416_, _26148_);
  or (_29016_, _26440_, _26439_);
  or (_26441_, _26416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_26442_, _26425_, _26032_);
  and (_29019_, _26442_, _26441_);
  not (_26443_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_26444_, _26036_, _26012_);
  nor (_26445_, _26444_, _26443_);
  and (_26446_, _26444_, _26054_);
  or (_29025_, _26446_, _26445_);
  or (_26447_, _26444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  not (_26448_, _26444_);
  or (_26449_, _26448_, _26071_);
  and (_29029_, _26449_, _26447_);
  not (_26450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor (_26451_, _26444_, _26450_);
  and (_26452_, _26444_, _26087_);
  or (_29033_, _26452_, _26451_);
  not (_26453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_26454_, _26444_, _26453_);
  and (_26455_, _26444_, _26103_);
  or (_29037_, _26455_, _26454_);
  not (_26456_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_26457_, _26444_, _26456_);
  and (_26458_, _26444_, _26118_);
  or (_29041_, _26458_, _26457_);
  not (_26459_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_26460_, _26444_, _26459_);
  and (_26461_, _26444_, _26133_);
  or (_29045_, _26461_, _26460_);
  not (_26463_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_26465_, _26444_, _26463_);
  and (_26467_, _26444_, _26148_);
  or (_29049_, _26467_, _26465_);
  nor (_26470_, _26444_, _25988_);
  and (_26472_, _26444_, _26032_);
  or (_29052_, _26472_, _26470_);
  not (_26475_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_26477_, _26153_, _26012_);
  nor (_26479_, _26477_, _26475_);
  and (_26481_, _26477_, _26054_);
  or (_29057_, _26481_, _26479_);
  not (_26484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_26486_, _26477_, _26484_);
  and (_26488_, _26477_, _26071_);
  or (_29061_, _26488_, _26486_);
  not (_26491_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_26493_, _26477_, _26491_);
  and (_26495_, _26477_, _26087_);
  or (_29065_, _26495_, _26493_);
  not (_26498_, _26477_);
  and (_26500_, _26498_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_26502_, _26477_, _26103_);
  or (_29069_, _26502_, _26500_);
  not (_26505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_26507_, _26477_, _26505_);
  and (_26509_, _26477_, _26118_);
  or (_29072_, _26509_, _26507_);
  or (_26511_, _26477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_26512_, _26498_, _26133_);
  and (_29074_, _26512_, _26511_);
  not (_26513_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_26514_, _26477_, _26513_);
  and (_26515_, _26477_, _26148_);
  or (_29078_, _26515_, _26514_);
  or (_26516_, _26477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_26517_, _26498_, _26032_);
  and (_29081_, _26517_, _26516_);
  not (_26518_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_26519_, _26178_, _26012_);
  nor (_26520_, _26519_, _26518_);
  and (_26521_, _26519_, _26054_);
  or (_29086_, _26521_, _26520_);
  or (_26522_, _26519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  not (_26523_, _26519_);
  or (_26524_, _26523_, _26071_);
  and (_29090_, _26524_, _26522_);
  not (_26525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_26526_, _26519_, _26525_);
  and (_26527_, _26519_, _26087_);
  or (_29094_, _26527_, _26526_);
  not (_26528_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_26529_, _26519_, _26528_);
  and (_26530_, _26519_, _26103_);
  or (_29098_, _26530_, _26529_);
  not (_26531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_26532_, _26519_, _26531_);
  and (_26533_, _26519_, _26118_);
  or (_29102_, _26533_, _26532_);
  or (_26534_, _26519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_26535_, _26523_, _26133_);
  and (_29106_, _26535_, _26534_);
  not (_26536_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_26537_, _26519_, _26536_);
  and (_26538_, _26519_, _26148_);
  or (_29110_, _26538_, _26537_);
  nor (_26539_, _26519_, _25994_);
  and (_26540_, _26519_, _26032_);
  or (_29113_, _26540_, _26539_);
  not (_26541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_26542_, _26013_, _26541_);
  and (_26543_, _26054_, _26013_);
  or (_29118_, _26543_, _26542_);
  not (_26544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_26545_, _26013_, _26544_);
  and (_26546_, _26071_, _26013_);
  or (_29122_, _26546_, _26545_);
  not (_26547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_26548_, _26013_, _26547_);
  and (_26549_, _26087_, _26013_);
  or (_29126_, _26549_, _26548_);
  and (_26550_, _26015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_26551_, _26103_, _26013_);
  or (_29130_, _26551_, _26550_);
  not (_26552_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_26553_, _26013_, _26552_);
  and (_26554_, _26118_, _26013_);
  or (_29134_, _26554_, _26553_);
  not (_26555_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_26556_, _26013_, _26555_);
  and (_26557_, _26133_, _26013_);
  or (_29138_, _26557_, _26556_);
  not (_26558_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_26559_, _26013_, _26558_);
  and (_26560_, _26148_, _26013_);
  or (_29142_, _26560_, _26559_);
  and (_26561_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_26562_, _25716_, _26152_);
  or (_26563_, _26562_, _26561_);
  and (_26564_, _26563_, _25890_);
  nor (_26565_, _25716_, _26200_);
  and (_26566_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_26567_, _26566_, _26565_);
  and (_26568_, _26567_, _25954_);
  or (_26569_, _26568_, _26564_);
  or (_26570_, _26569_, _25948_);
  and (_26571_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_26572_, _25716_, _26246_);
  or (_26573_, _26572_, _26571_);
  and (_26574_, _26573_, _25890_);
  nor (_26575_, _25716_, _26299_);
  and (_26576_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_26577_, _26576_, _26575_);
  and (_26578_, _26577_, _25954_);
  or (_26579_, _26578_, _26574_);
  or (_26580_, _26579_, _25800_);
  and (_26581_, _26580_, _25962_);
  and (_26582_, _26581_, _26570_);
  nand (_26583_, _25716_, _26323_);
  or (_26584_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_26585_, _26584_, _26583_);
  and (_26586_, _26585_, _25890_);
  or (_26587_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand (_26588_, _25716_, _26371_);
  and (_26589_, _26588_, _26587_);
  and (_26590_, _26589_, _25954_);
  or (_26591_, _26590_, _26586_);
  or (_26592_, _26591_, _25948_);
  nand (_26593_, _25716_, _26443_);
  or (_26594_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_26595_, _26594_, _26593_);
  and (_26596_, _26595_, _25890_);
  or (_26597_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand (_26598_, _25716_, _26518_);
  and (_26599_, _26598_, _26597_);
  and (_26600_, _26599_, _25954_);
  or (_26601_, _26600_, _26596_);
  or (_26602_, _26601_, _25800_);
  and (_26603_, _26602_, _25937_);
  and (_26604_, _26603_, _26592_);
  or (_26605_, _26604_, _26582_);
  or (_26606_, _26605_, _25947_);
  or (_26607_, _26004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_26608_, _26607_, _27053_);
  and (_00044_, _26608_, _26606_);
  or (_26609_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_26610_, _25716_, _26056_);
  and (_26611_, _26610_, _25890_);
  and (_26612_, _26611_, _26609_);
  and (_26613_, _25955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_26614_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_26615_, _26614_, _26613_);
  and (_26616_, _26615_, _25954_);
  or (_26617_, _26616_, _26612_);
  or (_26618_, _26617_, _25948_);
  and (_26619_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_26620_, _25716_, _26251_);
  or (_26621_, _26620_, _26619_);
  and (_26622_, _26621_, _25890_);
  or (_26623_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nand (_26624_, _25716_, _26278_);
  and (_26625_, _26624_, _26623_);
  and (_26626_, _26625_, _25954_);
  or (_26627_, _26626_, _26622_);
  or (_26628_, _26627_, _25800_);
  and (_26629_, _26628_, _25962_);
  and (_26630_, _26629_, _26618_);
  nand (_26631_, _25716_, _26328_);
  or (_26632_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_26633_, _26632_, _26631_);
  and (_26634_, _26633_, _25890_);
  or (_26635_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_26636_, _25955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_26637_, _26636_, _26635_);
  and (_26638_, _26637_, _25954_);
  or (_26639_, _26638_, _26634_);
  or (_26640_, _26639_, _25948_);
  and (_26641_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_26642_, _25716_, _26484_);
  or (_26643_, _26642_, _26641_);
  and (_26644_, _26643_, _25890_);
  and (_26645_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_26646_, _25716_, _26544_);
  or (_26647_, _26646_, _26645_);
  and (_26648_, _26647_, _25954_);
  or (_26649_, _26648_, _26644_);
  or (_26650_, _26649_, _25800_);
  and (_26651_, _26650_, _25937_);
  and (_26652_, _26651_, _26640_);
  or (_26653_, _26652_, _26630_);
  or (_26654_, _26653_, _25947_);
  or (_26655_, _26004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_26656_, _26655_, _27053_);
  and (_00046_, _26656_, _26654_);
  and (_26657_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_26658_, _25716_, _26160_);
  or (_26659_, _26658_, _26657_);
  and (_26660_, _26659_, _25890_);
  nor (_26661_, _25716_, _26207_);
  and (_26662_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_26663_, _26662_, _26661_);
  and (_26664_, _26663_, _25954_);
  or (_26665_, _26664_, _26660_);
  or (_26666_, _26665_, _25948_);
  and (_26667_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_26668_, _25716_, _26254_);
  or (_26669_, _26668_, _26667_);
  and (_26670_, _26669_, _25890_);
  nor (_26671_, _25716_, _26306_);
  and (_26672_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_26673_, _26672_, _26671_);
  and (_26674_, _26673_, _25954_);
  or (_26675_, _26674_, _26670_);
  or (_26676_, _26675_, _25800_);
  and (_26677_, _26676_, _25962_);
  and (_26678_, _26677_, _26666_);
  nand (_26679_, _25716_, _26331_);
  or (_26680_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_26681_, _26680_, _26679_);
  and (_26682_, _26681_, _25890_);
  or (_26683_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_26684_, _25716_, _26378_);
  and (_26685_, _26684_, _26683_);
  and (_26686_, _26685_, _25954_);
  or (_26687_, _26686_, _26682_);
  or (_26688_, _26687_, _25948_);
  nand (_26689_, _25716_, _26450_);
  or (_26690_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_26691_, _26690_, _26689_);
  and (_26692_, _26691_, _25890_);
  or (_26693_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_26694_, _25716_, _26525_);
  and (_26695_, _26694_, _26693_);
  and (_26696_, _26695_, _25954_);
  or (_26697_, _26696_, _26692_);
  or (_26698_, _26697_, _25800_);
  and (_26699_, _26698_, _25937_);
  and (_26700_, _26699_, _26688_);
  or (_26701_, _26700_, _26678_);
  or (_26702_, _26701_, _25947_);
  or (_26703_, _26004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_26704_, _26703_, _27053_);
  and (_00048_, _26704_, _26702_);
  and (_26705_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_26706_, _25716_, _26163_);
  or (_26707_, _26706_, _26705_);
  and (_26708_, _26707_, _25890_);
  and (_26709_, _25955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_26710_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_26711_, _26710_, _26709_);
  and (_26712_, _26711_, _25954_);
  or (_26713_, _26712_, _26708_);
  or (_26714_, _26713_, _25948_);
  and (_26715_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_26716_, _25716_, _26258_);
  or (_26717_, _26716_, _26715_);
  and (_26718_, _26717_, _25890_);
  nor (_26719_, _25716_, _26309_);
  and (_26720_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_26721_, _26720_, _26719_);
  and (_26722_, _26721_, _25954_);
  or (_26723_, _26722_, _26718_);
  or (_26724_, _26723_, _25800_);
  and (_26725_, _26724_, _25962_);
  and (_26726_, _26725_, _26714_);
  and (_26727_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_26728_, _25716_, _26358_);
  or (_26729_, _26728_, _26727_);
  and (_26730_, _26729_, _25890_);
  and (_26731_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_26732_, _25716_, _26430_);
  or (_26733_, _26732_, _26731_);
  and (_26734_, _26733_, _25954_);
  or (_26735_, _26734_, _26730_);
  or (_26736_, _26735_, _25948_);
  nand (_26737_, _25716_, _26453_);
  or (_26738_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_26739_, _26738_, _26737_);
  and (_26740_, _26739_, _25890_);
  or (_26741_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_26742_, _25716_, _26528_);
  and (_26743_, _26742_, _26741_);
  and (_26744_, _26743_, _25954_);
  or (_26745_, _26744_, _26740_);
  or (_26746_, _26745_, _25800_);
  and (_26747_, _26746_, _25937_);
  and (_26748_, _26747_, _26736_);
  or (_26749_, _26748_, _26726_);
  or (_26750_, _26749_, _25947_);
  or (_26751_, _26004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_26752_, _26751_, _27053_);
  and (_00049_, _26752_, _26750_);
  and (_26753_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_26754_, _25716_, _26166_);
  or (_26755_, _26754_, _26753_);
  and (_26756_, _26755_, _25890_);
  nor (_26757_, _25716_, _26212_);
  and (_26758_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_26759_, _26758_, _26757_);
  and (_26760_, _26759_, _25954_);
  or (_26761_, _26760_, _26756_);
  or (_26762_, _26761_, _25948_);
  and (_26763_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_26764_, _25716_, _26261_);
  or (_26765_, _26764_, _26763_);
  and (_26766_, _26765_, _25890_);
  nor (_26767_, _25716_, _26312_);
  and (_26768_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_26769_, _26768_, _26767_);
  and (_26770_, _26769_, _25954_);
  or (_26771_, _26770_, _26766_);
  or (_26772_, _26771_, _25800_);
  and (_26773_, _26772_, _25962_);
  and (_26774_, _26773_, _26762_);
  nand (_26775_, _25716_, _26337_);
  or (_26776_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_26777_, _26776_, _26775_);
  and (_26778_, _26777_, _25890_);
  or (_26779_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_26780_, _25716_, _26383_);
  and (_26781_, _26780_, _26779_);
  and (_26782_, _26781_, _25954_);
  or (_26783_, _26782_, _26778_);
  or (_26784_, _26783_, _25948_);
  nand (_26785_, _25716_, _26456_);
  or (_26786_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_26787_, _26786_, _26785_);
  and (_26788_, _26787_, _25890_);
  or (_26789_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_26790_, _25716_, _26531_);
  and (_26791_, _26790_, _26789_);
  and (_26792_, _26791_, _25954_);
  or (_26793_, _26792_, _26788_);
  or (_26794_, _26793_, _25800_);
  and (_26795_, _26794_, _25937_);
  and (_26796_, _26795_, _26784_);
  or (_26797_, _26796_, _26774_);
  or (_26798_, _26797_, _25947_);
  or (_26799_, _26004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_26800_, _26799_, _27053_);
  and (_00051_, _26800_, _26798_);
  and (_26801_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_26802_, _25716_, _26555_);
  or (_26803_, _26802_, _26801_);
  or (_26804_, _26803_, _25890_);
  nand (_26805_, _25716_, _26459_);
  or (_26806_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and (_26807_, _26806_, _26805_);
  or (_26808_, _26807_, _25954_);
  and (_26809_, _26808_, _25937_);
  and (_26810_, _26809_, _26804_);
  and (_26811_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_26812_, _25955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_26813_, _26812_, _25954_);
  or (_26814_, _26813_, _26811_);
  nor (_26815_, _25716_, _26315_);
  and (_26816_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_26817_, _26816_, _25890_);
  or (_26818_, _26817_, _26815_);
  and (_26819_, _26818_, _25962_);
  and (_26820_, _26819_, _26814_);
  or (_26821_, _26820_, _26810_);
  and (_26822_, _26821_, _25948_);
  or (_26823_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_26824_, _25716_, _26386_);
  and (_26825_, _26824_, _26823_);
  or (_26826_, _26825_, _25890_);
  nand (_26827_, _25716_, _26340_);
  or (_26828_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_26829_, _26828_, _26827_);
  or (_26830_, _26829_, _25954_);
  and (_26831_, _26830_, _25937_);
  and (_26832_, _26831_, _26826_);
  and (_26833_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_26834_, _25716_, _26169_);
  or (_26835_, _26834_, _25954_);
  or (_26836_, _26835_, _26833_);
  and (_26837_, _25955_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_26838_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_26839_, _26838_, _25890_);
  or (_26840_, _26839_, _26837_);
  and (_26841_, _26840_, _25962_);
  and (_26842_, _26841_, _26836_);
  or (_26843_, _26842_, _26832_);
  and (_26844_, _26843_, _25800_);
  or (_26845_, _26844_, _25947_);
  or (_26846_, _26845_, _26822_);
  or (_26847_, _26004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_26848_, _26847_, _27053_);
  and (_00053_, _26848_, _26846_);
  and (_26849_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_26850_, _25716_, _26172_);
  or (_26851_, _26850_, _26849_);
  and (_26852_, _26851_, _25890_);
  nor (_26853_, _25716_, _26217_);
  and (_26854_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_26855_, _26854_, _26853_);
  and (_26856_, _26855_, _25954_);
  or (_26857_, _26856_, _26852_);
  or (_26858_, _26857_, _25948_);
  and (_26859_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_26860_, _25716_, _26268_);
  or (_26861_, _26860_, _26859_);
  and (_26862_, _26861_, _25890_);
  nor (_26863_, _25716_, _26318_);
  and (_26864_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_26865_, _26864_, _26863_);
  and (_26866_, _26865_, _25954_);
  or (_26867_, _26866_, _26862_);
  or (_26868_, _26867_, _25800_);
  and (_26869_, _26868_, _25962_);
  and (_26870_, _26869_, _26858_);
  nand (_26871_, _25716_, _26343_);
  or (_26872_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_26873_, _26872_, _26871_);
  and (_26874_, _26873_, _25890_);
  or (_26875_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_26876_, _25716_, _26393_);
  and (_26877_, _26876_, _26875_);
  and (_26878_, _26877_, _25954_);
  or (_26879_, _26878_, _26874_);
  or (_26880_, _26879_, _25948_);
  nand (_26881_, _25716_, _26463_);
  or (_26882_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_26883_, _26882_, _26881_);
  and (_26884_, _26883_, _25890_);
  or (_26885_, _25716_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_26886_, _25716_, _26536_);
  and (_26887_, _26886_, _26885_);
  and (_26888_, _26887_, _25954_);
  or (_26889_, _26888_, _26884_);
  or (_26890_, _26889_, _25800_);
  and (_26891_, _26890_, _25937_);
  and (_26892_, _26891_, _26880_);
  or (_26893_, _26892_, _26870_);
  or (_26894_, _26893_, _25947_);
  or (_26895_, _26004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_26896_, _26895_, _27053_);
  and (_00055_, _26896_, _26894_);
  or (_26897_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_26898_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_26899_, _26898_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_26900_, _26899_, _26897_);
  nand (_26901_, _26900_, _27053_);
  or (_26902_, \oc8051_gm_cxrom_1.cell0.data [7], _27053_);
  and (_00062_, _26902_, _26901_);
  or (_26903_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_26904_, \oc8051_gm_cxrom_1.cell0.data [0], _26898_);
  nand (_26905_, _26904_, _26903_);
  nand (_26906_, _26905_, _27053_);
  or (_26907_, \oc8051_gm_cxrom_1.cell0.data [0], _27053_);
  and (_00088_, _26907_, _26906_);
  or (_26908_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_26909_, \oc8051_gm_cxrom_1.cell0.data [1], _26898_);
  nand (_26910_, _26909_, _26908_);
  nand (_26911_, _26910_, _27053_);
  or (_26912_, \oc8051_gm_cxrom_1.cell0.data [1], _27053_);
  and (_00090_, _26912_, _26911_);
  or (_26913_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_26914_, \oc8051_gm_cxrom_1.cell0.data [2], _26898_);
  nand (_26915_, _26914_, _26913_);
  nand (_26916_, _26915_, _27053_);
  or (_26917_, \oc8051_gm_cxrom_1.cell0.data [2], _27053_);
  and (_00092_, _26917_, _26916_);
  or (_26918_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_26919_, \oc8051_gm_cxrom_1.cell0.data [3], _26898_);
  nand (_26920_, _26919_, _26918_);
  nand (_26921_, _26920_, _27053_);
  or (_26922_, \oc8051_gm_cxrom_1.cell0.data [3], _27053_);
  and (_00094_, _26922_, _26921_);
  or (_26923_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_26924_, \oc8051_gm_cxrom_1.cell0.data [4], _26898_);
  nand (_26925_, _26924_, _26923_);
  nand (_26926_, _26925_, _27053_);
  or (_26927_, \oc8051_gm_cxrom_1.cell0.data [4], _27053_);
  and (_00096_, _26927_, _26926_);
  or (_26928_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_26929_, \oc8051_gm_cxrom_1.cell0.data [5], _26898_);
  nand (_26930_, _26929_, _26928_);
  nand (_26931_, _26930_, _27053_);
  or (_26932_, \oc8051_gm_cxrom_1.cell0.data [5], _27053_);
  and (_00098_, _26932_, _26931_);
  or (_26933_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_26934_, \oc8051_gm_cxrom_1.cell0.data [6], _26898_);
  nand (_26935_, _26934_, _26933_);
  nand (_26936_, _26935_, _27053_);
  or (_26937_, \oc8051_gm_cxrom_1.cell0.data [6], _27053_);
  and (_00100_, _26937_, _26936_);
  or (_26938_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_26939_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_26940_, _26939_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_26941_, _26940_, _26938_);
  nand (_26942_, _26941_, _27053_);
  or (_26943_, \oc8051_gm_cxrom_1.cell1.data [7], _27053_);
  and (_00108_, _26943_, _26942_);
  or (_26944_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_26945_, \oc8051_gm_cxrom_1.cell1.data [0], _26939_);
  nand (_26946_, _26945_, _26944_);
  nand (_26947_, _26946_, _27053_);
  or (_26948_, \oc8051_gm_cxrom_1.cell1.data [0], _27053_);
  and (_00140_, _26948_, _26947_);
  or (_26949_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_26950_, \oc8051_gm_cxrom_1.cell1.data [1], _26939_);
  nand (_26951_, _26950_, _26949_);
  nand (_26952_, _26951_, _27053_);
  or (_26953_, \oc8051_gm_cxrom_1.cell1.data [1], _27053_);
  and (_00142_, _26953_, _26952_);
  or (_26954_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_26955_, \oc8051_gm_cxrom_1.cell1.data [2], _26939_);
  nand (_26956_, _26955_, _26954_);
  nand (_26957_, _26956_, _27053_);
  or (_26958_, \oc8051_gm_cxrom_1.cell1.data [2], _27053_);
  and (_00144_, _26958_, _26957_);
  or (_26959_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_26960_, \oc8051_gm_cxrom_1.cell1.data [3], _26939_);
  nand (_26961_, _26960_, _26959_);
  nand (_26962_, _26961_, _27053_);
  or (_26963_, \oc8051_gm_cxrom_1.cell1.data [3], _27053_);
  and (_00146_, _26963_, _26962_);
  or (_26964_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_26965_, \oc8051_gm_cxrom_1.cell1.data [4], _26939_);
  nand (_26966_, _26965_, _26964_);
  nand (_26967_, _26966_, _27053_);
  or (_26968_, \oc8051_gm_cxrom_1.cell1.data [4], _27053_);
  and (_00148_, _26968_, _26967_);
  or (_26969_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_26970_, \oc8051_gm_cxrom_1.cell1.data [5], _26939_);
  nand (_26971_, _26970_, _26969_);
  nand (_26972_, _26971_, _27053_);
  or (_26973_, \oc8051_gm_cxrom_1.cell1.data [5], _27053_);
  and (_00149_, _26973_, _26972_);
  or (_26974_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_26975_, \oc8051_gm_cxrom_1.cell1.data [6], _26939_);
  nand (_26976_, _26975_, _26974_);
  nand (_26977_, _26976_, _27053_);
  or (_26978_, \oc8051_gm_cxrom_1.cell1.data [6], _27053_);
  and (_00151_, _26978_, _26977_);
  or (_26979_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_26980_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_26981_, _26980_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_26982_, _26981_, _26979_);
  nand (_26983_, _26982_, _27053_);
  or (_26984_, \oc8051_gm_cxrom_1.cell2.data [7], _27053_);
  and (_00158_, _26984_, _26983_);
  or (_26985_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_26986_, \oc8051_gm_cxrom_1.cell2.data [0], _26980_);
  nand (_26987_, _26986_, _26985_);
  nand (_26988_, _26987_, _27053_);
  or (_26989_, \oc8051_gm_cxrom_1.cell2.data [0], _27053_);
  and (_00190_, _26989_, _26988_);
  or (_26990_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_26991_, \oc8051_gm_cxrom_1.cell2.data [1], _26980_);
  nand (_26992_, _26991_, _26990_);
  nand (_26993_, _26992_, _27053_);
  or (_26994_, \oc8051_gm_cxrom_1.cell2.data [1], _27053_);
  and (_00192_, _26994_, _26993_);
  or (_26995_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_26996_, \oc8051_gm_cxrom_1.cell2.data [2], _26980_);
  nand (_26997_, _26996_, _26995_);
  nand (_26998_, _26997_, _27053_);
  or (_26999_, \oc8051_gm_cxrom_1.cell2.data [2], _27053_);
  and (_00194_, _26999_, _26998_);
  or (_27000_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_27001_, \oc8051_gm_cxrom_1.cell2.data [3], _26980_);
  nand (_27002_, _27001_, _27000_);
  nand (_27003_, _27002_, _27053_);
  or (_27004_, \oc8051_gm_cxrom_1.cell2.data [3], _27053_);
  and (_00196_, _27004_, _27003_);
  or (_27005_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_27006_, \oc8051_gm_cxrom_1.cell2.data [4], _26980_);
  nand (_27007_, _27006_, _27005_);
  nand (_27008_, _27007_, _27053_);
  or (_27009_, \oc8051_gm_cxrom_1.cell2.data [4], _27053_);
  and (_00198_, _27009_, _27008_);
  or (_27010_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_27011_, \oc8051_gm_cxrom_1.cell2.data [5], _26980_);
  nand (_27012_, _27011_, _27010_);
  nand (_27013_, _27012_, _27053_);
  or (_27014_, \oc8051_gm_cxrom_1.cell2.data [5], _27053_);
  and (_00200_, _27014_, _27013_);
  or (_27015_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_27016_, \oc8051_gm_cxrom_1.cell2.data [6], _26980_);
  nand (_27017_, _27016_, _27015_);
  nand (_27018_, _27017_, _27053_);
  or (_27019_, \oc8051_gm_cxrom_1.cell2.data [6], _27053_);
  and (_00202_, _27019_, _27018_);
  or (_27020_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_27021_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_27022_, _27021_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_27023_, _27022_, _27020_);
  nand (_27024_, _27023_, _27053_);
  or (_27025_, \oc8051_gm_cxrom_1.cell3.data [7], _27053_);
  and (_00210_, _27025_, _27024_);
  or (_27026_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_27027_, \oc8051_gm_cxrom_1.cell3.data [0], _27021_);
  nand (_27028_, _27027_, _27026_);
  nand (_27029_, _27028_, _27053_);
  or (_27030_, \oc8051_gm_cxrom_1.cell3.data [0], _27053_);
  and (_00241_, _27030_, _27029_);
  or (_27031_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_27032_, \oc8051_gm_cxrom_1.cell3.data [1], _27021_);
  nand (_27033_, _27032_, _27031_);
  nand (_27034_, _27033_, _27053_);
  or (_27035_, \oc8051_gm_cxrom_1.cell3.data [1], _27053_);
  and (_00243_, _27035_, _27034_);
  or (_27036_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_27037_, \oc8051_gm_cxrom_1.cell3.data [2], _27021_);
  nand (_27038_, _27037_, _27036_);
  nand (_27039_, _27038_, _27053_);
  or (_27040_, \oc8051_gm_cxrom_1.cell3.data [2], _27053_);
  and (_00245_, _27040_, _27039_);
  or (_27041_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_27042_, \oc8051_gm_cxrom_1.cell3.data [3], _27021_);
  nand (_27043_, _27042_, _27041_);
  nand (_27044_, _27043_, _27053_);
  or (_27045_, \oc8051_gm_cxrom_1.cell3.data [3], _27053_);
  and (_00247_, _27045_, _27044_);
  or (_27046_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_27047_, \oc8051_gm_cxrom_1.cell3.data [4], _27021_);
  nand (_27048_, _27047_, _27046_);
  nand (_27049_, _27048_, _27053_);
  or (_27050_, \oc8051_gm_cxrom_1.cell3.data [4], _27053_);
  and (_00249_, _27050_, _27049_);
  or (_27051_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_27052_, \oc8051_gm_cxrom_1.cell3.data [5], _27021_);
  nand (_27054_, _27052_, _27051_);
  nand (_27055_, _27054_, _27053_);
  or (_27057_, \oc8051_gm_cxrom_1.cell3.data [5], _27053_);
  and (_00251_, _27057_, _27055_);
  or (_27059_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_27060_, \oc8051_gm_cxrom_1.cell3.data [6], _27021_);
  nand (_27062_, _27060_, _27059_);
  nand (_27063_, _27062_, _27053_);
  or (_27065_, \oc8051_gm_cxrom_1.cell3.data [6], _27053_);
  and (_00253_, _27065_, _27063_);
  or (_27067_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_27069_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_27071_, _27069_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_27072_, _27071_, _27067_);
  nand (_27073_, _27072_, _27053_);
  or (_27074_, \oc8051_gm_cxrom_1.cell4.data [7], _27053_);
  and (_00261_, _27074_, _27073_);
  or (_27075_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_27076_, \oc8051_gm_cxrom_1.cell4.data [0], _27069_);
  nand (_27077_, _27076_, _27075_);
  nand (_27078_, _27077_, _27053_);
  or (_27079_, \oc8051_gm_cxrom_1.cell4.data [0], _27053_);
  and (_00292_, _27079_, _27078_);
  or (_27080_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_27081_, \oc8051_gm_cxrom_1.cell4.data [1], _27069_);
  nand (_27082_, _27081_, _27080_);
  nand (_27083_, _27082_, _27053_);
  or (_27084_, \oc8051_gm_cxrom_1.cell4.data [1], _27053_);
  and (_00294_, _27084_, _27083_);
  or (_27085_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_27086_, \oc8051_gm_cxrom_1.cell4.data [2], _27069_);
  nand (_27087_, _27086_, _27085_);
  nand (_27088_, _27087_, _27053_);
  or (_27089_, \oc8051_gm_cxrom_1.cell4.data [2], _27053_);
  and (_00296_, _27089_, _27088_);
  or (_27090_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_27091_, \oc8051_gm_cxrom_1.cell4.data [3], _27069_);
  nand (_27092_, _27091_, _27090_);
  nand (_27093_, _27092_, _27053_);
  or (_27094_, \oc8051_gm_cxrom_1.cell4.data [3], _27053_);
  and (_00298_, _27094_, _27093_);
  or (_27095_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_27096_, \oc8051_gm_cxrom_1.cell4.data [4], _27069_);
  nand (_27097_, _27096_, _27095_);
  nand (_27098_, _27097_, _27053_);
  or (_27099_, \oc8051_gm_cxrom_1.cell4.data [4], _27053_);
  and (_00300_, _27099_, _27098_);
  or (_27100_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_27101_, \oc8051_gm_cxrom_1.cell4.data [5], _27069_);
  nand (_27102_, _27101_, _27100_);
  nand (_27103_, _27102_, _27053_);
  or (_27104_, \oc8051_gm_cxrom_1.cell4.data [5], _27053_);
  and (_00302_, _27104_, _27103_);
  or (_27106_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_27108_, \oc8051_gm_cxrom_1.cell4.data [6], _27069_);
  nand (_27110_, _27108_, _27106_);
  nand (_27112_, _27110_, _27053_);
  or (_27114_, \oc8051_gm_cxrom_1.cell4.data [6], _27053_);
  and (_00304_, _27114_, _27112_);
  or (_27116_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_27118_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_27119_, _27118_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_27120_, _27119_, _27116_);
  nand (_27121_, _27120_, _27053_);
  or (_27122_, \oc8051_gm_cxrom_1.cell5.data [7], _27053_);
  and (_00312_, _27122_, _27121_);
  or (_27123_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_27124_, \oc8051_gm_cxrom_1.cell5.data [0], _27118_);
  nand (_27125_, _27124_, _27123_);
  nand (_27126_, _27125_, _27053_);
  or (_27127_, \oc8051_gm_cxrom_1.cell5.data [0], _27053_);
  and (_00343_, _27127_, _27126_);
  or (_27128_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_27129_, \oc8051_gm_cxrom_1.cell5.data [1], _27118_);
  nand (_27130_, _27129_, _27128_);
  nand (_27131_, _27130_, _27053_);
  or (_27132_, \oc8051_gm_cxrom_1.cell5.data [1], _27053_);
  and (_00345_, _27132_, _27131_);
  or (_27133_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_27134_, \oc8051_gm_cxrom_1.cell5.data [2], _27118_);
  nand (_27135_, _27134_, _27133_);
  nand (_27136_, _27135_, _27053_);
  or (_27137_, \oc8051_gm_cxrom_1.cell5.data [2], _27053_);
  and (_00347_, _27137_, _27136_);
  or (_27138_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_27139_, \oc8051_gm_cxrom_1.cell5.data [3], _27118_);
  nand (_27140_, _27139_, _27138_);
  nand (_27141_, _27140_, _27053_);
  or (_27142_, \oc8051_gm_cxrom_1.cell5.data [3], _27053_);
  and (_00349_, _27142_, _27141_);
  or (_27143_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_27144_, \oc8051_gm_cxrom_1.cell5.data [4], _27118_);
  nand (_27145_, _27144_, _27143_);
  nand (_27146_, _27145_, _27053_);
  or (_27147_, \oc8051_gm_cxrom_1.cell5.data [4], _27053_);
  and (_00351_, _27147_, _27146_);
  or (_27148_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_27149_, \oc8051_gm_cxrom_1.cell5.data [5], _27118_);
  nand (_27150_, _27149_, _27148_);
  nand (_27151_, _27150_, _27053_);
  or (_27152_, \oc8051_gm_cxrom_1.cell5.data [5], _27053_);
  and (_00352_, _27152_, _27151_);
  or (_27153_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_27154_, \oc8051_gm_cxrom_1.cell5.data [6], _27118_);
  nand (_27155_, _27154_, _27153_);
  nand (_27156_, _27155_, _27053_);
  or (_27157_, \oc8051_gm_cxrom_1.cell5.data [6], _27053_);
  and (_00354_, _27157_, _27156_);
  or (_27158_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_27159_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_27160_, _27159_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_27161_, _27160_, _27158_);
  nand (_27162_, _27161_, _27053_);
  or (_27163_, \oc8051_gm_cxrom_1.cell6.data [7], _27053_);
  and (_00362_, _27163_, _27162_);
  or (_27164_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_27165_, \oc8051_gm_cxrom_1.cell6.data [0], _27159_);
  nand (_27166_, _27165_, _27164_);
  nand (_27167_, _27166_, _27053_);
  or (_27168_, \oc8051_gm_cxrom_1.cell6.data [0], _27053_);
  and (_00395_, _27168_, _27167_);
  or (_27169_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_27170_, \oc8051_gm_cxrom_1.cell6.data [1], _27159_);
  nand (_27171_, _27170_, _27169_);
  nand (_27172_, _27171_, _27053_);
  or (_27173_, \oc8051_gm_cxrom_1.cell6.data [1], _27053_);
  and (_00397_, _27173_, _27172_);
  or (_27174_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_27175_, \oc8051_gm_cxrom_1.cell6.data [2], _27159_);
  nand (_27176_, _27175_, _27174_);
  nand (_27177_, _27176_, _27053_);
  or (_27178_, \oc8051_gm_cxrom_1.cell6.data [2], _27053_);
  and (_00399_, _27178_, _27177_);
  or (_27179_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_27180_, \oc8051_gm_cxrom_1.cell6.data [3], _27159_);
  nand (_27181_, _27180_, _27179_);
  nand (_27182_, _27181_, _27053_);
  or (_27183_, \oc8051_gm_cxrom_1.cell6.data [3], _27053_);
  and (_00401_, _27183_, _27182_);
  or (_27184_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_27185_, \oc8051_gm_cxrom_1.cell6.data [4], _27159_);
  nand (_27186_, _27185_, _27184_);
  nand (_27187_, _27186_, _27053_);
  or (_27188_, \oc8051_gm_cxrom_1.cell6.data [4], _27053_);
  and (_00403_, _27188_, _27187_);
  or (_27189_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_27190_, \oc8051_gm_cxrom_1.cell6.data [5], _27159_);
  nand (_27191_, _27190_, _27189_);
  nand (_27192_, _27191_, _27053_);
  or (_27193_, \oc8051_gm_cxrom_1.cell6.data [5], _27053_);
  and (_00405_, _27193_, _27192_);
  or (_27194_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_27195_, \oc8051_gm_cxrom_1.cell6.data [6], _27159_);
  nand (_27196_, _27195_, _27194_);
  nand (_27197_, _27196_, _27053_);
  or (_27198_, \oc8051_gm_cxrom_1.cell6.data [6], _27053_);
  and (_00407_, _27198_, _27197_);
  or (_27199_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_27200_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_27201_, _27200_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_27202_, _27201_, _27199_);
  nand (_27203_, _27202_, _27053_);
  or (_27204_, \oc8051_gm_cxrom_1.cell7.data [7], _27053_);
  and (_00415_, _27204_, _27203_);
  or (_27205_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_27206_, \oc8051_gm_cxrom_1.cell7.data [0], _27200_);
  nand (_27207_, _27206_, _27205_);
  nand (_27208_, _27207_, _27053_);
  or (_27209_, \oc8051_gm_cxrom_1.cell7.data [0], _27053_);
  and (_00448_, _27209_, _27208_);
  or (_27210_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_27211_, \oc8051_gm_cxrom_1.cell7.data [1], _27200_);
  nand (_27212_, _27211_, _27210_);
  nand (_27213_, _27212_, _27053_);
  or (_27214_, \oc8051_gm_cxrom_1.cell7.data [1], _27053_);
  and (_00450_, _27214_, _27213_);
  or (_27215_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_27216_, \oc8051_gm_cxrom_1.cell7.data [2], _27200_);
  nand (_27217_, _27216_, _27215_);
  nand (_27218_, _27217_, _27053_);
  or (_27219_, \oc8051_gm_cxrom_1.cell7.data [2], _27053_);
  and (_00452_, _27219_, _27218_);
  or (_27220_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_27221_, \oc8051_gm_cxrom_1.cell7.data [3], _27200_);
  nand (_27222_, _27221_, _27220_);
  nand (_27223_, _27222_, _27053_);
  or (_27224_, \oc8051_gm_cxrom_1.cell7.data [3], _27053_);
  and (_00454_, _27224_, _27223_);
  or (_27225_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_27226_, \oc8051_gm_cxrom_1.cell7.data [4], _27200_);
  nand (_27227_, _27226_, _27225_);
  nand (_27228_, _27227_, _27053_);
  or (_27229_, \oc8051_gm_cxrom_1.cell7.data [4], _27053_);
  and (_00456_, _27229_, _27228_);
  or (_27230_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_27231_, \oc8051_gm_cxrom_1.cell7.data [5], _27200_);
  nand (_27232_, _27231_, _27230_);
  nand (_27233_, _27232_, _27053_);
  or (_27234_, \oc8051_gm_cxrom_1.cell7.data [5], _27053_);
  and (_00458_, _27234_, _27233_);
  or (_27235_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_27236_, \oc8051_gm_cxrom_1.cell7.data [6], _27200_);
  nand (_27237_, _27236_, _27235_);
  nand (_27238_, _27237_, _27053_);
  or (_27239_, \oc8051_gm_cxrom_1.cell7.data [6], _27053_);
  and (_00460_, _27239_, _27238_);
  or (_27240_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_27241_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_27242_, _27241_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_27243_, _27242_, _27240_);
  nand (_27244_, _27243_, _27053_);
  or (_27245_, \oc8051_gm_cxrom_1.cell8.data [7], _27053_);
  and (_00467_, _27245_, _27244_);
  or (_27246_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_27247_, \oc8051_gm_cxrom_1.cell8.data [0], _27241_);
  nand (_27248_, _27247_, _27246_);
  nand (_27249_, _27248_, _27053_);
  or (_27250_, \oc8051_gm_cxrom_1.cell8.data [0], _27053_);
  and (_00499_, _27250_, _27249_);
  or (_27251_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_27252_, \oc8051_gm_cxrom_1.cell8.data [1], _27241_);
  nand (_27253_, _27252_, _27251_);
  nand (_27254_, _27253_, _27053_);
  or (_27255_, \oc8051_gm_cxrom_1.cell8.data [1], _27053_);
  and (_00501_, _27255_, _27254_);
  or (_27256_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_27257_, \oc8051_gm_cxrom_1.cell8.data [2], _27241_);
  nand (_27258_, _27257_, _27256_);
  nand (_27259_, _27258_, _27053_);
  or (_27260_, \oc8051_gm_cxrom_1.cell8.data [2], _27053_);
  and (_00503_, _27260_, _27259_);
  or (_27261_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_27262_, \oc8051_gm_cxrom_1.cell8.data [3], _27241_);
  nand (_27263_, _27262_, _27261_);
  nand (_27264_, _27263_, _27053_);
  or (_27265_, \oc8051_gm_cxrom_1.cell8.data [3], _27053_);
  and (_00505_, _27265_, _27264_);
  or (_27266_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_27267_, \oc8051_gm_cxrom_1.cell8.data [4], _27241_);
  nand (_27268_, _27267_, _27266_);
  nand (_27269_, _27268_, _27053_);
  or (_27270_, \oc8051_gm_cxrom_1.cell8.data [4], _27053_);
  and (_00507_, _27270_, _27269_);
  or (_27271_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_27272_, \oc8051_gm_cxrom_1.cell8.data [5], _27241_);
  nand (_27273_, _27272_, _27271_);
  nand (_27274_, _27273_, _27053_);
  or (_27275_, \oc8051_gm_cxrom_1.cell8.data [5], _27053_);
  and (_00509_, _27275_, _27274_);
  or (_27276_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_27277_, \oc8051_gm_cxrom_1.cell8.data [6], _27241_);
  nand (_27278_, _27277_, _27276_);
  nand (_27279_, _27278_, _27053_);
  or (_27280_, \oc8051_gm_cxrom_1.cell8.data [6], _27053_);
  and (_00511_, _27280_, _27279_);
  or (_27281_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_27282_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_27283_, _27282_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_27284_, _27283_, _27281_);
  nand (_27285_, _27284_, _27053_);
  or (_27286_, \oc8051_gm_cxrom_1.cell9.data [7], _27053_);
  and (_00519_, _27286_, _27285_);
  or (_27287_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_27288_, \oc8051_gm_cxrom_1.cell9.data [0], _27282_);
  nand (_27289_, _27288_, _27287_);
  nand (_27290_, _27289_, _27053_);
  or (_27291_, \oc8051_gm_cxrom_1.cell9.data [0], _27053_);
  and (_00551_, _27291_, _27290_);
  or (_27292_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_27293_, \oc8051_gm_cxrom_1.cell9.data [1], _27282_);
  nand (_27294_, _27293_, _27292_);
  nand (_27295_, _27294_, _27053_);
  or (_27296_, \oc8051_gm_cxrom_1.cell9.data [1], _27053_);
  and (_00553_, _27296_, _27295_);
  or (_27297_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_27298_, \oc8051_gm_cxrom_1.cell9.data [2], _27282_);
  nand (_27299_, _27298_, _27297_);
  nand (_27300_, _27299_, _27053_);
  or (_27301_, \oc8051_gm_cxrom_1.cell9.data [2], _27053_);
  and (_00555_, _27301_, _27300_);
  or (_27302_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_27303_, \oc8051_gm_cxrom_1.cell9.data [3], _27282_);
  nand (_27304_, _27303_, _27302_);
  nand (_27305_, _27304_, _27053_);
  or (_27306_, \oc8051_gm_cxrom_1.cell9.data [3], _27053_);
  and (_00557_, _27306_, _27305_);
  or (_27307_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_27308_, \oc8051_gm_cxrom_1.cell9.data [4], _27282_);
  nand (_27309_, _27308_, _27307_);
  nand (_27310_, _27309_, _27053_);
  or (_27311_, \oc8051_gm_cxrom_1.cell9.data [4], _27053_);
  and (_00559_, _27311_, _27310_);
  or (_27312_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_27313_, \oc8051_gm_cxrom_1.cell9.data [5], _27282_);
  nand (_27314_, _27313_, _27312_);
  nand (_27315_, _27314_, _27053_);
  or (_27316_, \oc8051_gm_cxrom_1.cell9.data [5], _27053_);
  and (_00561_, _27316_, _27315_);
  or (_27317_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_27318_, \oc8051_gm_cxrom_1.cell9.data [6], _27282_);
  nand (_27319_, _27318_, _27317_);
  nand (_27320_, _27319_, _27053_);
  or (_27321_, \oc8051_gm_cxrom_1.cell9.data [6], _27053_);
  and (_00563_, _27321_, _27320_);
  or (_27322_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_27323_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_27324_, _27323_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_27325_, _27324_, _27322_);
  nand (_27326_, _27325_, _27053_);
  or (_27327_, \oc8051_gm_cxrom_1.cell10.data [7], _27053_);
  and (_00571_, _27327_, _27326_);
  or (_27328_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_27329_, \oc8051_gm_cxrom_1.cell10.data [0], _27323_);
  nand (_27330_, _27329_, _27328_);
  nand (_27331_, _27330_, _27053_);
  or (_27332_, \oc8051_gm_cxrom_1.cell10.data [0], _27053_);
  and (_00603_, _27332_, _27331_);
  or (_27333_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_27334_, \oc8051_gm_cxrom_1.cell10.data [1], _27323_);
  nand (_27335_, _27334_, _27333_);
  nand (_27336_, _27335_, _27053_);
  or (_27337_, \oc8051_gm_cxrom_1.cell10.data [1], _27053_);
  and (_00605_, _27337_, _27336_);
  or (_27338_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_27339_, \oc8051_gm_cxrom_1.cell10.data [2], _27323_);
  nand (_27340_, _27339_, _27338_);
  nand (_27341_, _27340_, _27053_);
  or (_27342_, \oc8051_gm_cxrom_1.cell10.data [2], _27053_);
  and (_00607_, _27342_, _27341_);
  or (_27343_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_27344_, \oc8051_gm_cxrom_1.cell10.data [3], _27323_);
  nand (_27345_, _27344_, _27343_);
  nand (_27346_, _27345_, _27053_);
  or (_27347_, \oc8051_gm_cxrom_1.cell10.data [3], _27053_);
  and (_00609_, _27347_, _27346_);
  or (_27348_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_27349_, \oc8051_gm_cxrom_1.cell10.data [4], _27323_);
  nand (_27350_, _27349_, _27348_);
  nand (_27351_, _27350_, _27053_);
  or (_27352_, \oc8051_gm_cxrom_1.cell10.data [4], _27053_);
  and (_00611_, _27352_, _27351_);
  or (_27353_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_27354_, \oc8051_gm_cxrom_1.cell10.data [5], _27323_);
  nand (_27355_, _27354_, _27353_);
  nand (_27356_, _27355_, _27053_);
  or (_27357_, \oc8051_gm_cxrom_1.cell10.data [5], _27053_);
  and (_00613_, _27357_, _27356_);
  or (_27358_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_27359_, \oc8051_gm_cxrom_1.cell10.data [6], _27323_);
  nand (_27360_, _27359_, _27358_);
  nand (_27361_, _27360_, _27053_);
  or (_27362_, \oc8051_gm_cxrom_1.cell10.data [6], _27053_);
  and (_00615_, _27362_, _27361_);
  or (_27363_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_27364_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_27365_, _27364_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_27366_, _27365_, _27363_);
  nand (_27367_, _27366_, _27053_);
  or (_27368_, \oc8051_gm_cxrom_1.cell11.data [7], _27053_);
  and (_00623_, _27368_, _27367_);
  or (_27369_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_27370_, \oc8051_gm_cxrom_1.cell11.data [0], _27364_);
  nand (_27371_, _27370_, _27369_);
  nand (_27372_, _27371_, _27053_);
  or (_27373_, \oc8051_gm_cxrom_1.cell11.data [0], _27053_);
  and (_00655_, _27373_, _27372_);
  or (_27374_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_27375_, \oc8051_gm_cxrom_1.cell11.data [1], _27364_);
  nand (_27376_, _27375_, _27374_);
  nand (_27377_, _27376_, _27053_);
  or (_27378_, \oc8051_gm_cxrom_1.cell11.data [1], _27053_);
  and (_00657_, _27378_, _27377_);
  or (_27379_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_27380_, \oc8051_gm_cxrom_1.cell11.data [2], _27364_);
  nand (_27381_, _27380_, _27379_);
  nand (_27382_, _27381_, _27053_);
  or (_27383_, \oc8051_gm_cxrom_1.cell11.data [2], _27053_);
  and (_00659_, _27383_, _27382_);
  or (_27384_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_27385_, \oc8051_gm_cxrom_1.cell11.data [3], _27364_);
  nand (_27386_, _27385_, _27384_);
  nand (_27387_, _27386_, _27053_);
  or (_27388_, \oc8051_gm_cxrom_1.cell11.data [3], _27053_);
  and (_00661_, _27388_, _27387_);
  or (_27389_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_27390_, \oc8051_gm_cxrom_1.cell11.data [4], _27364_);
  nand (_27391_, _27390_, _27389_);
  nand (_27392_, _27391_, _27053_);
  or (_27393_, \oc8051_gm_cxrom_1.cell11.data [4], _27053_);
  and (_00663_, _27393_, _27392_);
  or (_27394_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_27395_, \oc8051_gm_cxrom_1.cell11.data [5], _27364_);
  nand (_27396_, _27395_, _27394_);
  nand (_27397_, _27396_, _27053_);
  or (_27398_, \oc8051_gm_cxrom_1.cell11.data [5], _27053_);
  and (_00665_, _27398_, _27397_);
  or (_27399_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_27400_, \oc8051_gm_cxrom_1.cell11.data [6], _27364_);
  nand (_27401_, _27400_, _27399_);
  nand (_27402_, _27401_, _27053_);
  or (_27403_, \oc8051_gm_cxrom_1.cell11.data [6], _27053_);
  and (_00667_, _27403_, _27402_);
  or (_27404_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_27405_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_27406_, _27405_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_27407_, _27406_, _27404_);
  nand (_27408_, _27407_, _27053_);
  or (_27409_, \oc8051_gm_cxrom_1.cell12.data [7], _27053_);
  and (_00675_, _27409_, _27408_);
  or (_27410_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_27411_, \oc8051_gm_cxrom_1.cell12.data [0], _27405_);
  nand (_27412_, _27411_, _27410_);
  nand (_27413_, _27412_, _27053_);
  or (_27414_, \oc8051_gm_cxrom_1.cell12.data [0], _27053_);
  and (_00707_, _27414_, _27413_);
  or (_27415_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_27416_, \oc8051_gm_cxrom_1.cell12.data [1], _27405_);
  nand (_27417_, _27416_, _27415_);
  nand (_27418_, _27417_, _27053_);
  or (_27419_, \oc8051_gm_cxrom_1.cell12.data [1], _27053_);
  and (_00709_, _27419_, _27418_);
  or (_27420_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_27421_, \oc8051_gm_cxrom_1.cell12.data [2], _27405_);
  nand (_27422_, _27421_, _27420_);
  nand (_27423_, _27422_, _27053_);
  or (_27424_, \oc8051_gm_cxrom_1.cell12.data [2], _27053_);
  and (_00711_, _27424_, _27423_);
  or (_27425_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_27426_, \oc8051_gm_cxrom_1.cell12.data [3], _27405_);
  nand (_27427_, _27426_, _27425_);
  nand (_27428_, _27427_, _27053_);
  or (_27429_, \oc8051_gm_cxrom_1.cell12.data [3], _27053_);
  and (_00713_, _27429_, _27428_);
  or (_27430_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_27431_, \oc8051_gm_cxrom_1.cell12.data [4], _27405_);
  nand (_27432_, _27431_, _27430_);
  nand (_27433_, _27432_, _27053_);
  or (_27434_, \oc8051_gm_cxrom_1.cell12.data [4], _27053_);
  and (_00715_, _27434_, _27433_);
  or (_27435_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_27436_, \oc8051_gm_cxrom_1.cell12.data [5], _27405_);
  nand (_27437_, _27436_, _27435_);
  nand (_27438_, _27437_, _27053_);
  or (_27439_, \oc8051_gm_cxrom_1.cell12.data [5], _27053_);
  and (_00717_, _27439_, _27438_);
  or (_27440_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_27441_, \oc8051_gm_cxrom_1.cell12.data [6], _27405_);
  nand (_27442_, _27441_, _27440_);
  nand (_27443_, _27442_, _27053_);
  or (_27444_, \oc8051_gm_cxrom_1.cell12.data [6], _27053_);
  and (_00719_, _27444_, _27443_);
  or (_27445_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_27446_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_27447_, _27446_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_27448_, _27447_, _27445_);
  nand (_27449_, _27448_, _27053_);
  or (_27450_, \oc8051_gm_cxrom_1.cell13.data [7], _27053_);
  and (_00727_, _27450_, _27449_);
  or (_27451_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_27452_, \oc8051_gm_cxrom_1.cell13.data [0], _27446_);
  nand (_27453_, _27452_, _27451_);
  nand (_27454_, _27453_, _27053_);
  or (_27455_, \oc8051_gm_cxrom_1.cell13.data [0], _27053_);
  and (_00759_, _27455_, _27454_);
  or (_27456_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_27457_, \oc8051_gm_cxrom_1.cell13.data [1], _27446_);
  nand (_27458_, _27457_, _27456_);
  nand (_27459_, _27458_, _27053_);
  or (_27460_, \oc8051_gm_cxrom_1.cell13.data [1], _27053_);
  and (_00761_, _27460_, _27459_);
  or (_27461_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_27462_, \oc8051_gm_cxrom_1.cell13.data [2], _27446_);
  nand (_27463_, _27462_, _27461_);
  nand (_27464_, _27463_, _27053_);
  or (_27465_, \oc8051_gm_cxrom_1.cell13.data [2], _27053_);
  and (_00763_, _27465_, _27464_);
  or (_27466_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_27467_, \oc8051_gm_cxrom_1.cell13.data [3], _27446_);
  nand (_27468_, _27467_, _27466_);
  nand (_27469_, _27468_, _27053_);
  or (_27470_, \oc8051_gm_cxrom_1.cell13.data [3], _27053_);
  and (_00765_, _27470_, _27469_);
  or (_27471_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_27472_, \oc8051_gm_cxrom_1.cell13.data [4], _27446_);
  nand (_27473_, _27472_, _27471_);
  nand (_27474_, _27473_, _27053_);
  or (_27475_, \oc8051_gm_cxrom_1.cell13.data [4], _27053_);
  and (_00767_, _27475_, _27474_);
  or (_27476_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_27477_, \oc8051_gm_cxrom_1.cell13.data [5], _27446_);
  nand (_27478_, _27477_, _27476_);
  nand (_27479_, _27478_, _27053_);
  or (_27480_, \oc8051_gm_cxrom_1.cell13.data [5], _27053_);
  and (_00769_, _27480_, _27479_);
  or (_27481_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_27482_, \oc8051_gm_cxrom_1.cell13.data [6], _27446_);
  nand (_27483_, _27482_, _27481_);
  nand (_27484_, _27483_, _27053_);
  or (_27485_, \oc8051_gm_cxrom_1.cell13.data [6], _27053_);
  and (_00771_, _27485_, _27484_);
  or (_27486_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_27487_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_27488_, _27487_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_27489_, _27488_, _27486_);
  nand (_27490_, _27489_, _27053_);
  or (_27491_, \oc8051_gm_cxrom_1.cell14.data [7], _27053_);
  and (_00779_, _27491_, _27490_);
  or (_27492_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_27493_, \oc8051_gm_cxrom_1.cell14.data [0], _27487_);
  nand (_27494_, _27493_, _27492_);
  nand (_27495_, _27494_, _27053_);
  or (_27496_, \oc8051_gm_cxrom_1.cell14.data [0], _27053_);
  and (_00811_, _27496_, _27495_);
  or (_27497_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_27498_, \oc8051_gm_cxrom_1.cell14.data [1], _27487_);
  nand (_27499_, _27498_, _27497_);
  nand (_27500_, _27499_, _27053_);
  or (_27501_, \oc8051_gm_cxrom_1.cell14.data [1], _27053_);
  and (_00813_, _27501_, _27500_);
  or (_27502_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_27503_, \oc8051_gm_cxrom_1.cell14.data [2], _27487_);
  nand (_27504_, _27503_, _27502_);
  nand (_27505_, _27504_, _27053_);
  or (_27506_, \oc8051_gm_cxrom_1.cell14.data [2], _27053_);
  and (_00815_, _27506_, _27505_);
  or (_27507_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_27508_, \oc8051_gm_cxrom_1.cell14.data [3], _27487_);
  nand (_27509_, _27508_, _27507_);
  nand (_27510_, _27509_, _27053_);
  or (_27511_, \oc8051_gm_cxrom_1.cell14.data [3], _27053_);
  and (_00817_, _27511_, _27510_);
  or (_27512_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_27513_, \oc8051_gm_cxrom_1.cell14.data [4], _27487_);
  nand (_27514_, _27513_, _27512_);
  nand (_27515_, _27514_, _27053_);
  or (_27516_, \oc8051_gm_cxrom_1.cell14.data [4], _27053_);
  and (_00819_, _27516_, _27515_);
  or (_27517_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_27518_, \oc8051_gm_cxrom_1.cell14.data [5], _27487_);
  nand (_27519_, _27518_, _27517_);
  nand (_27520_, _27519_, _27053_);
  or (_27521_, \oc8051_gm_cxrom_1.cell14.data [5], _27053_);
  and (_00821_, _27521_, _27520_);
  or (_27522_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_27523_, \oc8051_gm_cxrom_1.cell14.data [6], _27487_);
  nand (_27524_, _27523_, _27522_);
  nand (_27525_, _27524_, _27053_);
  or (_27526_, \oc8051_gm_cxrom_1.cell14.data [6], _27053_);
  and (_00823_, _27526_, _27525_);
  or (_27527_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_27528_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_27529_, _27528_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_27530_, _27529_, _27527_);
  nand (_27531_, _27530_, _27053_);
  or (_27532_, \oc8051_gm_cxrom_1.cell15.data [7], _27053_);
  and (_00831_, _27532_, _27531_);
  or (_27533_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_27534_, \oc8051_gm_cxrom_1.cell15.data [0], _27528_);
  nand (_27535_, _27534_, _27533_);
  nand (_27536_, _27535_, _27053_);
  or (_27537_, \oc8051_gm_cxrom_1.cell15.data [0], _27053_);
  and (_00863_, _27537_, _27536_);
  or (_27538_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_27539_, \oc8051_gm_cxrom_1.cell15.data [1], _27528_);
  nand (_27540_, _27539_, _27538_);
  nand (_27541_, _27540_, _27053_);
  or (_27542_, \oc8051_gm_cxrom_1.cell15.data [1], _27053_);
  and (_00865_, _27542_, _27541_);
  or (_27543_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_27544_, \oc8051_gm_cxrom_1.cell15.data [2], _27528_);
  nand (_27545_, _27544_, _27543_);
  nand (_27546_, _27545_, _27053_);
  or (_27547_, \oc8051_gm_cxrom_1.cell15.data [2], _27053_);
  and (_00867_, _27547_, _27546_);
  or (_27548_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_27549_, \oc8051_gm_cxrom_1.cell15.data [3], _27528_);
  nand (_27550_, _27549_, _27548_);
  nand (_27551_, _27550_, _27053_);
  or (_27552_, \oc8051_gm_cxrom_1.cell15.data [3], _27053_);
  and (_00869_, _27552_, _27551_);
  or (_27553_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_27554_, \oc8051_gm_cxrom_1.cell15.data [4], _27528_);
  nand (_27555_, _27554_, _27553_);
  nand (_27556_, _27555_, _27053_);
  or (_27557_, \oc8051_gm_cxrom_1.cell15.data [4], _27053_);
  and (_00871_, _27557_, _27556_);
  or (_27558_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_27559_, \oc8051_gm_cxrom_1.cell15.data [5], _27528_);
  nand (_27560_, _27559_, _27558_);
  nand (_27561_, _27560_, _27053_);
  or (_27562_, \oc8051_gm_cxrom_1.cell15.data [5], _27053_);
  and (_00873_, _27562_, _27561_);
  or (_27563_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_27564_, \oc8051_gm_cxrom_1.cell15.data [6], _27528_);
  nand (_27565_, _27564_, _27563_);
  nand (_27566_, _27565_, _27053_);
  or (_27567_, \oc8051_gm_cxrom_1.cell15.data [6], _27053_);
  and (_00875_, _27567_, _27566_);
  nor (_00906_, _21576_, rst);
  nor (_00910_, _25577_, rst);
  and (_27568_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and (_27569_, _19975_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_27570_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_27571_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_27572_, _27571_, _27570_);
  and (_27573_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_27574_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_27575_, _27574_, _27573_);
  and (_27576_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_27577_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_27578_, _27577_, _27576_);
  and (_27579_, _27578_, _27575_);
  and (_27580_, _27579_, _27572_);
  nor (_27581_, _27580_, _19975_);
  nor (_27582_, _27581_, _27569_);
  nor (_27583_, _27582_, _25561_);
  nor (_27584_, _27583_, _27568_);
  nor (_00914_, _27584_, rst);
  nor (_01036_, _20293_, rst);
  and (_01039_, _20567_, _27053_);
  nor (_01042_, _20819_, rst);
  nor (_01044_, _21061_, rst);
  and (_01047_, _21850_, _27053_);
  nor (_01050_, _22091_, rst);
  nor (_01053_, _21335_, rst);
  nor (_01056_, _25709_, rst);
  nor (_01059_, _25866_, rst);
  nor (_01062_, _25793_, rst);
  nor (_01065_, _25671_, rst);
  nor (_01068_, _25828_, rst);
  nor (_01071_, _25756_, rst);
  nor (_01074_, _25914_, rst);
  and (_27585_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and (_27586_, _19975_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_27587_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_27588_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_27589_, _27588_, _27587_);
  and (_27590_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_27591_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_27592_, _27591_, _27590_);
  and (_27593_, _27592_, _27589_);
  and (_27594_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_27595_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_27596_, _27595_, _27594_);
  and (_27597_, _27596_, _27593_);
  nor (_27598_, _27597_, _19975_);
  nor (_27599_, _27598_, _27586_);
  nor (_27600_, _27599_, _25561_);
  nor (_27601_, _27600_, _27585_);
  nor (_01077_, _27601_, rst);
  and (_27602_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and (_27603_, _19975_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_27604_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_27605_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_27606_, _27605_, _27604_);
  and (_27607_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_27608_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_27609_, _27608_, _27607_);
  and (_27610_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_27611_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_27612_, _27611_, _27610_);
  and (_27613_, _27612_, _27609_);
  and (_27614_, _27613_, _27606_);
  nor (_27615_, _27614_, _19975_);
  nor (_27616_, _27615_, _27603_);
  nor (_27617_, _27616_, _25561_);
  nor (_27618_, _27617_, _27602_);
  nor (_01080_, _27618_, rst);
  and (_27619_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and (_27620_, _19975_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_27621_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_27622_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_27623_, _27622_, _27621_);
  and (_27624_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_27625_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_27626_, _27625_, _27624_);
  and (_27627_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_27628_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_27629_, _27628_, _27627_);
  and (_27630_, _27629_, _27626_);
  and (_27631_, _27630_, _27623_);
  nor (_27632_, _27631_, _19975_);
  nor (_27633_, _27632_, _27620_);
  nor (_27634_, _27633_, _25561_);
  nor (_27635_, _27634_, _27619_);
  nor (_01083_, _27635_, rst);
  and (_27636_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and (_27637_, _19975_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_27638_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_27639_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_27640_, _27639_, _27638_);
  and (_27641_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_27642_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_27643_, _27642_, _27641_);
  and (_27644_, _27643_, _27640_);
  and (_27645_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_27646_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_27647_, _27646_, _27645_);
  and (_27648_, _27647_, _27644_);
  nor (_27649_, _27648_, _19975_);
  nor (_27650_, _27649_, _27637_);
  nor (_27651_, _27650_, _25561_);
  nor (_27652_, _27651_, _27636_);
  nor (_01086_, _27652_, rst);
  and (_27653_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and (_27654_, _19975_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_27655_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_27656_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_27657_, _27656_, _27655_);
  and (_27658_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_27659_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_27660_, _27659_, _27658_);
  and (_27661_, _27660_, _27657_);
  and (_27662_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_27663_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_27664_, _27663_, _27662_);
  and (_27665_, _27664_, _27661_);
  nor (_27666_, _27665_, _19975_);
  nor (_27667_, _27666_, _27654_);
  nor (_27668_, _27667_, _25561_);
  nor (_27669_, _27668_, _27653_);
  nor (_01089_, _27669_, rst);
  and (_27670_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and (_27671_, _19975_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_27672_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_27673_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_27674_, _27673_, _27672_);
  and (_27675_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_27676_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_27677_, _27676_, _27675_);
  and (_27678_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_27679_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_27680_, _27679_, _27678_);
  and (_27681_, _27680_, _27677_);
  and (_27682_, _27681_, _27674_);
  nor (_27683_, _27682_, _19975_);
  nor (_27684_, _27683_, _27671_);
  nor (_27685_, _27684_, _25561_);
  nor (_27686_, _27685_, _27670_);
  nor (_01091_, _27686_, rst);
  and (_27687_, _25561_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and (_27688_, _19975_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_27689_, _20084_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_27690_, _20194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_27691_, _27690_, _27689_);
  and (_27692_, _20150_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_27693_, _20007_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_27694_, _27693_, _27692_);
  and (_27695_, _20106_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_27696_, _20051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_27697_, _27696_, _27695_);
  and (_27698_, _27697_, _27694_);
  and (_27699_, _27698_, _27691_);
  nor (_27700_, _27699_, _19975_);
  nor (_27701_, _27700_, _27688_);
  nor (_27702_, _27701_, _25561_);
  nor (_27703_, _27702_, _27687_);
  nor (_01094_, _27703_, rst);
  nor (_27704_, _25849_, _25618_);
  and (_27705_, _25935_, _25762_);
  and (_27706_, _27705_, _27704_);
  and (_27707_, _27706_, _25676_);
  and (_27708_, _25935_, _25761_);
  and (_27709_, _27708_, _27704_);
  and (_27710_, _27709_, _25676_);
  nor (_27711_, _27710_, _27707_);
  nor (_27712_, _25850_, _25618_);
  and (_27713_, _27712_, _27705_);
  and (_27714_, _27713_, _25676_);
  and (_27715_, _27712_, _27708_);
  and (_27716_, _27715_, _25676_);
  nor (_27717_, _27716_, _27714_);
  and (_27718_, _27717_, _27711_);
  and (_27719_, _27706_, _25677_);
  and (_27720_, _25935_, _25677_);
  and (_27721_, _27720_, _27712_);
  nor (_27722_, _27721_, _27719_);
  and (_27723_, _25676_, _25850_);
  nor (_27724_, _25935_, _25618_);
  and (_27725_, _27724_, _25761_);
  and (_27726_, _27725_, _27723_);
  and (_27727_, _27724_, _25762_);
  and (_27728_, _27727_, _27723_);
  nor (_27729_, _27728_, _27726_);
  and (_27730_, _25676_, _25849_);
  and (_27731_, _27727_, _27730_);
  and (_27732_, _27709_, _25677_);
  nor (_27733_, _27732_, _27731_);
  and (_27734_, _27733_, _27729_);
  and (_27735_, _27734_, _27722_);
  and (_27736_, _27735_, _27718_);
  not (_27737_, _27736_);
  nor (_27738_, _22442_, _22289_);
  nor (_27739_, _27738_, _22245_);
  not (_27740_, _27739_);
  and (_27741_, _22793_, _23270_);
  nor (_27742_, _27741_, _23000_);
  and (_27743_, _27742_, _27740_);
  nor (_27744_, _23510_, _22848_);
  and (_27745_, _21872_, _21082_);
  and (_27746_, _27745_, _22343_);
  nor (_27747_, _27746_, _23433_);
  and (_27748_, _27747_, _27744_);
  and (_27749_, _27748_, _27743_);
  and (_27750_, _22618_, _22267_);
  nor (_27751_, _27750_, _22650_);
  and (_27752_, _23052_, _23270_);
  not (_27753_, _27752_);
  nor (_27754_, _23096_, _22881_);
  and (_27755_, _27754_, _27753_);
  and (_27756_, _27755_, _27751_);
  and (_27757_, _27756_, _27749_);
  and (_27758_, _27757_, _22563_);
  nor (_27759_, _27758_, _19843_);
  nor (_27760_, _27759_, _27718_);
  nor (_27761_, _25618_, _17307_);
  and (_27762_, _25618_, _17307_);
  nor (_27763_, _27762_, _27761_);
  nor (_27764_, _25849_, _17937_);
  and (_27765_, _25849_, _17937_);
  nor (_27766_, _27765_, _27764_);
  nor (_27767_, _27766_, _27763_);
  nor (_27768_, _25761_, _17448_);
  and (_27769_, _25761_, _17448_);
  nor (_27770_, _27769_, _27768_);
  nor (_27771_, _25935_, _17579_);
  and (_27772_, _25935_, _17579_);
  nor (_27773_, _27772_, _27771_);
  nor (_27774_, _27773_, _27770_);
  nor (_27775_, _25676_, _17742_);
  and (_27776_, _25676_, _17742_);
  nor (_27777_, _27776_, _27775_);
  not (_27778_, _27777_);
  and (_27779_, _27778_, _27774_);
  and (_27780_, _27779_, _27767_);
  and (_27781_, _27780_, _24445_);
  not (_27782_, _27781_);
  nor (_27783_, _27782_, _27760_);
  and (_27784_, _27783_, _27737_);
  and (_27785_, _27731_, _24522_);
  not (_27786_, _25888_);
  and (_27787_, _25714_, _27786_);
  and (_27788_, _19898_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_27789_, _27788_);
  and (_27790_, _27789_, p1in_reg[6]);
  and (_27791_, _27788_, p1_in[6]);
  nor (_27792_, _27791_, _27790_);
  nor (_27793_, _27792_, _27759_);
  and (_27794_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_27795_, _27794_, _27793_);
  not (_27796_, _27795_);
  nor (_27797_, _27796_, _25798_);
  and (_27798_, _27789_, p1in_reg[2]);
  and (_27799_, _27788_, p1_in[2]);
  nor (_27800_, _27799_, _27798_);
  not (_27801_, _27800_);
  nor (_27802_, _27801_, _27759_);
  and (_27803_, _27759_, _24813_);
  nor (_27804_, _27803_, _27802_);
  and (_27805_, _27804_, _25798_);
  or (_27806_, _27805_, _27797_);
  and (_27807_, _27806_, _27787_);
  and (_27808_, _27789_, p1in_reg[1]);
  and (_27809_, _27788_, p1_in[1]);
  nor (_27810_, _27809_, _27808_);
  nor (_27811_, _27810_, _27759_);
  and (_27812_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_27813_, _27812_, _27811_);
  not (_27814_, _27813_);
  nand (_27815_, _27814_, _25798_);
  nor (_27816_, _25714_, _27786_);
  and (_27817_, _27789_, p1in_reg[5]);
  and (_27818_, _27788_, p1_in[5]);
  nor (_27819_, _27818_, _27817_);
  not (_27820_, _27819_);
  nor (_27821_, _27820_, _27759_);
  and (_27822_, _27759_, _24855_);
  nor (_27823_, _27822_, _27821_);
  or (_27824_, _27823_, _25798_);
  and (_27825_, _27824_, _27816_);
  and (_27826_, _27825_, _27815_);
  nor (_27827_, _25714_, _25888_);
  and (_27828_, _27789_, p1in_reg[7]);
  and (_27829_, _27788_, p1_in[7]);
  nor (_27830_, _27829_, _27828_);
  nor (_27831_, _27830_, _27759_);
  and (_27832_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_27833_, _27832_, _27831_);
  not (_27834_, _27833_);
  nor (_27835_, _27834_, _25798_);
  and (_27836_, _27789_, p1in_reg[3]);
  and (_27837_, _27788_, p1_in[3]);
  nor (_27838_, _27837_, _27836_);
  not (_27839_, _27838_);
  nor (_27840_, _27839_, _27759_);
  and (_27841_, _27759_, _24827_);
  nor (_27842_, _27841_, _27840_);
  and (_27843_, _27842_, _25798_);
  or (_27844_, _27843_, _27835_);
  and (_27845_, _27844_, _27827_);
  and (_27846_, _27789_, p1in_reg[0]);
  and (_27847_, _27788_, p1_in[0]);
  nor (_27848_, _27847_, _27846_);
  nor (_27849_, _27848_, _27759_);
  and (_27850_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_27851_, _27850_, _27849_);
  not (_27852_, _27851_);
  nand (_27853_, _27852_, _25798_);
  and (_27854_, _25714_, _25888_);
  and (_27855_, _27789_, p1in_reg[4]);
  and (_27856_, _27788_, p1_in[4]);
  nor (_27857_, _27856_, _27855_);
  not (_27858_, _27857_);
  nor (_27859_, _27858_, _27759_);
  and (_27860_, _27759_, _24841_);
  nor (_27861_, _27860_, _27859_);
  or (_27862_, _27861_, _25798_);
  and (_27863_, _27862_, _27854_);
  and (_27864_, _27863_, _27853_);
  or (_27865_, _27864_, _27845_);
  or (_27866_, _27865_, _27826_);
  or (_27867_, _27866_, _27807_);
  and (_27868_, _27867_, _27710_);
  not (_27869_, _25798_);
  and (_27870_, _27869_, _24517_);
  and (_27871_, _25798_, _24471_);
  or (_27872_, _27871_, _27870_);
  and (_27873_, _27872_, _27787_);
  or (_27874_, _27869_, _24459_);
  or (_27875_, _25798_, _24504_);
  and (_27876_, _27875_, _27816_);
  and (_27877_, _27876_, _27874_);
  or (_27878_, _27869_, _24489_);
  or (_27879_, _25798_, _24451_);
  and (_27880_, _27879_, _27827_);
  and (_27881_, _27880_, _27878_);
  nor (_27882_, _24591_, _24580_);
  and (_27883_, _24591_, _24580_);
  nor (_27884_, _27883_, _27882_);
  and (_27885_, _24569_, _24556_);
  nor (_27886_, _24569_, _24556_);
  or (_27887_, _27886_, _27885_);
  nor (_27888_, _27887_, _27884_);
  and (_27889_, _27887_, _27884_);
  nor (_27890_, _27889_, _27888_);
  and (_27891_, _24603_, _24541_);
  nor (_27892_, _24603_, _24541_);
  or (_27893_, _27892_, _27891_);
  not (_27894_, _27893_);
  and (_27895_, _24625_, _24613_);
  nor (_27896_, _24625_, _24613_);
  or (_27897_, _27896_, _27895_);
  and (_27898_, _27897_, _27894_);
  nor (_27899_, _27897_, _27894_);
  nor (_27900_, _27899_, _27898_);
  nor (_27901_, _27900_, _27890_);
  and (_27902_, _27900_, _27890_);
  nor (_27903_, _27902_, _27901_);
  or (_27904_, _27903_, _27869_);
  or (_27905_, _25798_, _24496_);
  and (_27906_, _27905_, _27854_);
  and (_27907_, _27906_, _27904_);
  or (_27908_, _27907_, _27881_);
  or (_27909_, _27908_, _27877_);
  or (_27910_, _27909_, _27873_);
  and (_27911_, _27910_, _27726_);
  or (_27912_, _27911_, _27868_);
  nor (_27913_, _25798_, _19383_);
  and (_27914_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_27915_, _27914_, _27913_);
  and (_27916_, _27915_, _27854_);
  or (_27917_, _27869_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_27918_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_27919_, _27918_, _27827_);
  and (_27920_, _27919_, _27917_);
  and (_27921_, _27869_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_27922_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_27923_, _27922_, _27921_);
  and (_27924_, _27923_, _27816_);
  nand (_27925_, _25798_, _19021_);
  or (_27926_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_27927_, _27926_, _27787_);
  and (_27928_, _27927_, _27925_);
  or (_27929_, _27928_, _27924_);
  or (_27930_, _27929_, _27920_);
  or (_27931_, _27930_, _27916_);
  and (_27932_, _27931_, _27728_);
  nor (_27933_, _25798_, _24614_);
  and (_27934_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_27935_, _27934_, _27933_);
  and (_27936_, _27935_, _27787_);
  or (_27937_, _27869_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_27938_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_27939_, _27938_, _27816_);
  and (_27940_, _27939_, _27937_);
  nor (_27941_, _25798_, _24529_);
  and (_27942_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_27943_, _27942_, _27941_);
  and (_27944_, _27943_, _27827_);
  not (_27945_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nand (_27946_, _25798_, _27945_);
  or (_27947_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_27948_, _27947_, _27854_);
  and (_27949_, _27948_, _27946_);
  or (_27950_, _27949_, _27944_);
  or (_27951_, _27950_, _27940_);
  or (_27952_, _27951_, _27936_);
  and (_27953_, _27952_, _27731_);
  or (_27954_, _27953_, _27932_);
  or (_27955_, _27954_, _27912_);
  and (_27956_, _27869_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_27957_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_27958_, _27957_, _27956_);
  and (_27959_, _27958_, _27787_);
  nand (_27960_, _25798_, _25101_);
  or (_27961_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_27962_, _27961_, _27816_);
  and (_27963_, _27962_, _27960_);
  nand (_27964_, _25798_, _25106_);
  or (_27965_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_27966_, _27965_, _27827_);
  and (_27967_, _27966_, _27964_);
  nand (_27968_, _25798_, _25103_);
  or (_27969_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_27970_, _27969_, _27854_);
  and (_27971_, _27970_, _27968_);
  or (_27972_, _27971_, _27967_);
  or (_27973_, _27972_, _27963_);
  or (_27974_, _27973_, _27959_);
  and (_27975_, _27974_, _27719_);
  and (_27976_, _27789_, p2in_reg[6]);
  and (_27977_, _27788_, p2_in[6]);
  nor (_27978_, _27977_, _27976_);
  nor (_27979_, _27978_, _27759_);
  and (_27980_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_27981_, _27980_, _27979_);
  not (_27982_, _27981_);
  nor (_27983_, _27982_, _25798_);
  and (_27984_, _27789_, p2in_reg[2]);
  and (_27985_, _27788_, p2_in[2]);
  nor (_27986_, _27985_, _27984_);
  not (_27987_, _27986_);
  nor (_27988_, _27987_, _27759_);
  and (_27989_, _27759_, _24911_);
  nor (_27990_, _27989_, _27988_);
  and (_27991_, _27990_, _25798_);
  or (_27992_, _27991_, _27983_);
  and (_27994_, _27992_, _27787_);
  and (_27996_, _27789_, p2in_reg[1]);
  and (_27998_, _27788_, p2_in[1]);
  nor (_28000_, _27998_, _27996_);
  nor (_28002_, _28000_, _27759_);
  and (_28004_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_28006_, _28004_, _28002_);
  not (_28008_, _28006_);
  nand (_28010_, _28008_, _25798_);
  and (_28012_, _27789_, p2in_reg[5]);
  and (_28014_, _27788_, p2_in[5]);
  nor (_28016_, _28014_, _28012_);
  not (_28018_, _28016_);
  nor (_28020_, _28018_, _27759_);
  and (_28022_, _27759_, _24952_);
  nor (_28024_, _28022_, _28020_);
  or (_28026_, _28024_, _25798_);
  and (_28028_, _28026_, _27816_);
  and (_28030_, _28028_, _28010_);
  and (_28032_, _27789_, p2in_reg[7]);
  and (_28034_, _27788_, p2_in[7]);
  nor (_28036_, _28034_, _28032_);
  nor (_28038_, _28036_, _27759_);
  and (_28040_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_28042_, _28040_, _28038_);
  not (_28044_, _28042_);
  nor (_28046_, _28044_, _25798_);
  and (_28048_, _27789_, p2in_reg[3]);
  and (_28050_, _27788_, p2_in[3]);
  nor (_28052_, _28050_, _28048_);
  not (_28054_, _28052_);
  nor (_28055_, _28054_, _27759_);
  and (_28056_, _27759_, _24925_);
  nor (_28057_, _28056_, _28055_);
  and (_28058_, _28057_, _25798_);
  or (_28059_, _28058_, _28046_);
  and (_28060_, _28059_, _27827_);
  and (_28061_, _27789_, p2in_reg[0]);
  and (_28062_, _27788_, p2_in[0]);
  nor (_28063_, _28062_, _28061_);
  nor (_28064_, _28063_, _27759_);
  and (_28065_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_28066_, _28065_, _28064_);
  not (_28067_, _28066_);
  nand (_28068_, _28067_, _25798_);
  and (_28069_, _27789_, p2in_reg[4]);
  and (_28070_, _27788_, p2_in[4]);
  nor (_28071_, _28070_, _28069_);
  not (_28072_, _28071_);
  nor (_28073_, _28072_, _27759_);
  and (_28074_, _27759_, _24938_);
  nor (_28075_, _28074_, _28073_);
  or (_28076_, _28075_, _25798_);
  and (_28077_, _28076_, _27854_);
  and (_28078_, _28077_, _28068_);
  or (_28079_, _28078_, _28060_);
  or (_28080_, _28079_, _28030_);
  or (_28081_, _28080_, _27994_);
  and (_28082_, _28081_, _27714_);
  or (_28083_, _28082_, _27975_);
  and (_28084_, _27789_, p0in_reg[2]);
  and (_28085_, _27788_, p0_in[2]);
  nor (_28086_, _28085_, _28084_);
  nor (_28087_, _28086_, _27759_);
  and (_28088_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_28089_, _28088_, _28087_);
  not (_28090_, _28089_);
  nand (_28091_, _28090_, _25798_);
  and (_28092_, _27789_, p0in_reg[6]);
  and (_28093_, _27788_, p0_in[6]);
  nor (_28094_, _28093_, _28092_);
  not (_28095_, _28094_);
  nor (_28096_, _28095_, _27759_);
  and (_28097_, _27759_, _24778_);
  nor (_28098_, _28097_, _28096_);
  or (_28099_, _28098_, _25798_);
  and (_28100_, _28099_, _27787_);
  and (_28101_, _28100_, _28091_);
  and (_28102_, _27789_, p0in_reg[5]);
  and (_28103_, _27788_, p0_in[5]);
  nor (_28104_, _28103_, _28102_);
  nor (_28105_, _28104_, _27759_);
  and (_28106_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_28107_, _28106_, _28105_);
  not (_28108_, _28107_);
  nor (_28109_, _28108_, _25798_);
  and (_28110_, _27789_, p0in_reg[1]);
  and (_28111_, _27788_, p0_in[1]);
  nor (_28112_, _28111_, _28110_);
  not (_28113_, _28112_);
  nor (_28114_, _28113_, _27759_);
  and (_28115_, _27759_, _24715_);
  nor (_28116_, _28115_, _28114_);
  and (_28117_, _28116_, _25798_);
  or (_28118_, _28117_, _28109_);
  and (_28119_, _28118_, _27816_);
  and (_28120_, _27789_, p0in_reg[4]);
  and (_28121_, _27788_, p0_in[4]);
  nor (_28122_, _28121_, _28120_);
  nor (_28123_, _28122_, _27759_);
  and (_28124_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_28125_, _28124_, _28123_);
  not (_28126_, _28125_);
  nor (_28127_, _28126_, _25798_);
  and (_28128_, _27789_, p0in_reg[0]);
  and (_28129_, _27788_, p0_in[0]);
  nor (_28130_, _28129_, _28128_);
  not (_28131_, _28130_);
  nor (_28132_, _28131_, _27759_);
  and (_28133_, _27759_, _24699_);
  nor (_28134_, _28133_, _28132_);
  and (_28135_, _28134_, _25798_);
  or (_28136_, _28135_, _28127_);
  and (_28137_, _28136_, _27854_);
  and (_28139_, _27789_, p0in_reg[3]);
  and (_28140_, _27788_, p0_in[3]);
  nor (_28141_, _28140_, _28139_);
  nor (_28142_, _28141_, _27759_);
  and (_28143_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_28144_, _28143_, _28142_);
  not (_28145_, _28144_);
  nand (_28146_, _28145_, _25798_);
  and (_28147_, _27789_, p0in_reg[7]);
  and (_28148_, _27788_, p0_in[7]);
  nor (_28149_, _28148_, _28147_);
  not (_28151_, _28149_);
  nor (_28152_, _28151_, _27759_);
  and (_28153_, _27759_, _24631_);
  nor (_28154_, _28153_, _28152_);
  or (_28155_, _28154_, _25798_);
  and (_28156_, _28155_, _27827_);
  and (_28157_, _28156_, _28146_);
  or (_28158_, _28157_, _28137_);
  or (_28159_, _28158_, _28119_);
  or (_28160_, _28159_, _28101_);
  and (_28161_, _28160_, _27716_);
  and (_28162_, _27789_, p3in_reg[4]);
  and (_28163_, _27788_, p3_in[4]);
  nor (_28164_, _28163_, _28162_);
  nor (_28165_, _28164_, _27759_);
  and (_28166_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_28167_, _28166_, _28165_);
  not (_28168_, _28167_);
  nor (_28169_, _28168_, _25798_);
  and (_28170_, _27789_, p3in_reg[0]);
  and (_28171_, _27788_, p3_in[0]);
  nor (_28172_, _28171_, _28170_);
  not (_28173_, _28172_);
  nor (_28174_, _28173_, _27759_);
  and (_28175_, _27759_, _24981_);
  nor (_28176_, _28175_, _28174_);
  and (_28177_, _28176_, _25798_);
  or (_28178_, _28177_, _28169_);
  and (_28179_, _28178_, _27854_);
  and (_28180_, _27789_, p3in_reg[7]);
  and (_28182_, _27788_, p3_in[7]);
  nor (_28183_, _28182_, _28180_);
  nor (_28184_, _28183_, _27759_);
  and (_28185_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_28186_, _28185_, _28184_);
  not (_28187_, _28186_);
  nor (_28188_, _28187_, _25798_);
  and (_28189_, _27789_, p3in_reg[3]);
  and (_28190_, _27788_, p3_in[3]);
  nor (_28191_, _28190_, _28189_);
  not (_28192_, _28191_);
  nor (_28193_, _28192_, _27759_);
  and (_28194_, _27759_, _25022_);
  nor (_28195_, _28194_, _28193_);
  and (_28196_, _28195_, _25798_);
  or (_28197_, _28196_, _28188_);
  and (_28198_, _28197_, _27827_);
  or (_28199_, _28198_, _28179_);
  and (_28200_, _27789_, p3in_reg[6]);
  and (_28201_, _27788_, p3_in[6]);
  nor (_28203_, _28201_, _28200_);
  nor (_28204_, _28203_, _27759_);
  and (_28205_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_28206_, _28205_, _28204_);
  not (_28207_, _28206_);
  nor (_28208_, _28207_, _25798_);
  and (_28209_, _27789_, p3in_reg[2]);
  and (_28210_, _27788_, p3_in[2]);
  nor (_28211_, _28210_, _28209_);
  not (_28212_, _28211_);
  nor (_28213_, _28212_, _27759_);
  and (_28214_, _27759_, _25008_);
  nor (_28215_, _28214_, _28213_);
  and (_28216_, _28215_, _25798_);
  or (_28217_, _28216_, _28208_);
  and (_28218_, _28217_, _27787_);
  and (_28219_, _27789_, p3in_reg[5]);
  and (_28220_, _27788_, p3_in[5]);
  nor (_28221_, _28220_, _28219_);
  nor (_28222_, _28221_, _27759_);
  and (_28223_, _27759_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_28224_, _28223_, _28222_);
  not (_28225_, _28224_);
  nor (_28226_, _28225_, _25798_);
  and (_28227_, _27789_, p3in_reg[1]);
  and (_28228_, _27788_, p3_in[1]);
  nor (_28229_, _28228_, _28227_);
  not (_28230_, _28229_);
  nor (_28231_, _28230_, _27759_);
  and (_28232_, _27759_, _24994_);
  nor (_28233_, _28232_, _28231_);
  and (_28234_, _28233_, _25798_);
  or (_28235_, _28234_, _28226_);
  and (_28236_, _28235_, _27816_);
  or (_28237_, _28236_, _28218_);
  or (_28238_, _28237_, _28199_);
  and (_28239_, _28238_, _27707_);
  or (_28240_, _28239_, _28161_);
  or (_28241_, _28240_, _28083_);
  nor (_28242_, _25798_, _18081_);
  and (_28243_, _25798_, _18081_);
  nor (_28244_, _28243_, _28242_);
  nor (_28245_, _28244_, _27777_);
  nor (_28246_, _25888_, _18333_);
  and (_28247_, _25888_, _18333_);
  nor (_28248_, _28247_, _28246_);
  nor (_28249_, _25714_, _18212_);
  and (_28250_, _25714_, _18212_);
  nor (_28251_, _28250_, _28249_);
  nor (_28252_, _28251_, _28248_);
  and (_28253_, _28252_, _28245_);
  and (_28254_, _27774_, _27767_);
  and (_28255_, _28254_, _28253_);
  nand (_28256_, _28255_, _16959_);
  nor (_28257_, _28256_, _27736_);
  and (_28258_, _27827_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_28259_, _27787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_28260_, _28259_, _25798_);
  or (_28261_, _28260_, _28258_);
  and (_28262_, _27827_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_28263_, _27787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_28264_, _28263_, _27869_);
  or (_28265_, _28264_, _28262_);
  and (_28266_, _28265_, _28261_);
  or (_28267_, _27869_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_28268_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_28269_, _28268_, _27854_);
  and (_28270_, _28269_, _28267_);
  and (_28271_, _27869_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_28272_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_28273_, _28272_, _28271_);
  and (_28274_, _28273_, _27816_);
  or (_28275_, _28274_, _25761_);
  or (_28276_, _28275_, _28270_);
  or (_28277_, _28276_, _28266_);
  and (_28278_, _27869_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_28279_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_28280_, _28279_, _28278_);
  and (_28281_, _28280_, _27816_);
  or (_28282_, _28281_, _25762_);
  nand (_28283_, _25798_, _25216_);
  or (_28284_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_28285_, _28284_, _27854_);
  and (_28286_, _28285_, _28283_);
  or (_28287_, _27869_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_28288_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_28289_, _28288_, _27827_);
  and (_28290_, _28289_, _28287_);
  and (_28291_, _27869_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_28292_, _25798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_28293_, _28292_, _28291_);
  and (_28294_, _28293_, _27787_);
  or (_28295_, _28294_, _28290_);
  or (_28296_, _28295_, _28286_);
  or (_28297_, _28296_, _28282_);
  and (_28298_, _28297_, _27721_);
  and (_28299_, _28298_, _28277_);
  or (_28300_, _28299_, _28257_);
  or (_28301_, _28300_, _28241_);
  or (_28302_, _28301_, _27955_);
  nand (_28303_, _28257_, _18388_);
  and (_28304_, _28303_, _28302_);
  or (_28305_, _28304_, _27785_);
  nand (_28306_, _27869_, _24603_);
  nand (_28307_, _25798_, _24556_);
  and (_28308_, _28307_, _27854_);
  and (_28309_, _28308_, _28306_);
  nor (_28310_, _27869_, _24580_);
  nor (_28311_, _25798_, _24625_);
  or (_28312_, _28311_, _28310_);
  and (_28313_, _28312_, _27787_);
  or (_28314_, _28313_, _28309_);
  nand (_28315_, _27869_, _24541_);
  nand (_28316_, _25798_, _24591_);
  and (_28317_, _28316_, _27827_);
  and (_28318_, _28317_, _28315_);
  nor (_28319_, _27869_, _24569_);
  nor (_28320_, _25798_, _24613_);
  or (_28321_, _28320_, _28319_);
  and (_28322_, _28321_, _27816_);
  or (_28323_, _28322_, _28318_);
  nor (_28324_, _28323_, _28314_);
  nand (_28325_, _28324_, _27785_);
  and (_28326_, _28325_, _28305_);
  or (_28327_, _28326_, _27784_);
  nor (_28328_, _25798_, _24502_);
  and (_28329_, _25798_, ABINPUT[4]);
  or (_28330_, _28329_, _28328_);
  and (_28331_, _28330_, _27816_);
  nand (_28332_, _25798_, _25445_);
  or (_28333_, _25798_, ABINPUT[9]);
  and (_28334_, _28333_, _27787_);
  and (_28335_, _28334_, _28332_);
  nor (_28336_, _25798_, _25247_);
  and (_28337_, _25798_, ABINPUT[6]);
  or (_28338_, _28337_, _28336_);
  and (_28339_, _28338_, _27827_);
  nand (_28340_, _25798_, _25437_);
  or (_28341_, _25798_, ABINPUT[7]);
  and (_28342_, _28341_, _27854_);
  and (_28343_, _28342_, _28340_);
  or (_28344_, _28343_, _28339_);
  or (_28345_, _28344_, _28335_);
  nor (_28346_, _28345_, _28331_);
  nand (_28347_, _28346_, _27784_);
  and (_28348_, _28347_, _27053_);
  and (_01506_, _28348_, _28327_);
  and (_28349_, _27854_, _25798_);
  and (_28350_, _28349_, _27731_);
  and (_28351_, _28350_, _24519_);
  not (_28352_, _24439_);
  and (_28353_, _28349_, _27726_);
  and (_28354_, _28353_, _28352_);
  nor (_28355_, _28354_, _28351_);
  not (_28356_, _24334_);
  and (_28357_, _25676_, _25798_);
  and (_28358_, _28357_, _27827_);
  nand (_28359_, _28358_, _27715_);
  or (_28360_, _28359_, _28356_);
  and (_28361_, _28360_, _28355_);
  nor (_28362_, _28361_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_28363_, _24432_);
  and (_28364_, _27827_, _27869_);
  nor (_28365_, _28364_, _28363_);
  and (_28366_, _28365_, _27780_);
  nor (_28367_, _24047_, _17307_);
  and (_28368_, _28367_, _28255_);
  and (_28369_, _28349_, _27785_);
  or (_28370_, _28369_, _28368_);
  or (_28371_, _28370_, _28366_);
  or (_28372_, _28371_, _28362_);
  and (_28373_, _28357_, _27715_);
  and (_28374_, _28373_, _27787_);
  nand (_28375_, _28374_, _24334_);
  and (_28376_, _28375_, _27053_);
  and (_01508_, _28376_, _28372_);
  and (_28377_, _28372_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_28378_, _28349_, _25677_);
  and (_28379_, _28378_, _27706_);
  nand (_28380_, _28379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand (_28381_, _28374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_28382_, _28381_, _28380_);
  and (_28383_, _28378_, _27715_);
  nand (_28384_, _28383_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_28385_, _28378_, _27713_);
  nand (_28386_, _28385_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_28387_, _28386_, _28384_);
  and (_28388_, _28387_, _28382_);
  and (_28389_, _28349_, _27728_);
  nand (_28390_, _28389_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  not (_28391_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_28392_, _28359_, _28391_);
  and (_28393_, _28392_, _28390_);
  not (_28394_, _27706_);
  nand (_28395_, _28357_, _27854_);
  or (_28396_, _28395_, _28394_);
  or (_28397_, _28396_, _28187_);
  not (_28398_, _27715_);
  nand (_28399_, _28357_, _27816_);
  or (_28400_, _28399_, _28398_);
  or (_28401_, _28400_, _24288_);
  and (_28402_, _28401_, _28397_);
  and (_28403_, _28402_, _28393_);
  and (_28404_, _28403_, _28388_);
  nand (_28405_, _28350_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand (_28406_, _28349_, _27714_);
  or (_28407_, _28406_, _28044_);
  not (_28408_, _27709_);
  or (_28409_, _28395_, _28408_);
  or (_28410_, _28409_, _27834_);
  and (_28411_, _28410_, _28407_);
  not (_28412_, _28154_);
  or (_28413_, _28395_, _28398_);
  or (_28414_, _28413_, _28412_);
  nand (_28415_, _28353_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_28416_, _28415_, _28414_);
  and (_28417_, _28416_, _28411_);
  and (_28418_, _28417_, _28405_);
  and (_28419_, _28418_, _28404_);
  or (_28420_, _28419_, _28372_);
  nand (_28421_, _28420_, _28375_);
  or (_28422_, _28421_, _28377_);
  or (_28423_, _28375_, ABINPUT[26]);
  and (_28424_, _28423_, _27053_);
  and (_01510_, _28424_, _28422_);
  nor (_01513_, _25636_, rst);
  and (_28425_, _28372_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_28426_, _28379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nand (_28427_, _28374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_28428_, _28427_, _28426_);
  nand (_28429_, _28383_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_28430_, _28385_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_28431_, _28430_, _28429_);
  and (_28432_, _28431_, _28428_);
  nand (_28433_, _28389_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not (_28434_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_28435_, _28359_, _28434_);
  and (_28436_, _28435_, _28433_);
  not (_28437_, _28176_);
  or (_28439_, _28396_, _28437_);
  or (_28440_, _28400_, _24296_);
  and (_28441_, _28440_, _28439_);
  and (_28442_, _28441_, _28436_);
  and (_28443_, _28442_, _28432_);
  nand (_28445_, _28350_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_28446_, _28406_, _28067_);
  or (_28447_, _28409_, _27852_);
  and (_28448_, _28447_, _28446_);
  not (_28449_, _28134_);
  or (_28451_, _28413_, _28449_);
  nand (_28452_, _28353_, _27903_);
  and (_28453_, _28452_, _28451_);
  and (_28454_, _28453_, _28448_);
  and (_28455_, _28454_, _28445_);
  and (_28457_, _28455_, _28443_);
  or (_28458_, _28457_, _28372_);
  nand (_28459_, _28458_, _28375_);
  or (_28460_, _28459_, _28425_);
  or (_28461_, _28375_, ABINPUT[19]);
  and (_28463_, _28461_, _27053_);
  and (_02181_, _28463_, _28460_);
  and (_28464_, _28372_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_28465_, _28379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nand (_28466_, _28374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_28468_, _28466_, _28465_);
  nand (_28469_, _28383_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand (_28470_, _28385_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_28471_, _28470_, _28469_);
  and (_28472_, _28471_, _28468_);
  nand (_28474_, _28389_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  not (_28475_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_28477_, _28359_, _28475_);
  and (_28478_, _28477_, _28474_);
  not (_28479_, _28233_);
  or (_28480_, _28396_, _28479_);
  or (_28481_, _28400_, _24302_);
  and (_28482_, _28481_, _28480_);
  and (_28483_, _28482_, _28478_);
  and (_28485_, _28483_, _28472_);
  nand (_28486_, _28350_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_28487_, _28406_, _28008_);
  or (_28489_, _28409_, _27814_);
  and (_28490_, _28489_, _28487_);
  not (_28491_, _28116_);
  or (_28493_, _28413_, _28491_);
  nand (_28494_, _28353_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_28495_, _28494_, _28493_);
  and (_28497_, _28495_, _28490_);
  and (_28498_, _28497_, _28486_);
  and (_28499_, _28498_, _28485_);
  or (_28501_, _28499_, _28372_);
  nand (_28502_, _28501_, _28375_);
  or (_28503_, _28502_, _28464_);
  or (_28505_, _28375_, ABINPUT[20]);
  and (_28506_, _28505_, _27053_);
  and (_02183_, _28506_, _28503_);
  and (_28508_, _28372_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_28509_, _28379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nand (_28511_, _28374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_28512_, _28511_, _28509_);
  nand (_28513_, _28383_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand (_28514_, _28385_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_28515_, _28514_, _28513_);
  and (_28516_, _28515_, _28512_);
  nand (_28517_, _28389_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_28519_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_28520_, _28359_, _28519_);
  and (_28521_, _28520_, _28517_);
  not (_28523_, _28215_);
  or (_28524_, _28396_, _28523_);
  or (_28525_, _28400_, _24308_);
  and (_28527_, _28525_, _28524_);
  and (_28528_, _28527_, _28521_);
  and (_28529_, _28528_, _28516_);
  nand (_28531_, _28350_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not (_28532_, _27990_);
  or (_28533_, _28406_, _28532_);
  not (_28535_, _27804_);
  or (_28536_, _28409_, _28535_);
  and (_28537_, _28536_, _28533_);
  nand (_28539_, _28353_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_28540_, _28413_, _28090_);
  and (_28541_, _28540_, _28539_);
  and (_28543_, _28541_, _28537_);
  and (_28544_, _28543_, _28531_);
  and (_28546_, _28544_, _28529_);
  or (_28547_, _28546_, _28372_);
  nand (_28548_, _28547_, _28375_);
  or (_28549_, _28548_, _28508_);
  or (_28550_, _28375_, ABINPUT[21]);
  and (_28552_, _28550_, _27053_);
  and (_02185_, _28552_, _28549_);
  and (_28553_, _28372_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_28555_, _28379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nand (_28556_, _28374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_28557_, _28556_, _28555_);
  nand (_28559_, _28383_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand (_28560_, _28385_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_28561_, _28560_, _28559_);
  and (_28563_, _28561_, _28557_);
  nand (_28564_, _28389_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not (_28565_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_28567_, _28359_, _28565_);
  and (_28568_, _28567_, _28564_);
  not (_28569_, _28195_);
  or (_28571_, _28396_, _28569_);
  or (_28572_, _28400_, _24314_);
  and (_28573_, _28572_, _28571_);
  and (_28575_, _28573_, _28568_);
  and (_28576_, _28575_, _28563_);
  nand (_28578_, _28350_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  not (_28579_, _28057_);
  or (_28580_, _28406_, _28579_);
  not (_28581_, _27842_);
  or (_28582_, _28409_, _28581_);
  and (_28583_, _28582_, _28580_);
  or (_28584_, _28413_, _28145_);
  nand (_28586_, _28353_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_28587_, _28586_, _28584_);
  and (_28588_, _28587_, _28583_);
  and (_28590_, _28588_, _28578_);
  and (_28591_, _28590_, _28576_);
  or (_28592_, _28591_, _28372_);
  nand (_28594_, _28592_, _28375_);
  or (_28595_, _28594_, _28553_);
  or (_28596_, _28375_, ABINPUT[22]);
  and (_28598_, _28596_, _27053_);
  and (_02187_, _28598_, _28595_);
  and (_28599_, _28372_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_28601_, _28379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nand (_28602_, _28374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_28603_, _28602_, _28601_);
  nand (_28605_, _28383_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand (_28606_, _28385_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_28607_, _28606_, _28605_);
  and (_28609_, _28607_, _28603_);
  nand (_28610_, _28389_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_28612_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_28613_, _28359_, _28612_);
  and (_28614_, _28613_, _28610_);
  or (_28615_, _28396_, _28168_);
  or (_28617_, _28400_, _24320_);
  and (_28618_, _28617_, _28615_);
  and (_28619_, _28618_, _28614_);
  and (_28621_, _28619_, _28609_);
  nand (_28622_, _28350_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not (_28623_, _28075_);
  or (_28625_, _28406_, _28623_);
  not (_28626_, _27861_);
  or (_28627_, _28409_, _28626_);
  and (_28629_, _28627_, _28625_);
  or (_28630_, _28413_, _28126_);
  nand (_28631_, _28353_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_28633_, _28631_, _28630_);
  and (_28634_, _28633_, _28629_);
  and (_28635_, _28634_, _28622_);
  and (_28637_, _28635_, _28621_);
  or (_28638_, _28637_, _28372_);
  nand (_28639_, _28638_, _28375_);
  or (_28641_, _28639_, _28599_);
  or (_28642_, _28375_, ABINPUT[23]);
  and (_28644_, _28642_, _27053_);
  and (_02189_, _28644_, _28641_);
  and (_28645_, _28372_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_28646_, _28374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand (_28648_, _28379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_28649_, _28648_, _28646_);
  nand (_28650_, _28383_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  nand (_28652_, _28385_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_28653_, _28652_, _28650_);
  and (_28654_, _28653_, _28649_);
  nand (_28656_, _28389_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_28657_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_28658_, _28359_, _28657_);
  and (_28660_, _28658_, _28656_);
  or (_28661_, _28396_, _28225_);
  or (_28662_, _28400_, _24326_);
  and (_28664_, _28662_, _28661_);
  and (_28665_, _28664_, _28660_);
  and (_28666_, _28665_, _28654_);
  nand (_28668_, _28350_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not (_28669_, _28024_);
  or (_28670_, _28406_, _28669_);
  not (_28672_, _27823_);
  or (_28673_, _28409_, _28672_);
  and (_28675_, _28673_, _28670_);
  or (_28676_, _28413_, _28108_);
  nand (_28677_, _28353_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_28678_, _28677_, _28676_);
  and (_28680_, _28678_, _28675_);
  and (_28681_, _28680_, _28668_);
  and (_28682_, _28681_, _28666_);
  or (_28684_, _28682_, _28372_);
  nand (_28685_, _28684_, _28375_);
  or (_28686_, _28685_, _28645_);
  or (_28688_, _28375_, ABINPUT[24]);
  and (_28689_, _28688_, _27053_);
  and (_02191_, _28689_, _28686_);
  and (_28691_, _28372_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_28692_, _28374_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  nand (_28693_, _28379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_28695_, _28693_, _28692_);
  nand (_28696_, _28383_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nand (_28697_, _28385_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_28699_, _28697_, _28696_);
  and (_28700_, _28699_, _28695_);
  nand (_28701_, _28389_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  not (_28703_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_28704_, _28359_, _28703_);
  and (_28706_, _28704_, _28701_);
  or (_28707_, _28396_, _28207_);
  or (_28708_, _28400_, _24332_);
  and (_28709_, _28708_, _28707_);
  and (_28710_, _28709_, _28706_);
  and (_28711_, _28710_, _28700_);
  nand (_28712_, _28350_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_28714_, _28406_, _27982_);
  or (_28715_, _28409_, _27796_);
  and (_28716_, _28715_, _28714_);
  nand (_28718_, _28353_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  not (_28719_, _28098_);
  or (_28720_, _28413_, _28719_);
  and (_28722_, _28720_, _28718_);
  and (_28723_, _28722_, _28716_);
  and (_28724_, _28723_, _28712_);
  and (_28726_, _28724_, _28711_);
  or (_28727_, _28726_, _28372_);
  nand (_28728_, _28727_, _28375_);
  or (_28730_, _28728_, _28691_);
  or (_28731_, _28375_, ABINPUT[25]);
  and (_28732_, _28731_, _27053_);
  and (_02193_, _28732_, _28730_);
  or (_28734_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_28735_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_28737_, _27788_, _28735_);
  and (_28738_, _28737_, _27053_);
  and (_02749_, _28738_, _28734_);
  and (_28740_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_28741_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  or (_28742_, _28741_, _28740_);
  and (_02753_, _28742_, _27053_);
  nor (_03131_, _25618_, rst);
  nor (_03138_, _25811_, rst);
  nor (_03142_, _25610_, rst);
  and (_28745_, _23291_, _22168_);
  nor (_28747_, _25634_, _22977_);
  not (_28748_, _28747_);
  nor (_28749_, _22977_, _19843_);
  nor (_28751_, _28745_, _28749_);
  and (_28752_, _28751_, _28748_);
  nor (_28753_, _28752_, _28745_);
  nor (_28755_, _24047_, _18355_);
  and (_28756_, _28755_, _28753_);
  and (_28757_, _28756_, _27780_);
  not (_28759_, _28757_);
  nor (_28760_, ABINPUT[28], ABINPUT[27]);
  nor (_28761_, ABINPUT[30], ABINPUT[29]);
  and (_28765_, _28761_, _28760_);
  nor (_28766_, ABINPUT[32], ABINPUT[31]);
  nor (_28774_, ABINPUT[33], ABINPUT[34]);
  and (_28775_, _28774_, _28766_);
  and (_28782_, _28775_, _28765_);
  not (_28790_, _23291_);
  and (_28792_, _28752_, _28790_);
  and (_28793_, _28792_, _28782_);
  and (_28806_, _28745_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_28811_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_28812_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_28819_, _28812_, _28811_);
  nor (_28828_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_28829_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_28837_, _28829_, _28828_);
  and (_28839_, _28837_, _28819_);
  and (_28840_, _28839_, _23807_);
  or (_28848_, _28840_, _28806_);
  nor (_28857_, _28848_, _28793_);
  not (_28858_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_28865_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _28858_);
  and (_28870_, _26110_, _26109_);
  and (_28871_, _26079_, _26077_);
  nor (_28884_, _28871_, _28870_);
  and (_28890_, _26051_, _26047_);
  and (_28891_, _26096_, _26095_);
  nor (_28903_, _28891_, _28890_);
  and (_28904_, _28903_, _28884_);
  and (_28911_, _26125_, _26124_);
  and (_28920_, _26063_, _26060_);
  nor (_28929_, _28920_, _28911_);
  and (_28930_, _26025_, _26024_);
  and (_28938_, _26140_, _26139_);
  nor (_28947_, _28938_, _28930_);
  and (_28948_, _28947_, _28929_);
  and (_28956_, _28948_, _28904_);
  nor (_28962_, _28956_, _28865_);
  and (_28963_, _28865_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_28977_, _28963_, _28962_);
  not (_28984_, _28977_);
  and (_28985_, _28984_, _28753_);
  not (_28997_, _28985_);
  and (_29002_, _28997_, _28857_);
  and (_29003_, _23280_, _22157_);
  nor (_29011_, _29003_, _23248_);
  or (_29013_, _29011_, _29002_);
  and (_29014_, _27745_, _22190_);
  not (_29015_, _29014_);
  and (_29017_, _22267_, _22135_);
  nor (_29018_, _29017_, _22453_);
  and (_29020_, _29018_, _29015_);
  and (_29021_, _23422_, _22387_);
  and (_29022_, _27745_, _22387_);
  nor (_29023_, _29022_, _29021_);
  and (_29024_, _29023_, _29020_);
  or (_29026_, _22954_, _22486_);
  or (_29027_, _29026_, _22618_);
  and (_29028_, _29027_, _22409_);
  not (_29030_, _29028_);
  and (_29031_, _29030_, _29024_);
  not (_29032_, _29031_);
  and (_29034_, _29032_, _29002_);
  and (_29035_, _22596_, _22409_);
  nor (_29036_, _29035_, _23631_);
  not (_29038_, _29036_);
  nor (_29039_, _29038_, _29034_);
  and (_29040_, _29039_, _29013_);
  nor (_29042_, _29040_, _25634_);
  nand (_29043_, _20600_, _20315_);
  nor (_29044_, _29043_, _21093_);
  and (_29046_, _22289_, _21115_);
  nor (_29047_, _29046_, _29044_);
  nor (_29048_, _29047_, _19843_);
  nor (_29050_, _29048_, _23302_);
  not (_29051_, _29050_);
  nor (_29053_, _29051_, _29042_);
  or (_29054_, _24474_, _28352_);
  nor (_29055_, _29054_, _24433_);
  not (_29056_, _29055_);
  and (_29058_, _29056_, _28745_);
  not (_29059_, _23807_);
  nor (_29060_, _24558_, _24547_);
  nor (_29062_, _29060_, _29059_);
  nor (_29063_, _29062_, _29058_);
  not (_29064_, _29063_);
  nor (_29066_, _29064_, _29053_);
  not (_29067_, _29066_);
  nor (_29068_, _29067_, _28368_);
  and (_29070_, _29068_, _28759_);
  nor (_29071_, _23313_, rst);
  and (_03151_, _29071_, _29070_);
  and (_03155_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _27053_);
  and (_03158_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _27053_);
  not (_29073_, _27584_);
  and (_29075_, _29023_, _29018_);
  nor (_29076_, _29075_, _25634_);
  not (_29077_, _29076_);
  not (_29079_, _19843_);
  and (_29080_, _22409_, _29079_);
  and (_29082_, _29080_, _22672_);
  and (_29083_, _23216_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_29084_, _29083_, _22782_);
  and (_29085_, _29046_, _29079_);
  or (_29087_, _29085_, _29084_);
  nor (_29088_, _29087_, _29082_);
  and (_29089_, _29088_, _29077_);
  and (_29091_, _29089_, _28748_);
  nor (_29092_, _29091_, _29073_);
  and (_29093_, _29091_, _25577_);
  nor (_29095_, _29093_, _29092_);
  not (_29096_, _29095_);
  and (_29097_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_29099_, _29097_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_29100_, _29095_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_29101_, _29095_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_29103_, _27703_);
  nor (_29104_, _29091_, _29103_);
  and (_29105_, _29091_, _25914_);
  nor (_29107_, _29105_, _29104_);
  and (_29108_, _29107_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_29109_, _29107_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_29111_, _29109_, _29108_);
  not (_29112_, _27686_);
  nor (_29114_, _29091_, _29112_);
  and (_29115_, _29091_, _25756_);
  nor (_29116_, _29115_, _29114_);
  and (_29117_, _29116_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_29119_, _29116_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_29120_, _27669_);
  nor (_29121_, _29091_, _29120_);
  and (_29123_, _29091_, _25828_);
  nor (_29124_, _29123_, _29121_);
  nand (_29125_, _29124_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_29127_, _27652_);
  nor (_29128_, _29091_, _29127_);
  and (_29129_, _29091_, _25671_);
  nor (_29131_, _29129_, _29128_);
  and (_29132_, _29131_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_29133_, _29131_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_29135_, _27635_);
  nor (_29136_, _29091_, _29135_);
  and (_29137_, _29091_, _25793_);
  nor (_29139_, _29137_, _29136_);
  and (_29140_, _29139_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_29141_, _27618_);
  nor (_29143_, _29091_, _29141_);
  and (_29144_, _29091_, _25866_);
  nor (_29145_, _29144_, _29143_);
  and (_29146_, _29145_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_29147_, _27601_);
  nor (_29148_, _29091_, _29147_);
  and (_29149_, _29091_, _25709_);
  nor (_29150_, _29149_, _29148_);
  and (_29151_, _29150_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_29152_, _29145_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_29153_, _29152_, _29146_);
  and (_29154_, _29153_, _29151_);
  nor (_29155_, _29154_, _29146_);
  not (_29156_, _29155_);
  nor (_29157_, _29139_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_29158_, _29157_, _29140_);
  and (_29159_, _29158_, _29156_);
  nor (_29160_, _29159_, _29140_);
  nor (_29161_, _29160_, _29133_);
  or (_29162_, _29161_, _29132_);
  or (_29163_, _29124_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_29164_, _29163_, _29125_);
  nand (_29165_, _29164_, _29162_);
  and (_29166_, _29165_, _29125_);
  nor (_29167_, _29166_, _29119_);
  or (_29168_, _29167_, _29117_);
  and (_29169_, _29168_, _29111_);
  nor (_29170_, _29169_, _29108_);
  nor (_29171_, _29170_, _29101_);
  or (_29172_, _29171_, _29100_);
  and (_29173_, _29172_, _29099_);
  and (_29174_, _29173_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_29175_, _29174_, _29096_);
  and (_29176_, _29175_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_29177_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_29178_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_29179_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_29180_, _29172_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_29181_, _29180_, _29179_);
  and (_29182_, _29181_, _29178_);
  not (_29183_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_29184_, _29095_, _29183_);
  and (_29185_, _29184_, _29182_);
  and (_29186_, _29185_, _29177_);
  nor (_29187_, _29186_, _29176_);
  nor (_29188_, _29095_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_29189_, _29095_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_29190_, _29189_, _29188_);
  not (_29191_, _29190_);
  nor (_29192_, _29191_, _29187_);
  nor (_29193_, _29095_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_29194_, _29095_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_29195_, _29194_, _29193_);
  nand (_29196_, _29195_, _29192_);
  nand (_29197_, _29196_, _28735_);
  or (_29198_, _29196_, _28735_);
  and (_29199_, _29036_, _29024_);
  nor (_29200_, _29199_, _25634_);
  not (_29201_, _29200_);
  and (_29202_, _22936_, _29079_);
  nor (_29203_, _29202_, _23291_);
  and (_29204_, _29203_, _28748_);
  and (_29205_, _29204_, _29201_);
  not (_29206_, _29205_);
  and (_29207_, _23631_, _23227_);
  nor (_29208_, _29207_, _29048_);
  not (_29209_, _29208_);
  nand (_29210_, _29209_, _29091_);
  and (_29211_, _29210_, _29206_);
  and (_29212_, _29211_, _29198_);
  and (_29213_, _29212_, _29197_);
  and (_29214_, _29205_, _29089_);
  and (_29215_, _29214_, _29208_);
  and (_29216_, _29215_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_29217_, _29207_, ABINPUT[18]);
  and (_29218_, _23313_, ABINPUT[26]);
  or (_29219_, _29218_, _29217_);
  or (_29220_, _29219_, _29216_);
  and (_29221_, _29085_, _25578_);
  and (_29222_, _29214_, _29209_);
  and (_29223_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_29224_, _29223_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_29225_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_29226_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_29227_, _29226_, _29225_);
  and (_29228_, _29227_, _29224_);
  and (_29229_, _29228_, _29099_);
  and (_29230_, _29229_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_29231_, _29230_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_29232_, _29231_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_29233_, _29232_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_29234_, _29233_, _28735_);
  and (_29235_, _29233_, _28735_);
  or (_29236_, _29235_, _29234_);
  and (_29237_, _29236_, _29222_);
  or (_29238_, _29237_, _29221_);
  nor (_29239_, _29238_, _29220_);
  nand (_29240_, _29239_, _29070_);
  or (_29241_, _29240_, _29213_);
  and (_29242_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_29243_, _20139_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_29244_, _29243_, _25561_);
  nor (_29245_, _29244_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_29246_, _29245_);
  and (_29247_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_29248_, _29247_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_29249_, _29248_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_29250_, _29249_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_29251_, _29250_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_29252_, _29251_, _29246_);
  and (_29253_, _29252_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_29254_, _29253_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_29255_, _29254_, _29242_);
  and (_29256_, _29255_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_29257_, _29256_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_29258_, _29257_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_29259_, _29258_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_29260_, _29258_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_29261_, _29260_, _29259_);
  or (_29262_, _29261_, _29070_);
  and (_29263_, _29262_, _27053_);
  and (_03161_, _29263_, _29241_);
  and (_29264_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _27053_);
  and (_29265_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_29266_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_29267_, _19887_, _29266_);
  not (_29268_, _29267_);
  not (_29269_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_29270_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_29271_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_29272_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_29273_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_29274_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_29275_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_29276_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_29277_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_29278_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_29279_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_29280_, _29279_, _29278_);
  and (_29281_, _29280_, _29277_);
  and (_29282_, _29281_, _29276_);
  and (_29283_, _29282_, _29275_);
  and (_29284_, _29283_, _29274_);
  and (_29285_, _29284_, _29273_);
  and (_29286_, _29285_, _29272_);
  and (_29287_, _29286_, _29271_);
  and (_29288_, _29287_, _29270_);
  nor (_29289_, _29288_, _29269_);
  and (_29290_, _29288_, _29269_);
  nor (_29291_, _29290_, _29289_);
  nor (_29292_, _29287_, _29270_);
  or (_29293_, _29292_, _29288_);
  and (_29294_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_29295_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_29296_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_29297_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_29298_, _29297_, _29295_);
  and (_29299_, _29298_, _29296_);
  nor (_29300_, _29299_, _29295_);
  nor (_29301_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_29302_, _29301_, _29294_);
  not (_29303_, _29302_);
  nor (_29304_, _29303_, _29300_);
  nor (_29305_, _29304_, _29294_);
  not (_29306_, _29305_);
  and (_29307_, _29306_, _29285_);
  and (_29308_, _29307_, _29272_);
  and (_29309_, _29308_, _29271_);
  and (_29310_, _29309_, _29293_);
  nor (_29311_, _29309_, _29293_);
  or (_29312_, _29311_, _29310_);
  not (_29313_, _29312_);
  and (_29314_, _29305_, _29287_);
  and (_29315_, _29305_, _29286_);
  nor (_29316_, _29315_, _29271_);
  nor (_29317_, _29316_, _29314_);
  not (_29318_, _29317_);
  and (_29319_, _29305_, _29285_);
  and (_29320_, _29305_, _29283_);
  and (_29321_, _29320_, _29274_);
  nor (_29322_, _29321_, _29273_);
  nor (_29323_, _29322_, _29319_);
  not (_29324_, _29323_);
  nor (_29325_, _29320_, _29274_);
  or (_29326_, _29325_, _29321_);
  not (_29327_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_29328_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_29329_, _29305_, _29282_);
  and (_29330_, _29329_, _29328_);
  nor (_29331_, _29330_, _29327_);
  nor (_29332_, _29331_, _29320_);
  not (_29333_, _29332_);
  and (_29334_, _29305_, _29280_);
  and (_29335_, _29334_, _29277_);
  nor (_29336_, _29335_, _29276_);
  nor (_29337_, _29336_, _29329_);
  not (_29338_, _29337_);
  nor (_29339_, _29334_, _29277_);
  or (_29340_, _29339_, _29335_);
  and (_29341_, _29305_, _29279_);
  nor (_29342_, _29341_, _29278_);
  nor (_29343_, _29342_, _29334_);
  not (_29344_, _29343_);
  not (_29345_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_29346_, _29305_, _29345_);
  nor (_29347_, _29305_, _29345_);
  nor (_29348_, _29347_, _29346_);
  not (_29349_, _29348_);
  and (_29350_, _21061_, _20819_);
  not (_29351_, _20567_);
  and (_29352_, _29351_, _20293_);
  and (_29353_, _29352_, _29350_);
  not (_29354_, _21335_);
  and (_29355_, _21576_, _29354_);
  not (_29356_, _21850_);
  and (_29357_, _22091_, _29356_);
  and (_29358_, _29357_, _29355_);
  and (_29359_, _29358_, _29353_);
  and (_29360_, _20819_, _20567_);
  and (_29361_, _29360_, _21061_);
  and (_29362_, _29361_, _20293_);
  not (_29363_, _21576_);
  and (_29364_, _29363_, _21335_);
  and (_29365_, _29364_, _29357_);
  and (_29366_, _29365_, _29362_);
  nor (_29367_, _29366_, _29359_);
  and (_29368_, _29364_, _29362_);
  not (_29369_, _22091_);
  and (_29370_, _29369_, _21850_);
  nor (_29371_, _29370_, _29357_);
  and (_29372_, _29371_, _29368_);
  and (_29373_, _22091_, _21850_);
  and (_29374_, _29373_, _29355_);
  not (_29375_, _29374_);
  not (_29376_, _20819_);
  and (_29377_, _21061_, _29351_);
  and (_29378_, _29377_, _29376_);
  nor (_29379_, _29378_, _29362_);
  nor (_29380_, _29379_, _29375_);
  nor (_29381_, _29380_, _29372_);
  and (_29382_, _29381_, _29367_);
  and (_29383_, _29365_, _29353_);
  and (_29384_, _29355_, _29369_);
  and (_29385_, _29384_, _29353_);
  nor (_29386_, _29385_, _29383_);
  and (_29387_, _29370_, _29355_);
  and (_29388_, _29378_, _20293_);
  and (_29389_, _29388_, _29387_);
  not (_29390_, _21061_);
  nor (_29391_, _21576_, _21335_);
  and (_29392_, _29391_, _29373_);
  and (_29393_, _29392_, _29390_);
  nor (_29394_, _29393_, _29389_);
  and (_29395_, _29394_, _29386_);
  and (_29396_, _29395_, _29382_);
  and (_29397_, _29370_, _29364_);
  and (_29398_, _29397_, _29388_);
  not (_29399_, _29398_);
  and (_29400_, _21576_, _21335_);
  and (_29401_, _29400_, _29371_);
  and (_29402_, _29401_, _29353_);
  not (_29403_, _20293_);
  and (_29404_, _29378_, _29403_);
  and (_29405_, _29404_, _29392_);
  nor (_29406_, _29405_, _29402_);
  and (_29407_, _29406_, _29399_);
  not (_29408_, _29407_);
  not (_29409_, _29362_);
  not (_29410_, _29392_);
  and (_29411_, _29391_, _29357_);
  nor (_29412_, _29397_, _29387_);
  not (_29413_, _29412_);
  nor (_29414_, _29413_, _29411_);
  and (_29415_, _29414_, _29410_);
  nor (_29416_, _29415_, _29409_);
  nor (_29417_, _29416_, _29408_);
  and (_29418_, _29417_, _29396_);
  not (_29420_, _29404_);
  nor (_29421_, _29387_, _29365_);
  nor (_29422_, _29421_, _29420_);
  and (_29423_, _29400_, _22091_);
  and (_29424_, _29423_, _29362_);
  nor (_29425_, _29424_, _29422_);
  not (_29426_, _29397_);
  nor (_29427_, _29353_, _29390_);
  nor (_29428_, _29427_, _29426_);
  not (_29429_, _29428_);
  and (_29431_, _29429_, _29425_);
  and (_29432_, _29374_, _29353_);
  and (_29433_, _29400_, _29370_);
  and (_29434_, _29433_, _29353_);
  nor (_29435_, _29434_, _29432_);
  not (_29436_, _29435_);
  not (_29437_, _29388_);
  and (_29438_, _29373_, _29364_);
  and (_29439_, _29400_, _29369_);
  nor (_29440_, _29439_, _29438_);
  nor (_29442_, _29440_, _29437_);
  nor (_29443_, _29442_, _29436_);
  and (_29444_, _29443_, _29431_);
  nor (_29445_, _22091_, _21850_);
  and (_29446_, _29445_, _29355_);
  nor (_29447_, _29378_, _29361_);
  not (_29448_, _29447_);
  and (_29449_, _29448_, _29446_);
  and (_29450_, _29445_, _29364_);
  nor (_29451_, _29387_, _29450_);
  nor (_29453_, _29451_, _21061_);
  nor (_29454_, _29453_, _29449_);
  not (_29455_, _29353_);
  nor (_29456_, _29369_, _21576_);
  and (_29457_, _29456_, _29354_);
  nor (_29458_, _29457_, _29450_);
  nor (_29459_, _29458_, _29455_);
  and (_29460_, _29404_, _29400_);
  nor (_29461_, _29460_, _29459_);
  and (_29462_, _29461_, _29454_);
  nor (_29464_, _29411_, _29438_);
  nor (_29465_, _29464_, _29420_);
  not (_29466_, _29465_);
  and (_29467_, _29364_, _29356_);
  nor (_29468_, _20819_, _29351_);
  and (_29469_, _29468_, _21061_);
  and (_29470_, _29469_, _29467_);
  and (_29471_, _29469_, _29413_);
  nor (_29472_, _29471_, _29470_);
  and (_29473_, _29365_, _29390_);
  nor (_29475_, _20567_, _20293_);
  and (_29476_, _29475_, _29350_);
  nor (_29477_, _29476_, _29473_);
  and (_29478_, _29477_, _29472_);
  and (_29479_, _29478_, _29466_);
  and (_29480_, _29479_, _29462_);
  and (_29481_, _29480_, _29444_);
  and (_29482_, _29391_, _29370_);
  and (_29483_, _29482_, _29404_);
  nor (_29484_, _29483_, _29358_);
  nor (_29486_, _29484_, _29379_);
  not (_29487_, _29486_);
  and (_29488_, _29404_, _29397_);
  and (_29489_, _29361_, _29403_);
  and (_29490_, _29489_, _29374_);
  nor (_29491_, _29490_, _29488_);
  and (_29492_, _29391_, _29445_);
  and (_29493_, _29492_, _29404_);
  not (_29494_, _29493_);
  and (_29495_, _29489_, _29358_);
  and (_29497_, _29438_, _29353_);
  nor (_29498_, _29497_, _29495_);
  and (_29499_, _29498_, _29494_);
  and (_29500_, _29499_, _29491_);
  and (_29501_, _29500_, _29487_);
  and (_29502_, _29501_, _29481_);
  and (_29503_, _29502_, _29418_);
  not (_29504_, _29503_);
  nor (_29505_, _29298_, _29296_);
  nor (_29506_, _29505_, _29299_);
  nand (_29508_, _29506_, _29504_);
  and (_29509_, _29489_, _29446_);
  or (_29510_, _29468_, _29390_);
  and (_29511_, _29510_, _29397_);
  or (_29512_, _29511_, _29509_);
  nor (_29513_, _29512_, _29434_);
  nand (_29514_, _29513_, _29425_);
  nand (_29515_, _29498_, _29491_);
  or (_29516_, _29515_, _29514_);
  or (_29517_, _29516_, _29408_);
  nor (_29519_, _29517_, _29503_);
  not (_29520_, _29519_);
  nor (_29521_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_29522_, _29521_, _29296_);
  and (_29523_, _29522_, _29520_);
  or (_29524_, _29506_, _29504_);
  and (_29525_, _29524_, _29508_);
  nand (_29526_, _29525_, _29523_);
  and (_29527_, _29526_, _29508_);
  not (_29528_, _29527_);
  and (_29530_, _29303_, _29300_);
  nor (_29531_, _29530_, _29304_);
  and (_29532_, _29531_, _29528_);
  and (_29533_, _29532_, _29349_);
  not (_29534_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_29535_, _29346_, _29534_);
  or (_29536_, _29535_, _29341_);
  and (_29537_, _29536_, _29533_);
  and (_29538_, _29537_, _29344_);
  and (_29539_, _29538_, _29340_);
  and (_29541_, _29539_, _29338_);
  nor (_29542_, _29329_, _29328_);
  or (_29543_, _29542_, _29330_);
  and (_29544_, _29543_, _29541_);
  and (_29545_, _29544_, _29333_);
  and (_29546_, _29545_, _29326_);
  and (_29547_, _29546_, _29324_);
  nor (_29548_, _29319_, _29272_);
  or (_29549_, _29548_, _29315_);
  and (_29550_, _29549_, _29547_);
  and (_29552_, _29550_, _29318_);
  and (_29553_, _29552_, _29313_);
  or (_29554_, _29553_, _29310_);
  nor (_29555_, _29554_, _29291_);
  and (_29556_, _29554_, _29291_);
  or (_29557_, _29556_, _29555_);
  or (_29558_, _29557_, _29268_);
  or (_29559_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_29560_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_29561_, _29560_, _29559_);
  and (_29563_, _29561_, _29558_);
  or (_03164_, _29563_, _29265_);
  nor (_29564_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_03169_, _29564_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_03172_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _27053_);
  nor (_29565_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_29566_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_29567_, _29566_, _29565_);
  nor (_29568_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_29569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_29570_, _29569_, _29568_);
  and (_29571_, _29570_, _29567_);
  nor (_29572_, _29571_, rst);
  and (_29573_, \oc8051_top_1.oc8051_rom1.ea_int , _19854_);
  nand (_29574_, _29573_, _19887_);
  and (_29575_, _29574_, _03172_);
  or (_03175_, _29575_, _29572_);
  and (_29576_, _29571_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_29577_, _29576_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_03178_, _29577_, _27053_);
  nor (_29578_, _29245_, _25561_);
  or (_29579_, _29503_, _20172_);
  nor (_29580_, _29519_, _20029_);
  nand (_29581_, _29503_, _20172_);
  and (_29582_, _29581_, _29579_);
  nand (_29583_, _29582_, _29580_);
  and (_29584_, _29583_, _29579_);
  nor (_29585_, _29584_, _25561_);
  and (_29586_, _29585_, _19986_);
  nor (_29587_, _29585_, _19986_);
  nor (_29588_, _29587_, _29586_);
  nor (_29589_, _29588_, _29578_);
  and (_29590_, _20183_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_29591_, _29590_, _29578_);
  and (_29592_, _29591_, _29517_);
  or (_29593_, _29592_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_29594_, _29593_, _29589_);
  and (_03180_, _29594_, _27053_);
  not (_29595_, _20501_);
  and (_29596_, _21280_, _29595_);
  not (_29597_, _21784_);
  and (_29598_, _21521_, _29597_);
  and (_29599_, _29598_, _29596_);
  and (_29600_, _19887_, _27053_);
  and (_29601_, _29600_, _19876_);
  nand (_29602_, _29601_, _20764_);
  nor (_29603_, _29602_, _21017_);
  not (_29604_, _22047_);
  nor (_29605_, _29604_, _20249_);
  and (_29606_, _29605_, _29603_);
  and (_03188_, _29606_, _29599_);
  nor (_29607_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_29608_, _29607_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_29609_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_03193_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _27053_);
  and (_29610_, _03193_, _29609_);
  or (_03190_, _29610_, _29608_);
  not (_29611_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_29612_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_29613_, _29612_, _29611_);
  and (_29614_, _29612_, _29611_);
  nor (_29615_, _29614_, _29613_);
  not (_29616_, _29615_);
  and (_29617_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_29618_, _29617_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_29619_, _29617_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_29620_, _29619_, _29618_);
  or (_29621_, _29620_, _29612_);
  and (_29622_, _29621_, _29616_);
  nor (_29623_, _29613_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_29624_, _29613_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_29625_, _29624_, _29623_);
  or (_29626_, _29618_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_03199_, _29626_, _27053_);
  and (_29627_, _03199_, _29625_);
  and (_03196_, _29627_, _29622_);
  not (_29628_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_29629_, _29245_, _29628_);
  and (_29630_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_29631_, _29629_);
  and (_29632_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_29633_, _29632_, _29630_);
  and (_03202_, _29633_, _27053_);
  and (_29634_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_29635_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_29636_, _29635_, _29634_);
  and (_03204_, _29636_, _27053_);
  and (_29637_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_29638_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_29639_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _29638_);
  and (_29640_, _29639_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_29641_, _29640_, _29637_);
  and (_03206_, _29641_, _27053_);
  and (_29642_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_29643_, _29642_, _29639_);
  and (_03208_, _29643_, _27053_);
  or (_29644_, _29638_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_03210_, _29644_, _27053_);
  not (_29645_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_29646_, _29645_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_29647_, _29646_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_29648_, _29638_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_29649_, _29648_, _27053_);
  and (_03212_, _29649_, _29647_);
  or (_29650_, _29638_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_03214_, _29650_, _27053_);
  nor (_29651_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_29652_, _29651_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_29653_, _29652_, _27053_);
  and (_29654_, _03193_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_03216_, _29654_, _29653_);
  and (_29655_, _29628_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_29656_, _29655_, _29652_);
  and (_03218_, _29656_, _27053_);
  or (_29657_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  nand (_29658_, _29652_, _24342_);
  and (_29659_, _29658_, _27053_);
  and (_03220_, _29659_, _29657_);
  or (_29660_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_29661_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_29662_, _27788_, _29661_);
  and (_29663_, _29662_, _27053_);
  and (_03604_, _29663_, _29660_);
  or (_29664_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_29665_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_29666_, _27788_, _29665_);
  and (_29667_, _29666_, _27053_);
  and (_03606_, _29667_, _29664_);
  or (_29668_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_29669_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_29670_, _27788_, _29669_);
  and (_29671_, _29670_, _27053_);
  and (_03608_, _29671_, _29668_);
  or (_29672_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_29673_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_29674_, _27788_, _29673_);
  and (_29675_, _29674_, _27053_);
  and (_03610_, _29675_, _29672_);
  or (_29676_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not (_29677_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_29678_, _27788_, _29677_);
  and (_29679_, _29678_, _27053_);
  and (_03612_, _29679_, _29676_);
  or (_29680_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_29681_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_29682_, _27788_, _29681_);
  and (_29683_, _29682_, _27053_);
  and (_03614_, _29683_, _29680_);
  or (_29684_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_29685_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_29686_, _27788_, _29685_);
  and (_29687_, _29686_, _27053_);
  and (_03616_, _29687_, _29684_);
  or (_29688_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_29689_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_29690_, _27788_, _29689_);
  and (_29691_, _29690_, _27053_);
  and (_03618_, _29691_, _29688_);
  or (_29692_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  not (_29693_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nand (_29694_, _27788_, _29693_);
  and (_29695_, _29694_, _27053_);
  and (_03620_, _29695_, _29692_);
  or (_29696_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_29697_, _27788_, _29179_);
  and (_29698_, _29697_, _27053_);
  and (_03622_, _29698_, _29696_);
  or (_29699_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_29700_, _27788_, _29178_);
  and (_29701_, _29700_, _27053_);
  and (_03624_, _29701_, _29699_);
  or (_29702_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_29703_, _27788_, _29183_);
  and (_29704_, _29703_, _27053_);
  and (_03626_, _29704_, _29702_);
  or (_29705_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_29706_, _27788_, _29177_);
  and (_29707_, _29706_, _27053_);
  and (_03628_, _29707_, _29705_);
  or (_29708_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_29709_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_29710_, _29709_, _27053_);
  and (_03630_, _29710_, _29708_);
  or (_29711_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  not (_29712_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_29713_, _27788_, _29712_);
  and (_29714_, _29713_, _27053_);
  and (_03632_, _29714_, _29711_);
  and (_29715_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_29716_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_29717_, _29716_, _29715_);
  and (_03664_, _29717_, _27053_);
  and (_29718_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_29719_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_29720_, _29719_, _29718_);
  and (_03666_, _29720_, _27053_);
  and (_29721_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_29722_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_29723_, _29722_, _29721_);
  and (_03668_, _29723_, _27053_);
  and (_29724_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_29725_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_29726_, _29725_, _29724_);
  and (_03670_, _29726_, _27053_);
  and (_29727_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_29728_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_29729_, _29728_, _29727_);
  and (_03672_, _29729_, _27053_);
  and (_29730_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_29731_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or (_29732_, _29731_, _29730_);
  and (_03674_, _29732_, _27053_);
  and (_29733_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_29734_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or (_29735_, _29734_, _29733_);
  and (_03676_, _29735_, _27053_);
  and (_29736_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_29737_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_29738_, _29737_, _29736_);
  and (_03678_, _29738_, _27053_);
  and (_29739_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_29740_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  or (_29741_, _29740_, _29739_);
  and (_03680_, _29741_, _27053_);
  and (_29742_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_29743_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  or (_29744_, _29743_, _29742_);
  and (_03682_, _29744_, _27053_);
  and (_29745_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_29746_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  or (_29747_, _29746_, _29745_);
  and (_03684_, _29747_, _27053_);
  and (_29748_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_29749_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or (_29750_, _29749_, _29748_);
  and (_03686_, _29750_, _27053_);
  and (_29751_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_29752_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  or (_29753_, _29752_, _29751_);
  and (_03688_, _29753_, _27053_);
  and (_29754_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_29755_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_29756_, _29755_, _29754_);
  and (_03690_, _29756_, _27053_);
  and (_29757_, _27789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and (_29758_, _27788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_29759_, _29758_, _29757_);
  and (_03692_, _29759_, _27053_);
  and (_29760_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_29761_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_29762_, _29761_, _29760_);
  and (_05565_, _29762_, _27053_);
  and (_29763_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_29764_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_29765_, _29764_, _29763_);
  and (_05567_, _29765_, _27053_);
  and (_29766_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_29767_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_29768_, _29767_, _29766_);
  and (_05569_, _29768_, _27053_);
  and (_29769_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_29770_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_29771_, _29770_, _29629_);
  or (_29772_, _29771_, _29769_);
  and (_05571_, _29772_, _27053_);
  and (_29773_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_29774_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_29775_, _29774_, _29773_);
  and (_05573_, _29775_, _27053_);
  and (_29776_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_29777_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_29778_, _29777_, _29776_);
  and (_05575_, _29778_, _27053_);
  and (_29779_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_29780_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_29781_, _29780_, _29779_);
  and (_05577_, _29781_, _27053_);
  and (_29782_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_29783_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or (_29784_, _29783_, _29782_);
  and (_05579_, _29784_, _27053_);
  and (_29785_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_29786_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_29787_, _29786_, _29785_);
  and (_05581_, _29787_, _27053_);
  and (_29788_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_29789_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_29790_, _29789_, _29788_);
  and (_05583_, _29790_, _27053_);
  and (_29791_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_29792_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_29793_, _29792_, _29791_);
  and (_05585_, _29793_, _27053_);
  and (_29794_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_29795_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_29796_, _29795_, _29794_);
  and (_05587_, _29796_, _27053_);
  and (_29797_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_29798_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_29799_, _29798_, _29797_);
  and (_05589_, _29799_, _27053_);
  and (_29800_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_29801_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_29802_, _29801_, _29800_);
  and (_05591_, _29802_, _27053_);
  and (_29803_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_29804_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_29805_, _29804_, _29803_);
  and (_05593_, _29805_, _27053_);
  and (_29806_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_29807_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_29808_, _29807_, _29806_);
  and (_05595_, _29808_, _27053_);
  and (_29809_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_29810_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_29811_, _29810_, _29809_);
  and (_05597_, _29811_, _27053_);
  and (_29812_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_29813_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_29814_, _29813_, _29812_);
  and (_05599_, _29814_, _27053_);
  and (_29815_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_29816_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_29817_, _29816_, _29815_);
  and (_05601_, _29817_, _27053_);
  and (_29818_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_29819_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_29820_, _29819_, _29818_);
  and (_05603_, _29820_, _27053_);
  and (_29821_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_29822_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_29823_, _29822_, _29821_);
  and (_05605_, _29823_, _27053_);
  and (_29824_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_29825_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_29826_, _29825_, _29824_);
  and (_05607_, _29826_, _27053_);
  and (_29827_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_29828_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_29829_, _29828_, _29827_);
  and (_05609_, _29829_, _27053_);
  and (_29830_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_29831_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_29832_, _29831_, _29830_);
  and (_05611_, _29832_, _27053_);
  and (_29833_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_29834_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_29835_, _29834_, _29833_);
  and (_05613_, _29835_, _27053_);
  and (_29836_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_29837_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_29838_, _29837_, _29836_);
  and (_05615_, _29838_, _27053_);
  and (_29839_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_29840_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_29841_, _29840_, _29839_);
  and (_05617_, _29841_, _27053_);
  and (_29842_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_29843_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_29844_, _29843_, _29842_);
  and (_05619_, _29844_, _27053_);
  and (_29845_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_29846_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_29847_, _29846_, _29845_);
  and (_05621_, _29847_, _27053_);
  and (_29848_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_29849_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_29850_, _29849_, _29848_);
  and (_05623_, _29850_, _27053_);
  and (_29851_, _29629_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_29852_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_29853_, _29852_, _29851_);
  and (_05625_, _29853_, _27053_);
  and (_05628_, _20315_, _27053_);
  and (_05631_, _20589_, _27053_);
  and (_05634_, _20841_, _27053_);
  nor (_05636_, _25585_, rst);
  nor (_05639_, _25688_, rst);
  nor (_05642_, _25879_, rst);
  nor (_05645_, _25777_, rst);
  nor (_05648_, _25648_, rst);
  nor (_05651_, _25845_, rst);
  nor (_05654_, _25733_, rst);
  nor (_05657_, _25929_, rst);
  and (_05687_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _27053_);
  and (_05689_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _27053_);
  and (_05691_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _27053_);
  and (_05693_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _27053_);
  and (_05695_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _27053_);
  and (_05697_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _27053_);
  and (_05699_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _27053_);
  or (_29854_, _29215_, _29207_);
  nand (_29855_, _29854_, ABINPUT[19]);
  nand (_29856_, _29084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_29857_, _29222_, _25710_);
  and (_29858_, _29085_, _29147_);
  nor (_29859_, _29858_, _29857_);
  not (_29860_, _25620_);
  and (_29861_, _25624_, _29860_);
  nor (_29862_, _25634_, _29861_);
  not (_29863_, _29023_);
  or (_29864_, _29863_, _23280_);
  nor (_29865_, _29864_, _29038_);
  nand (_29866_, _29865_, _29020_);
  and (_29867_, _29866_, _23227_);
  or (_29868_, _29867_, _29862_);
  or (_29869_, _29868_, _29082_);
  and (_29870_, _29869_, _29210_);
  or (_29871_, _29150_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_29872_, _29871_, _29870_);
  or (_29873_, _29872_, _29151_);
  and (_29874_, _29873_, _29859_);
  and (_29875_, _29874_, _29856_);
  and (_29876_, _29875_, _29855_);
  nand (_29877_, _29876_, _29070_);
  or (_29878_, _29070_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_29879_, _29878_, _27053_);
  and (_05701_, _29879_, _29877_);
  and (_29880_, _29854_, ABINPUT[20]);
  and (_29881_, _29222_, _25867_);
  and (_29882_, _29085_, _29141_);
  and (_29883_, _23313_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_29884_, _29883_, _29882_);
  or (_29885_, _29884_, _29881_);
  or (_29886_, _29885_, _29880_);
  nor (_29887_, _29153_, _29151_);
  nor (_29888_, _29887_, _29154_);
  and (_29889_, _29888_, _29870_);
  nor (_29890_, _29889_, _29886_);
  nand (_29891_, _29890_, _29070_);
  or (_29892_, _29070_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_29893_, _29892_, _27053_);
  and (_05703_, _29893_, _29891_);
  and (_29894_, _29084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_29895_, _29854_, ABINPUT[21]);
  and (_29896_, _29222_, _25794_);
  and (_29897_, _29085_, _29135_);
  or (_29898_, _29897_, _29896_);
  or (_29899_, _29898_, _29895_);
  nor (_29900_, _29158_, _29156_);
  nor (_29901_, _29900_, _29159_);
  and (_29902_, _29901_, _29870_);
  or (_29903_, _29902_, _29899_);
  or (_29904_, _29903_, _29894_);
  and (_29905_, _29904_, _29070_);
  not (_29906_, _29070_);
  not (_29907_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_29908_, _29245_, _29907_);
  and (_29909_, _29245_, _29907_);
  nor (_29910_, _29909_, _29908_);
  and (_29911_, _29910_, _29906_);
  or (_29912_, _29911_, _29905_);
  and (_05705_, _29912_, _27053_);
  or (_29913_, _29133_, _29132_);
  or (_29914_, _29913_, _29160_);
  nand (_29915_, _29913_, _29160_);
  and (_29916_, _29915_, _29211_);
  and (_29917_, _29916_, _29914_);
  and (_29918_, _29854_, ABINPUT[22]);
  and (_29919_, _29085_, _29127_);
  and (_29920_, _29222_, _25672_);
  and (_29921_, _23313_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_29922_, _29921_, _29920_);
  or (_29923_, _29922_, _29919_);
  or (_29924_, _29923_, _29918_);
  or (_29925_, _29924_, _29917_);
  and (_29926_, _29925_, _29070_);
  and (_29927_, _29908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_29928_, _29908_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_29929_, _29928_, _29927_);
  and (_29930_, _29929_, _29906_);
  or (_29931_, _29930_, _29926_);
  and (_05707_, _29931_, _27053_);
  and (_29932_, _29084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_29933_, _29854_, ABINPUT[23]);
  and (_29934_, _29085_, _29120_);
  and (_29935_, _29222_, _25829_);
  or (_29936_, _29935_, _29934_);
  or (_29937_, _29936_, _29933_);
  or (_29938_, _29937_, _29932_);
  or (_29939_, _29164_, _29162_);
  and (_29940_, _29939_, _29165_);
  and (_29941_, _29940_, _29870_);
  or (_29942_, _29941_, _29938_);
  and (_29943_, _29942_, _29070_);
  and (_29944_, _29908_, _29247_);
  nor (_29945_, _29927_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_29946_, _29945_, _29944_);
  nor (_29947_, _29946_, _29070_);
  or (_29948_, _29947_, _29943_);
  and (_05709_, _29948_, _27053_);
  and (_29949_, _29084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_29950_, _29854_, ABINPUT[24]);
  and (_29951_, _29085_, _29112_);
  and (_29952_, _29222_, _25757_);
  or (_29953_, _29952_, _29951_);
  or (_29954_, _29953_, _29950_);
  or (_29955_, _29954_, _29949_);
  or (_29956_, _29119_, _29117_);
  nand (_29957_, _29956_, _29166_);
  or (_29958_, _29956_, _29166_);
  and (_29959_, _29958_, _29957_);
  and (_29960_, _29959_, _29870_);
  or (_29961_, _29960_, _29955_);
  and (_29962_, _29961_, _29070_);
  and (_29963_, _29944_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_29964_, _29944_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_29965_, _29964_, _29963_);
  nor (_29966_, _29965_, _29070_);
  or (_29967_, _29966_, _29962_);
  and (_05711_, _29967_, _27053_);
  and (_29968_, _29084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_29969_, _29854_, ABINPUT[25]);
  and (_29970_, _29085_, _29103_);
  and (_29971_, _29222_, _25915_);
  or (_29972_, _29971_, _29970_);
  or (_29973_, _29972_, _29969_);
  or (_29974_, _29973_, _29968_);
  nor (_29975_, _29168_, _29111_);
  nor (_29976_, _29975_, _29169_);
  and (_29977_, _29976_, _29870_);
  or (_29978_, _29977_, _29974_);
  and (_29979_, _29978_, _29070_);
  and (_29980_, _29963_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_29981_, _29963_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_29982_, _29981_, _29980_);
  nor (_29983_, _29982_, _29070_);
  or (_29984_, _29983_, _29979_);
  and (_05713_, _29984_, _27053_);
  and (_29985_, _29084_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_29986_, _29854_, ABINPUT[26]);
  and (_29987_, _29085_, _29073_);
  and (_29988_, _29222_, _25578_);
  or (_29989_, _29988_, _29987_);
  or (_29990_, _29989_, _29986_);
  or (_29991_, _29990_, _29985_);
  or (_29992_, _29100_, _29101_);
  nand (_29993_, _29992_, _29170_);
  or (_29994_, _29992_, _29170_);
  and (_29995_, _29994_, _29993_);
  and (_29996_, _29995_, _29211_);
  or (_29997_, _29996_, _29991_);
  and (_29998_, _29997_, _29070_);
  or (_29999_, _29980_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_30000_, _29252_, _29070_);
  and (_30001_, _30000_, _29999_);
  or (_30002_, _30001_, _29998_);
  and (_05715_, _30002_, _27053_);
  and (_30003_, _29172_, _29693_);
  nor (_30004_, _29172_, _29693_);
  nor (_30005_, _30004_, _30003_);
  or (_30006_, _30005_, _29096_);
  nand (_30007_, _30005_, _29096_);
  and (_30008_, _30007_, _29211_);
  and (_30009_, _30008_, _30006_);
  and (_30010_, _29215_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_30011_, _29207_, ABINPUT[11]);
  and (_30012_, _23313_, ABINPUT[19]);
  or (_30013_, _30012_, _30011_);
  nor (_30014_, _30013_, _30010_);
  and (_30015_, _29085_, _25710_);
  and (_30016_, _29222_, _29369_);
  nor (_30017_, _30016_, _30015_);
  and (_30018_, _30017_, _30014_);
  nand (_30019_, _30018_, _29070_);
  or (_30020_, _30019_, _30009_);
  nor (_30021_, _29252_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_30022_, _30021_, _29253_);
  or (_30023_, _30022_, _29070_);
  and (_30024_, _30023_, _27053_);
  and (_05717_, _30024_, _30020_);
  and (_30025_, _29172_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_30026_, _30025_, _29096_);
  and (_30027_, _29180_, _29095_);
  nor (_30028_, _30027_, _30026_);
  nand (_30029_, _30028_, _29179_);
  or (_30030_, _30028_, _29179_);
  and (_30031_, _30030_, _29211_);
  and (_30032_, _30031_, _30029_);
  and (_30033_, _29215_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_30034_, _29207_, ABINPUT[12]);
  and (_30035_, _23313_, ABINPUT[20]);
  or (_30036_, _30035_, _30034_);
  nor (_30037_, _30036_, _30033_);
  and (_30038_, _29085_, _25867_);
  and (_30039_, _29222_, _29354_);
  nor (_30040_, _30039_, _30038_);
  and (_30041_, _30040_, _30037_);
  nand (_30042_, _30041_, _29070_);
  or (_30043_, _30042_, _30032_);
  and (_30044_, _29251_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_30045_, _30044_, _29246_);
  nor (_30046_, _30045_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_30047_, _30045_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_30048_, _30047_, _30046_);
  or (_30049_, _30048_, _29070_);
  and (_30050_, _30049_, _27053_);
  and (_05719_, _30050_, _30043_);
  and (_30051_, _29181_, _29095_);
  and (_30052_, _30026_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_30053_, _30052_, _30051_);
  nand (_30054_, _30053_, _29178_);
  or (_30055_, _30053_, _29178_);
  and (_30056_, _30055_, _29211_);
  and (_30057_, _30056_, _30054_);
  and (_30058_, _29215_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_30059_, _29207_, ABINPUT[13]);
  and (_30060_, _23313_, ABINPUT[21]);
  or (_30061_, _30060_, _30059_);
  nor (_30062_, _30061_, _30058_);
  and (_30063_, _29085_, _25794_);
  and (_30064_, _29222_, _29363_);
  nor (_30065_, _30064_, _30063_);
  and (_30066_, _30065_, _30062_);
  nand (_30067_, _30066_, _29070_);
  or (_30068_, _30067_, _30057_);
  nor (_30069_, _30047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_30070_, _30047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_30071_, _30070_, _30069_);
  or (_30072_, _30071_, _29070_);
  and (_30073_, _30072_, _27053_);
  and (_05721_, _30073_, _30068_);
  and (_30074_, _29173_, _29096_);
  and (_30075_, _29182_, _29095_);
  nor (_30076_, _30075_, _30074_);
  nand (_30077_, _30076_, _29183_);
  or (_30078_, _30076_, _29183_);
  and (_30079_, _30078_, _29211_);
  and (_30080_, _30079_, _30077_);
  nor (_30081_, _29229_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_30082_, _30081_, _29230_);
  and (_30083_, _30082_, _29222_);
  and (_30084_, _29215_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_30085_, _30084_, _30083_);
  and (_30086_, _29085_, _25672_);
  and (_30087_, _29207_, ABINPUT[14]);
  and (_30088_, _23313_, ABINPUT[22]);
  or (_30089_, _30088_, _30087_);
  or (_30090_, _30089_, _30086_);
  nor (_30091_, _30090_, _30085_);
  nand (_30092_, _30091_, _29070_);
  or (_30093_, _30092_, _30080_);
  nor (_30094_, _30070_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_30095_, _30094_, _29255_);
  or (_30096_, _30095_, _29070_);
  and (_30097_, _30096_, _27053_);
  and (_05723_, _30097_, _30093_);
  nor (_30098_, _29185_, _29175_);
  nand (_30099_, _30098_, _29177_);
  or (_30100_, _30098_, _29177_);
  and (_30101_, _30100_, _29211_);
  and (_30102_, _30101_, _30099_);
  and (_30103_, _29215_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_30104_, _29207_, ABINPUT[15]);
  and (_30105_, _23313_, ABINPUT[23]);
  or (_30106_, _30105_, _30104_);
  nor (_30107_, _30106_, _30103_);
  nor (_30108_, _29230_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_30109_, _30108_, _29231_);
  and (_30110_, _30109_, _29222_);
  and (_30111_, _29085_, _25829_);
  nor (_30112_, _30111_, _30110_);
  and (_30113_, _30112_, _30107_);
  nand (_30114_, _30113_, _29070_);
  or (_30115_, _30114_, _30102_);
  nor (_30116_, _29255_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_30117_, _30116_, _29256_);
  or (_30118_, _30117_, _29070_);
  and (_30119_, _30118_, _27053_);
  and (_05725_, _30119_, _30115_);
  and (_30120_, _29215_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_30121_, _29085_, _25757_);
  and (_30122_, _29084_, ABINPUT[24]);
  or (_30123_, _30122_, _30121_);
  or (_30124_, _30123_, _30120_);
  nor (_30125_, _29187_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_30126_, _29187_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_30127_, _30126_, _30125_);
  and (_30128_, _30127_, _29870_);
  or (_30129_, _30128_, _30124_);
  nor (_30130_, _29231_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_30131_, _30130_, _29232_);
  and (_30132_, _30131_, _29222_);
  and (_30133_, _29207_, ABINPUT[16]);
  nor (_30134_, _30133_, _30132_);
  nand (_30135_, _30134_, _29070_);
  or (_30136_, _30135_, _30129_);
  nor (_30137_, _29256_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_30138_, _30137_, _29257_);
  or (_30139_, _30138_, _29070_);
  and (_30140_, _30139_, _27053_);
  and (_05727_, _30140_, _30136_);
  nor (_30141_, _29192_, _29712_);
  and (_30142_, _29192_, _29712_);
  or (_30143_, _30142_, _30141_);
  and (_30144_, _30143_, _29211_);
  and (_30145_, _29085_, _25915_);
  and (_30146_, _29207_, ABINPUT[17]);
  and (_30147_, _23313_, ABINPUT[25]);
  or (_30148_, _30147_, _30146_);
  or (_30149_, _30148_, _30145_);
  nor (_30150_, _29232_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_30151_, _30150_, _29233_);
  and (_30152_, _30151_, _29222_);
  and (_30153_, _29215_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_30154_, _30153_, _30152_);
  or (_30155_, _30154_, _30149_);
  or (_30156_, _30155_, _30144_);
  or (_30157_, _30156_, _29906_);
  nor (_30158_, _29257_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_30159_, _30158_, _29258_);
  or (_30160_, _30159_, _29070_);
  and (_30161_, _30160_, _27053_);
  and (_05729_, _30161_, _30157_);
  and (_30162_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_30163_, _29522_, _29520_);
  nor (_30164_, _30163_, _29523_);
  or (_30165_, _30164_, _29268_);
  or (_30166_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_30167_, _30166_, _29560_);
  and (_30168_, _30167_, _30165_);
  or (_05731_, _30168_, _30162_);
  or (_30169_, _29525_, _29523_);
  and (_30170_, _30169_, _29526_);
  or (_30171_, _30170_, _29268_);
  or (_30172_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_30173_, _30172_, _29560_);
  and (_30174_, _30173_, _30171_);
  and (_30175_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_05733_, _30175_, _30174_);
  and (_30176_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_30177_, _29531_, _29528_);
  nor (_30178_, _30177_, _29532_);
  or (_30179_, _30178_, _29268_);
  or (_30180_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_30181_, _30180_, _29560_);
  and (_30182_, _30181_, _30179_);
  or (_05735_, _30182_, _30176_);
  nor (_30183_, _29532_, _29349_);
  nor (_30184_, _30183_, _29533_);
  or (_30185_, _30184_, _29268_);
  or (_30186_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_30187_, _30186_, _29560_);
  and (_30188_, _30187_, _30185_);
  and (_30189_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_05737_, _30189_, _30188_);
  and (_30190_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_30191_, _29536_, _29533_);
  nor (_30192_, _30191_, _29537_);
  or (_30193_, _30192_, _29268_);
  or (_30194_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_30195_, _30194_, _29560_);
  and (_30196_, _30195_, _30193_);
  or (_05739_, _30196_, _30190_);
  and (_30197_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_30198_, _29537_, _29344_);
  nor (_30199_, _30198_, _29538_);
  or (_30200_, _30199_, _29268_);
  or (_30201_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_30202_, _30201_, _29560_);
  and (_30203_, _30202_, _30200_);
  or (_05741_, _30203_, _30197_);
  nor (_30204_, _29538_, _29340_);
  nor (_30205_, _30204_, _29539_);
  or (_30206_, _30205_, _29268_);
  or (_30207_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_30208_, _30207_, _29560_);
  and (_30209_, _30208_, _30206_);
  and (_30210_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_05743_, _30210_, _30209_);
  nor (_30211_, _29539_, _29338_);
  nor (_30212_, _30211_, _29541_);
  or (_30213_, _30212_, _29268_);
  or (_30214_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_30215_, _30214_, _29560_);
  and (_30216_, _30215_, _30213_);
  and (_30217_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_05745_, _30217_, _30216_);
  nor (_30218_, _29543_, _29541_);
  nor (_30219_, _30218_, _29544_);
  or (_30220_, _30219_, _29268_);
  or (_30221_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_30222_, _30221_, _29560_);
  and (_30223_, _30222_, _30220_);
  and (_30224_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_05747_, _30224_, _30223_);
  nor (_30225_, _29544_, _29333_);
  nor (_30226_, _30225_, _29545_);
  or (_30227_, _30226_, _29268_);
  or (_30228_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_30229_, _30228_, _29560_);
  and (_30230_, _30229_, _30227_);
  and (_30231_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_05749_, _30231_, _30230_);
  nor (_30232_, _29545_, _29326_);
  nor (_30233_, _30232_, _29546_);
  or (_30234_, _30233_, _29268_);
  or (_30235_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_30236_, _30235_, _29560_);
  and (_30237_, _30236_, _30234_);
  and (_30238_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_05751_, _30238_, _30237_);
  nor (_30239_, _29546_, _29324_);
  nor (_30240_, _30239_, _29547_);
  or (_30241_, _30240_, _29268_);
  or (_30242_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_30243_, _30242_, _29560_);
  and (_30244_, _30243_, _30241_);
  and (_30245_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_05753_, _30245_, _30244_);
  or (_30246_, _29549_, _29547_);
  nor (_30247_, _29268_, _29550_);
  and (_30248_, _30247_, _30246_);
  nor (_30249_, _29267_, _29177_);
  or (_30250_, _30249_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_30251_, _30250_, _30248_);
  or (_30252_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _19854_);
  and (_30253_, _30252_, _27053_);
  and (_05755_, _30253_, _30251_);
  nor (_30254_, _29550_, _29318_);
  nor (_30255_, _30254_, _29552_);
  or (_30256_, _30255_, _29268_);
  or (_30257_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_30258_, _30257_, _29560_);
  and (_30259_, _30258_, _30256_);
  and (_30260_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_05757_, _30260_, _30259_);
  nor (_30261_, _29552_, _29313_);
  nor (_30262_, _30261_, _29553_);
  or (_30263_, _30262_, _29268_);
  or (_30264_, _29267_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_30265_, _30264_, _29560_);
  and (_30266_, _30265_, _30263_);
  and (_30267_, _29264_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_05759_, _30267_, _30266_);
  and (_30268_, _29571_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_30269_, _30268_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_05761_, _30269_, _27053_);
  and (_30270_, _29571_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_30271_, _30270_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_05763_, _30271_, _27053_);
  and (_30272_, _29571_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_30273_, _30272_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_05765_, _30273_, _27053_);
  and (_30274_, _29571_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_30275_, _30274_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_05767_, _30275_, _27053_);
  and (_30276_, _29571_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_30277_, _30276_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_05769_, _30277_, _27053_);
  and (_30278_, _29571_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_30279_, _30278_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_05771_, _30279_, _27053_);
  and (_30280_, _29571_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_30281_, _30280_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_05773_, _30281_, _27053_);
  nor (_30282_, _29519_, _25561_);
  nand (_30283_, _30282_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_30284_, _30282_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30285_, _30284_, _29560_);
  and (_05775_, _30285_, _30283_);
  or (_30286_, _29582_, _29580_);
  and (_30287_, _30286_, _29583_);
  or (_30288_, _30287_, _25561_);
  or (_30289_, _19887_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_30290_, _30289_, _29560_);
  and (_05777_, _30290_, _30288_);
  and (_30291_, _29607_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_30292_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_30293_, _30292_, _03193_);
  or (_05807_, _30293_, _30291_);
  and (_30294_, _29607_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_30295_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_30296_, _30295_, _03193_);
  or (_05809_, _30296_, _30294_);
  and (_30297_, _29607_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_30298_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_30299_, _30298_, _03193_);
  or (_05811_, _30299_, _30297_);
  and (_30300_, _29607_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_30301_, _29770_, _03193_);
  or (_05813_, _30301_, _30300_);
  and (_30302_, _29607_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_30303_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_30304_, _30303_, _03193_);
  or (_05815_, _30304_, _30302_);
  and (_30305_, _29607_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_30306_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_30307_, _30306_, _03193_);
  or (_05817_, _30307_, _30305_);
  and (_30308_, _29607_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_30309_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_30310_, _30309_, _03193_);
  or (_05819_, _30310_, _30308_);
  and (_05821_, _29615_, _27053_);
  nor (_05823_, _29625_, rst);
  and (_05825_, _29621_, _27053_);
  and (_30311_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_30312_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_30313_, _30312_, _30311_);
  and (_05827_, _30313_, _27053_);
  and (_30314_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_30315_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_30316_, _30315_, _30314_);
  and (_05829_, _30316_, _27053_);
  and (_30317_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_30318_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_30319_, _30318_, _30317_);
  and (_05831_, _30319_, _27053_);
  and (_30320_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_30321_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_30322_, _30321_, _30320_);
  and (_05833_, _30322_, _27053_);
  and (_30323_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_30324_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_30325_, _30324_, _30323_);
  and (_05835_, _30325_, _27053_);
  and (_30326_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_30327_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_30328_, _30327_, _30326_);
  and (_05837_, _30328_, _27053_);
  and (_30329_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_30330_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_30331_, _30330_, _30329_);
  and (_05839_, _30331_, _27053_);
  and (_30332_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_30333_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_30334_, _30333_, _30332_);
  and (_05841_, _30334_, _27053_);
  and (_30335_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_30336_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_30337_, _30336_, _30335_);
  and (_05843_, _30337_, _27053_);
  and (_30338_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_30339_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_30340_, _30339_, _30338_);
  and (_05845_, _30340_, _27053_);
  and (_30341_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_30342_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_30343_, _30342_, _30341_);
  and (_05847_, _30343_, _27053_);
  and (_30344_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_30345_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_30346_, _30345_, _30344_);
  and (_05849_, _30346_, _27053_);
  and (_30347_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_30348_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_30349_, _30348_, _30347_);
  and (_05851_, _30349_, _27053_);
  and (_30350_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_30351_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_30352_, _30351_, _30350_);
  and (_05853_, _30352_, _27053_);
  and (_30353_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_30354_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_30355_, _30354_, _30353_);
  and (_05855_, _30355_, _27053_);
  and (_30356_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_30357_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_30358_, _30357_, _30356_);
  and (_05857_, _30358_, _27053_);
  and (_30359_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_30360_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_30361_, _30360_, _30359_);
  and (_05859_, _30361_, _27053_);
  and (_30362_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_30363_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_30364_, _30363_, _30362_);
  and (_05861_, _30364_, _27053_);
  and (_30365_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_30366_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_30367_, _30366_, _30365_);
  and (_05863_, _30367_, _27053_);
  and (_30368_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_30369_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_30370_, _30369_, _30368_);
  and (_05865_, _30370_, _27053_);
  and (_30371_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_30372_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_30373_, _30372_, _30371_);
  and (_05867_, _30373_, _27053_);
  and (_30374_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_30375_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_30376_, _30375_, _30374_);
  and (_05869_, _30376_, _27053_);
  and (_30377_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_30378_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_30379_, _30378_, _30377_);
  and (_05871_, _30379_, _27053_);
  and (_30380_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_30381_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_30382_, _30381_, _30380_);
  and (_05873_, _30382_, _27053_);
  and (_30383_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_30384_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_30385_, _30384_, _30383_);
  and (_05875_, _30385_, _27053_);
  and (_30386_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_30387_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_30388_, _30387_, _30386_);
  and (_05877_, _30388_, _27053_);
  and (_30389_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_30390_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_30391_, _30390_, _30389_);
  and (_05879_, _30391_, _27053_);
  and (_30392_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_30393_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_30394_, _30393_, _30392_);
  and (_05881_, _30394_, _27053_);
  and (_30395_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_30396_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_30397_, _30396_, _30395_);
  and (_05882_, _30397_, _27053_);
  and (_30398_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_30399_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_30400_, _30399_, _30398_);
  and (_05884_, _30400_, _27053_);
  and (_30401_, _29629_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_30402_, _29631_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_30403_, _30402_, _30401_);
  and (_05886_, _30403_, _27053_);
  and (_30404_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_30405_, _29639_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_30406_, _30405_, _30404_);
  and (_05888_, _30406_, _27053_);
  and (_30407_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_30408_, _29639_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_30409_, _30408_, _30407_);
  and (_05890_, _30409_, _27053_);
  and (_30410_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_30411_, _29639_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_30412_, _30411_, _30410_);
  and (_05892_, _30412_, _27053_);
  and (_30413_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_30414_, _29639_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_30415_, _30414_, _30413_);
  and (_05894_, _30415_, _27053_);
  and (_30416_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_30417_, _29639_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_30418_, _30417_, _30416_);
  and (_05896_, _30418_, _27053_);
  and (_30419_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_30420_, _29639_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_30421_, _30420_, _30419_);
  and (_05898_, _30421_, _27053_);
  and (_30422_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_30423_, _29639_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_30424_, _30423_, _30422_);
  and (_05900_, _30424_, _27053_);
  and (_30425_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_30426_, _25688_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_30427_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_30428_, _30427_, _29638_);
  and (_30429_, _30428_, _30426_);
  or (_30430_, _30429_, _30425_);
  and (_05902_, _30430_, _27053_);
  and (_30431_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_30432_, _25879_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_30433_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_30434_, _30433_, _29638_);
  and (_30435_, _30434_, _30432_);
  or (_30436_, _30435_, _30431_);
  and (_05904_, _30436_, _27053_);
  and (_30437_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_30438_, _25777_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_30439_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_30440_, _30439_, _29638_);
  and (_30441_, _30440_, _30438_);
  or (_30442_, _30441_, _30437_);
  and (_05906_, _30442_, _27053_);
  and (_30443_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_30444_, _25648_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_30445_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_30446_, _30445_, _29638_);
  and (_30447_, _30446_, _30444_);
  or (_30448_, _30447_, _30443_);
  and (_05908_, _30448_, _27053_);
  and (_30449_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_30450_, _25845_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_30451_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_30452_, _30451_, _29638_);
  and (_30453_, _30452_, _30450_);
  or (_30454_, _30453_, _30449_);
  and (_05910_, _30454_, _27053_);
  and (_30455_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_30456_, _25733_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_30457_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_30458_, _30457_, _29638_);
  and (_30459_, _30458_, _30456_);
  or (_30460_, _30459_, _30455_);
  and (_05912_, _30460_, _27053_);
  and (_30461_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_30462_, _25929_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_30463_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_30464_, _30463_, _29638_);
  and (_30465_, _30464_, _30462_);
  or (_30466_, _30465_, _30461_);
  and (_05914_, _30466_, _27053_);
  and (_30467_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_30468_, _25610_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_30469_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_30470_, _30469_, _29638_);
  and (_30471_, _30470_, _30468_);
  or (_30472_, _30471_, _30467_);
  and (_05916_, _30472_, _27053_);
  and (_30473_, _29645_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_30474_, _30473_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_30475_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _29638_);
  and (_30476_, _30475_, _27053_);
  and (_05918_, _30476_, _30474_);
  and (_30477_, _29645_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_30478_, _30477_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_30479_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _29638_);
  and (_30480_, _30479_, _27053_);
  and (_05920_, _30480_, _30478_);
  and (_30481_, _29645_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_30482_, _30481_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_30483_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _29638_);
  and (_30484_, _30483_, _27053_);
  and (_05922_, _30484_, _30482_);
  and (_30485_, _29645_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_30486_, _30485_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_30487_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _29638_);
  and (_30488_, _30487_, _27053_);
  and (_05924_, _30488_, _30486_);
  and (_30489_, _29645_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_30490_, _30489_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_30491_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _29638_);
  and (_30492_, _30491_, _27053_);
  and (_05926_, _30492_, _30490_);
  and (_30493_, _29645_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_30494_, _30493_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_30495_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _29638_);
  and (_30496_, _30495_, _27053_);
  and (_05928_, _30496_, _30494_);
  and (_30497_, _29645_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_30498_, _30497_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_30499_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _29638_);
  and (_30500_, _30499_, _27053_);
  and (_05930_, _30500_, _30498_);
  not (_30501_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor (_30502_, _29652_, _30501_);
  and (_30503_, _29652_, ABINPUT[19]);
  or (_30504_, _30503_, _30502_);
  and (_05932_, _30504_, _27053_);
  not (_30505_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nor (_30506_, _29652_, _30505_);
  and (_30507_, _29652_, ABINPUT[20]);
  or (_30508_, _30507_, _30506_);
  and (_05934_, _30508_, _27053_);
  not (_30509_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor (_30510_, _29652_, _30509_);
  and (_30511_, _29652_, ABINPUT[21]);
  or (_30512_, _30511_, _30510_);
  and (_05936_, _30512_, _27053_);
  not (_30513_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor (_30514_, _29652_, _30513_);
  and (_30515_, _29652_, ABINPUT[22]);
  or (_30516_, _30515_, _30514_);
  and (_05938_, _30516_, _27053_);
  or (_30517_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  nand (_30518_, _29652_, _24386_);
  and (_30519_, _30518_, _27053_);
  and (_05940_, _30519_, _30517_);
  or (_30520_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  nand (_30521_, _29652_, _19560_);
  and (_30522_, _30521_, _27053_);
  and (_05942_, _30522_, _30520_);
  or (_30523_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  nand (_30524_, _29652_, _24401_);
  and (_30525_, _30524_, _27053_);
  and (_05944_, _30525_, _30523_);
  or (_30526_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  nand (_30527_, _29652_, _18454_);
  and (_30528_, _30527_, _27053_);
  and (_05946_, _30528_, _30526_);
  or (_30529_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  nand (_30530_, _29652_, _24360_);
  and (_30531_, _30530_, _27053_);
  and (_05948_, _30531_, _30529_);
  or (_30532_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  nand (_30533_, _29652_, _24367_);
  and (_30534_, _30533_, _27053_);
  and (_05950_, _30534_, _30532_);
  or (_30535_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  nand (_30536_, _29652_, _24375_);
  and (_30537_, _30536_, _27053_);
  and (_05952_, _30537_, _30535_);
  or (_30538_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  nand (_30539_, _29652_, _24382_);
  and (_30540_, _30539_, _27053_);
  and (_05954_, _30540_, _30538_);
  or (_30541_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  nand (_30542_, _29652_, _24390_);
  and (_30543_, _30542_, _27053_);
  and (_05956_, _30543_, _30541_);
  or (_30544_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  nand (_30545_, _29652_, _24397_);
  and (_30546_, _30545_, _27053_);
  and (_05958_, _30546_, _30544_);
  or (_30547_, _29652_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  nand (_30548_, _29652_, _24405_);
  and (_30549_, _30548_, _27053_);
  and (_05960_, _30549_, _30547_);
  and (_08268_, _25947_, _27053_);
  and (_08271_, _26031_, _27053_);
  nor (_08277_, _25798_, rst);
  and (_08429_, _26053_, _27053_);
  and (_08431_, _26070_, _27053_);
  and (_08433_, _26086_, _27053_);
  and (_08435_, _26102_, _27053_);
  and (_08437_, _26117_, _27053_);
  and (_08439_, _26132_, _27053_);
  and (_08441_, _26147_, _27053_);
  nor (_08443_, _25714_, rst);
  nor (_08445_, _25888_, rst);
  nor (_12105_, _23983_, rst);
  nand (_30550_, _29600_, _23708_);
  nor (_30551_, _22409_, _21104_);
  or (_12108_, _30551_, _30550_);
  and (_30552_, _29397_, _29378_);
  and (_30553_, _29489_, _29387_);
  and (_30554_, _29391_, _29369_);
  and (_30555_, _30554_, _29361_);
  or (_30556_, _30555_, _30553_);
  or (_30557_, _30556_, _30552_);
  or (_30558_, _29476_, _29424_);
  and (_30559_, _29433_, _29362_);
  or (_30560_, _30559_, _29511_);
  or (_30561_, _30560_, _30558_);
  or (_30562_, _30561_, _30557_);
  nand (_30563_, _29435_, _29406_);
  or (_30564_, _30563_, _30562_);
  and (_30565_, _29388_, _29467_);
  and (_30566_, _29400_, _29445_);
  and (_30567_, _30566_, _29362_);
  and (_30568_, _29456_, _21335_);
  and (_30569_, _29489_, _30568_);
  or (_30570_, _30569_, _30567_);
  and (_30571_, _30554_, _29353_);
  or (_30572_, _30571_, _30570_);
  or (_30573_, _30572_, _30565_);
  nor (_30574_, _29393_, _29359_);
  nand (_30575_, _30574_, _29386_);
  or (_30576_, _30575_, _30573_);
  or (_30577_, _30576_, _30564_);
  and (_30578_, _30577_, _19898_);
  not (_30579_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_30580_, _19876_, _16893_);
  and (_30581_, _30580_, _23206_);
  nor (_30582_, _30581_, _30579_);
  or (_30583_, _30582_, rst);
  or (_12111_, _30583_, _30578_);
  nand (_30584_, _21576_, _19832_);
  or (_30585_, _19832_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_30586_, _30585_, _27053_);
  and (_12114_, _30586_, _30584_);
  and (_30587_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _27053_);
  and (_30588_, _30587_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_30589_, _23598_, _22442_);
  or (_30590_, _30589_, _22881_);
  nor (_30591_, _30590_, _22212_);
  nand (_30592_, _30591_, _29861_);
  and (_30593_, _23873_, _23019_);
  and (_30594_, _22596_, _23598_);
  or (_30595_, _30594_, _30593_);
  and (_30596_, _23598_, _22201_);
  or (_30597_, _30596_, _29035_);
  or (_30598_, _30597_, _23280_);
  or (_30599_, _30598_, _30595_);
  or (_30600_, _30599_, _30592_);
  and (_30601_, _30600_, _29600_);
  or (_12117_, _30601_, _30588_);
  and (_30602_, _22716_, _22409_);
  or (_30603_, _30602_, _23609_);
  and (_30604_, _22793_, _22190_);
  or (_30605_, _30604_, _23675_);
  or (_30606_, _30605_, _23007_);
  or (_30607_, _30606_, _30603_);
  and (_30608_, _30607_, _19887_);
  nor (_30609_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_30610_, _30609_, \oc8051_top_1.oc8051_decoder1.state [0]);
  not (_30611_, _23906_);
  and (_30612_, _30611_, _30610_);
  and (_30613_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_30614_, _30613_, _30612_);
  or (_30615_, _30614_, _30608_);
  and (_12120_, _30615_, _27053_);
  and (_30616_, \oc8051_top_1.oc8051_sfr1.wait_data , _27053_);
  and (_30617_, _30616_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  or (_30618_, _29022_, _27739_);
  and (_30619_, _23873_, _22716_);
  or (_30620_, _30619_, _30618_);
  and (_30621_, _23873_, _23085_);
  or (_30622_, _23096_, _22453_);
  or (_30623_, _30622_, _30621_);
  or (_30624_, _30623_, _22311_);
  nand (_30625_, _29017_, _20326_);
  nand (_30626_, _30625_, _23532_);
  or (_30627_, _30626_, _30603_);
  or (_30628_, _30627_, _30624_);
  or (_30629_, _30628_, _30620_);
  and (_30630_, _30629_, _29600_);
  or (_12123_, _30630_, _30617_);
  and (_30631_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_30632_, _22738_, _19887_);
  or (_30633_, _30632_, _30631_);
  or (_30634_, _30633_, _30612_);
  and (_12126_, _30634_, _27053_);
  and (_30635_, _22585_, _23598_);
  not (_30636_, _23019_);
  nor (_30637_, _30551_, _30636_);
  nor (_30638_, _30637_, _30635_);
  not (_30639_, _30638_);
  and (_30640_, _30639_, _30610_);
  or (_30641_, _30640_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_30642_, _22300_, _21115_);
  and (_30643_, _29044_, _21872_);
  or (_30644_, _30643_, _30642_);
  or (_30645_, _30644_, _30594_);
  and (_30646_, _30644_, _23227_);
  or (_30647_, _30646_, _29079_);
  and (_30648_, _30647_, _30645_);
  or (_30649_, _30648_, _30641_);
  or (_30650_, _16893_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_30651_, _30650_, _27053_);
  and (_12129_, _30651_, _30649_);
  and (_30652_, _30616_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_30653_, _23609_, _22453_);
  and (_30654_, _22387_, _21115_);
  and (_30655_, _22442_, _21104_);
  or (_30656_, _30655_, _22311_);
  or (_30657_, _30656_, _30654_);
  or (_30658_, _30657_, _30653_);
  and (_30659_, _22365_, _22201_);
  or (_30660_, _30604_, _30659_);
  or (_30661_, _22289_, _22190_);
  and (_30662_, _30661_, _27745_);
  or (_30663_, _22300_, _22201_);
  and (_30664_, _30663_, _23041_);
  or (_30665_, _30664_, _30662_);
  or (_30666_, _30665_, _30660_);
  or (_30667_, _30666_, _30658_);
  and (_30668_, _30667_, _29600_);
  or (_12132_, _30668_, _30652_);
  and (_30669_, _30616_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_30670_, _23873_, _22354_);
  or (_30671_, _30670_, _22530_);
  and (_30672_, _23052_, _22179_);
  or (_30673_, _30672_, _23554_);
  and (_30674_, _23041_, _22442_);
  or (_30675_, _30674_, _30673_);
  and (_30676_, _22793_, _22179_);
  and (_30677_, _27741_, _22113_);
  or (_30678_, _30677_, _30676_);
  or (_30679_, _30678_, _23007_);
  and (_30680_, _23598_, _22278_);
  and (_30681_, _22837_, _22267_);
  or (_30682_, _30681_, _30680_);
  or (_30683_, _30682_, _30679_);
  or (_30684_, _30683_, _30675_);
  or (_30685_, _30684_, _30671_);
  and (_30686_, _27740_, _22431_);
  nand (_30687_, _30686_, _27744_);
  or (_30688_, _30687_, _30624_);
  or (_30689_, _30688_, _30685_);
  and (_30690_, _30689_, _29600_);
  or (_12135_, _30690_, _30669_);
  and (_30691_, _27745_, _22585_);
  or (_30692_, _30691_, _23444_);
  and (_30693_, _22672_, _22267_);
  and (_30694_, _22672_, _21082_);
  or (_30695_, _30694_, _23686_);
  or (_30696_, _30695_, _30693_);
  or (_30697_, _30696_, _30692_);
  and (_30698_, _22716_, _22267_);
  or (_30699_, _30698_, _30697_);
  and (_30700_, _30699_, _19887_);
  nand (_30701_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_00010_, _30701_, _23939_);
  or (_00011_, _00010_, _30700_);
  and (_12138_, _00011_, _27053_);
  nand (_00012_, _22859_, _22749_);
  or (_00013_, _30622_, _30642_);
  or (_00014_, _00013_, _00012_);
  or (_00015_, _23010_, _22881_);
  and (_00016_, _22464_, _21872_);
  and (_00017_, _00016_, _22365_);
  and (_00018_, _22596_, _21082_);
  or (_00019_, _00018_, _22508_);
  nor (_00020_, _00019_, _00017_);
  nand (_00021_, _00020_, _22333_);
  or (_00022_, _00021_, _00015_);
  or (_00023_, _00022_, _00014_);
  and (_00024_, _27745_, _22464_);
  or (_00025_, _00024_, _22804_);
  or (_00026_, _00025_, _30605_);
  or (_00027_, _00026_, _27739_);
  and (_00028_, _00016_, _23041_);
  or (_00029_, _00028_, _23510_);
  or (_00030_, _00029_, _23063_);
  or (_00031_, _30643_, _23488_);
  or (_00032_, _00031_, _22629_);
  or (_00033_, _00032_, _00030_);
  or (_00034_, _00033_, _00027_);
  or (_00035_, _00034_, _00023_);
  and (_00036_, _00035_, _19887_);
  and (_00037_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00038_, _30646_, _30612_);
  and (_00039_, _23227_, _23237_);
  or (_00040_, _00039_, _00038_);
  or (_00041_, _00040_, _00037_);
  or (_00042_, _00041_, _00036_);
  and (_12141_, _00042_, _27053_);
  nor (_12189_, _23829_, rst);
  nor (_12191_, _23345_, rst);
  nand (_12194_, _30639_, _29600_);
  nand (_00043_, _30635_, _29600_);
  not (_00045_, _22409_);
  or (_00047_, _30550_, _00045_);
  and (_12197_, _00047_, _00043_);
  or (_00050_, _30559_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_00052_, _00050_, _30570_);
  or (_00054_, _00052_, _30565_);
  and (_00056_, _00054_, _30581_);
  nor (_00057_, _30580_, _23206_);
  or (_00058_, _00057_, rst);
  or (_12200_, _00058_, _00056_);
  nand (_00059_, _20293_, _19832_);
  or (_00060_, _19832_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_00061_, _00060_, _27053_);
  and (_12203_, _00061_, _00059_);
  not (_00063_, _19832_);
  or (_00065_, _20567_, _00063_);
  or (_00066_, _19832_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_00067_, _00066_, _27053_);
  and (_12206_, _00067_, _00065_);
  nand (_00068_, _20819_, _19832_);
  or (_00069_, _19832_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_00070_, _00069_, _27053_);
  and (_12209_, _00070_, _00068_);
  nand (_00071_, _21061_, _19832_);
  or (_00072_, _19832_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_00073_, _00072_, _27053_);
  and (_12212_, _00073_, _00071_);
  or (_00074_, _21850_, _00063_);
  or (_00075_, _19832_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_00076_, _00075_, _27053_);
  and (_12215_, _00076_, _00074_);
  nand (_00077_, _22091_, _19832_);
  or (_00078_, _19832_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_00079_, _00078_, _27053_);
  and (_12218_, _00079_, _00077_);
  nand (_00080_, _21335_, _19832_);
  or (_00081_, _19832_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_00082_, _00081_, _27053_);
  and (_12221_, _00082_, _00080_);
  or (_00083_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _16893_);
  and (_00084_, _00083_, _30641_);
  or (_00085_, _30694_, _27746_);
  or (_00086_, _30677_, _23686_);
  or (_00087_, _30698_, _30693_);
  or (_00089_, _00087_, _00086_);
  or (_00091_, _00089_, _00085_);
  or (_00093_, _30670_, _22376_);
  or (_00095_, _00093_, _30602_);
  not (_00097_, _27738_);
  and (_00099_, _00097_, _23873_);
  or (_00101_, _00099_, _00095_);
  or (_00102_, _00101_, _00091_);
  or (_00103_, _30692_, _30681_);
  and (_00104_, _00016_, _23873_);
  and (_00105_, _23719_, _22793_);
  or (_00106_, _00105_, _00104_);
  or (_00107_, _00106_, _00103_);
  and (_00109_, _23041_, _22618_);
  or (_00110_, _27750_, _00109_);
  or (_00112_, _30680_, _30593_);
  or (_00113_, _00112_, _00110_);
  or (_00114_, _23609_, _23554_);
  or (_00115_, _23730_, _23030_);
  or (_00116_, _00115_, _00114_);
  or (_00117_, _00116_, _00113_);
  or (_00118_, _00117_, _00107_);
  or (_00119_, _00118_, _00102_);
  and (_00120_, _00119_, _19887_);
  or (_00121_, _00120_, _00084_);
  and (_25347_, _00121_, _27053_);
  and (_00122_, _30616_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_00123_, _23873_, _22837_);
  and (_00124_, _22135_, _21082_);
  or (_00125_, _00124_, _23521_);
  or (_00126_, _30678_, _00125_);
  or (_00127_, _00126_, _00123_);
  or (_00128_, _00127_, _23011_);
  and (_00129_, _30635_, _22157_);
  or (_00130_, _00129_, _30593_);
  or (_00131_, _30675_, _00130_);
  or (_00132_, _00131_, _00128_);
  or (_00133_, _30693_, _22848_);
  or (_00134_, _00133_, _22508_);
  and (_00135_, _00134_, _20326_);
  and (_00136_, _23873_, _21872_);
  or (_00137_, _22343_, _22387_);
  and (_00138_, _00137_, _00136_);
  or (_00139_, _00095_, _30619_);
  or (_00141_, _00139_, _00138_);
  or (_00143_, _00141_, _00135_);
  or (_00145_, _00143_, _00132_);
  and (_00147_, _00145_, _29600_);
  or (_25348_, _00147_, _00122_);
  or (_00150_, _00032_, _00023_);
  and (_00152_, _00150_, _19887_);
  and (_00153_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00154_, _00153_, _00040_);
  or (_00155_, _00154_, _00152_);
  and (_25349_, _00155_, _27053_);
  and (_00156_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00157_, _00156_, _00038_);
  and (_00159_, _00157_, _27053_);
  and (_00160_, _22826_, _22157_);
  or (_00162_, _00160_, _23675_);
  or (_00163_, _00162_, _00030_);
  or (_00164_, _00163_, _30644_);
  and (_00165_, _00164_, _29600_);
  or (_25350_, _00165_, _00159_);
  or (_00166_, _30640_, _23950_);
  and (_00167_, _30693_, _22157_);
  or (_00168_, _00167_, _00123_);
  and (_00169_, _22618_, _21115_);
  and (_00170_, _23873_, _22486_);
  or (_00171_, _00170_, _00169_);
  or (_00172_, _00171_, _00168_);
  or (_00173_, _00172_, _30644_);
  or (_00174_, _30691_, _23455_);
  or (_00175_, _27750_, _23895_);
  and (_00176_, _22954_, _22267_);
  or (_00177_, _00176_, _30635_);
  or (_00178_, _00177_, _00175_);
  or (_00179_, _00178_, _00174_);
  or (_00180_, _00179_, _00173_);
  and (_00181_, _23873_, _22201_);
  or (_00182_, _30698_, _30680_);
  or (_00183_, _00182_, _00181_);
  or (_00184_, _00183_, _00085_);
  or (_00185_, _00099_, _23884_);
  or (_00186_, _30593_, _29017_);
  and (_00187_, _00104_, _21598_);
  or (_00188_, _00187_, _00186_);
  or (_00189_, _00188_, _00185_);
  and (_00191_, _00017_, _21598_);
  or (_00193_, _00028_, _23686_);
  or (_00195_, _00193_, _00024_);
  or (_00197_, _30670_, _23631_);
  or (_00199_, _00197_, _00195_);
  or (_00201_, _00199_, _00191_);
  or (_00203_, _00201_, _00189_);
  or (_00204_, _00203_, _00184_);
  or (_00205_, _00204_, _00180_);
  and (_00206_, _00205_, _19887_);
  or (_00207_, _00206_, _00166_);
  and (_00208_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_00209_, _00208_, _00207_);
  and (_25351_, _00209_, _27053_);
  nand (_00211_, _23642_, _22705_);
  or (_00213_, _22837_, _22354_);
  and (_00214_, _00213_, _23598_);
  or (_00215_, _00028_, _00024_);
  and (_00216_, _00215_, _21598_);
  or (_00217_, _00216_, _00214_);
  or (_00218_, _00217_, _00211_);
  or (_00219_, _00017_, _22629_);
  or (_00220_, _30602_, _23686_);
  or (_00221_, _00220_, _23895_);
  or (_00222_, _00221_, _00219_);
  or (_00223_, _00222_, _00174_);
  or (_00224_, _00223_, _00218_);
  or (_00225_, _00189_, _00184_);
  or (_00226_, _00225_, _00224_);
  and (_00227_, _00226_, _19887_);
  or (_00228_, _00227_, _00166_);
  and (_00229_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or (_00230_, _00229_, _00228_);
  and (_25352_, _00230_, _27053_);
  and (_00231_, _30616_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_00232_, _23598_, _22300_);
  or (_00233_, _00232_, _30589_);
  and (_00234_, _00136_, _30661_);
  or (_00235_, _00234_, _22322_);
  or (_00236_, _00235_, _00015_);
  or (_00237_, _00236_, _00233_);
  not (_00238_, _25629_);
  and (_00239_, _22954_, _21093_);
  or (_00240_, _30698_, _23686_);
  or (_00242_, _00240_, _00239_);
  or (_00244_, _00242_, _00238_);
  and (_00246_, _22420_, _22157_);
  or (_00248_, _00246_, _22497_);
  or (_00250_, _30653_, _00248_);
  or (_00252_, _00250_, _00244_);
  and (_00254_, _23598_, _22135_);
  or (_00255_, _00254_, _22727_);
  and (_00256_, _22954_, _23598_);
  or (_00257_, _30691_, _30604_);
  or (_00258_, _00257_, _00256_);
  or (_00259_, _00258_, _00255_);
  or (_00260_, _00259_, _30665_);
  or (_00262_, _00260_, _00252_);
  or (_00263_, _00262_, _00237_);
  and (_00265_, _00263_, _29600_);
  or (_25353_, _00265_, _00231_);
  and (_00266_, _00136_, _22190_);
  or (_00267_, _00266_, _00256_);
  or (_00268_, _00178_, _30671_);
  or (_00269_, _00268_, _00267_);
  nand (_00270_, _23466_, _22639_);
  or (_00271_, _00085_, _00232_);
  or (_00272_, _00271_, _00270_);
  or (_00273_, _30672_, _22376_);
  or (_00274_, _00167_, _30674_);
  or (_00275_, _00274_, _00273_);
  or (_00276_, _30676_, _23609_);
  or (_00277_, _23631_, _23007_);
  or (_00278_, _00277_, _00276_);
  or (_00279_, _00278_, _00275_);
  or (_00280_, _00279_, _00272_);
  or (_00281_, _00280_, _00269_);
  and (_00282_, _00281_, _29600_);
  and (_00283_, _30616_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_00284_, _19843_, _27053_);
  and (_00285_, _00284_, _23895_);
  or (_00286_, _00285_, _00283_);
  or (_25354_, _00286_, _00282_);
  and (_00287_, _22672_, _23598_);
  or (_00288_, _00257_, _00246_);
  nor (_00289_, _00288_, _00287_);
  nand (_00290_, _00289_, _27751_);
  and (_00291_, _22135_, _21104_);
  or (_00293_, _00291_, _00187_);
  or (_00295_, _00293_, _30618_);
  or (_00297_, _00295_, _00290_);
  or (_00299_, _30698_, _23543_);
  not (_00301_, _23697_);
  or (_00303_, _00301_, _23007_);
  or (_00305_, _00303_, _00299_);
  not (_00306_, _27747_);
  or (_00307_, _00186_, _00306_);
  or (_00308_, _00307_, _00305_);
  or (_00309_, _00308_, _30624_);
  or (_00310_, _00309_, _00297_);
  and (_00311_, _00310_, _19887_);
  and (_00313_, _23895_, _16893_);
  and (_00314_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00316_, _00314_, _00313_);
  or (_00317_, _00316_, _00311_);
  and (_25355_, _00317_, _27053_);
  or (_00318_, _00235_, _30660_);
  or (_00319_, _00318_, _00293_);
  nand (_00320_, _27740_, _22639_);
  or (_00321_, _00320_, _00306_);
  or (_00322_, _23675_, _23510_);
  or (_00323_, _00322_, _25628_);
  and (_00324_, _23598_, _22289_);
  or (_00325_, _00324_, _27750_);
  or (_00326_, _00325_, _00323_);
  or (_00327_, _00326_, _30623_);
  or (_00328_, _00327_, _00321_);
  or (_00329_, _00328_, _00319_);
  and (_00330_, _00329_, _29600_);
  and (_00331_, _23884_, _16893_);
  and (_00332_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_00333_, _00332_, _00331_);
  and (_00334_, _00333_, _27053_);
  or (_25356_, _00334_, _00330_);
  and (_00335_, _30616_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_00336_, _30698_, _29017_);
  or (_00337_, _00336_, _22914_);
  or (_00338_, _00337_, _00238_);
  or (_00339_, _00338_, _00248_);
  or (_00340_, _30596_, _00125_);
  or (_00341_, _00340_, _00254_);
  or (_00342_, _00341_, _30697_);
  or (_00344_, _00267_, _00233_);
  or (_00346_, _00344_, _00342_);
  or (_00348_, _00346_, _00339_);
  and (_00350_, _00348_, _29600_);
  or (_25358_, _00350_, _00335_);
  not (_00353_, _27530_);
  nor (_00355_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00356_, _30501_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_00357_, _00356_, _00355_);
  nor (_00358_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00359_, _30505_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_00360_, _00359_, _00358_);
  nor (_00361_, _00360_, _00357_);
  nor (_00363_, _29910_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00364_, _30509_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_00366_, _00364_, _00363_);
  and (_00367_, _00366_, _00361_);
  nor (_00368_, _29929_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_00369_, _30513_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_00370_, _00369_, _00368_);
  and (_00371_, _00370_, _00367_);
  and (_00372_, _00371_, _00353_);
  not (_00373_, _27448_);
  not (_00374_, _00360_);
  nor (_00375_, _00374_, _00357_);
  not (_00376_, _00361_);
  and (_00377_, _00366_, _00376_);
  nor (_00378_, _00366_, _00376_);
  nor (_00379_, _00378_, _00377_);
  and (_00380_, _00370_, _00379_);
  and (_00381_, _00380_, _00375_);
  and (_00382_, _00381_, _00373_);
  not (_00383_, _27489_);
  and (_00384_, _00360_, _00357_);
  and (_00385_, _00380_, _00384_);
  and (_00386_, _00385_, _00383_);
  or (_00387_, _00386_, _00382_);
  not (_00388_, _27366_);
  and (_00389_, _00370_, _00378_);
  and (_00390_, _00389_, _00388_);
  not (_00391_, _27407_);
  and (_00392_, _00374_, _00357_);
  and (_00393_, _00380_, _00392_);
  and (_00394_, _00393_, _00391_);
  or (_00396_, _00394_, _00390_);
  or (_00398_, _00396_, _00387_);
  not (_00400_, _27325_);
  not (_00402_, _00379_);
  and (_00404_, _00370_, _00377_);
  nor (_00406_, _00370_, _00377_);
  nor (_00408_, _00406_, _00404_);
  and (_00409_, _00408_, _00402_);
  and (_00410_, _00409_, _00384_);
  and (_00411_, _00410_, _00400_);
  not (_00412_, _27284_);
  and (_00413_, _00375_, _00409_);
  and (_00414_, _00413_, _00412_);
  or (_00416_, _00414_, _00411_);
  not (_00417_, _27243_);
  and (_00419_, _00409_, _00392_);
  and (_00420_, _00419_, _00417_);
  not (_00421_, _27202_);
  nor (_00422_, _00370_, _00402_);
  and (_00423_, _00422_, _00361_);
  and (_00424_, _00423_, _00421_);
  or (_00425_, _00424_, _00420_);
  or (_00426_, _00425_, _00416_);
  or (_00427_, _00426_, _00398_);
  not (_00428_, _27120_);
  and (_00429_, _00422_, _00375_);
  and (_00430_, _00429_, _00428_);
  not (_00431_, _27161_);
  and (_00432_, _00384_, _00406_);
  and (_00433_, _00432_, _00431_);
  or (_00434_, _00433_, _00430_);
  not (_00435_, _27023_);
  nor (_00436_, _00408_, _00379_);
  and (_00437_, _00436_, _00361_);
  and (_00438_, _00437_, _00435_);
  not (_00439_, _27072_);
  and (_00440_, _00406_, _00392_);
  and (_00441_, _00440_, _00439_);
  or (_00442_, _00441_, _00438_);
  or (_00443_, _00442_, _00434_);
  not (_00444_, _26900_);
  and (_00445_, _00436_, _00392_);
  and (_00446_, _00445_, _00444_);
  not (_00447_, _26982_);
  and (_00449_, _00384_, _00436_);
  and (_00451_, _00449_, _00447_);
  not (_00453_, _26941_);
  and (_00455_, _00375_, _00436_);
  and (_00457_, _00455_, _00453_);
  or (_00459_, _00457_, _00451_);
  or (_00461_, _00459_, _00446_);
  or (_00462_, _00461_, _00443_);
  or (_00463_, _00462_, _00427_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _00463_, _00372_);
  and (_00464_, _00455_, _00353_);
  and (_00465_, _00389_, _00412_);
  and (_00466_, _00393_, _00400_);
  or (_00468_, _00466_, _00465_);
  and (_00469_, _00410_, _00417_);
  and (_00471_, _00413_, _00421_);
  or (_00472_, _00471_, _00469_);
  or (_00473_, _00472_, _00468_);
  and (_00474_, _00385_, _00391_);
  and (_00475_, _00381_, _00388_);
  or (_00476_, _00475_, _00474_);
  and (_00477_, _00445_, _00383_);
  and (_00478_, _00371_, _00373_);
  or (_00479_, _00478_, _00477_);
  or (_00480_, _00479_, _00476_);
  or (_00481_, _00480_, _00473_);
  and (_00482_, _00429_, _00435_);
  and (_00483_, _00432_, _00439_);
  or (_00484_, _00483_, _00482_);
  and (_00485_, _00419_, _00431_);
  and (_00486_, _00423_, _00428_);
  or (_00487_, _00486_, _00485_);
  or (_00488_, _00487_, _00484_);
  and (_00489_, _00449_, _00444_);
  and (_00490_, _00437_, _00453_);
  and (_00491_, _00440_, _00447_);
  or (_00492_, _00491_, _00490_);
  or (_00493_, _00492_, _00489_);
  or (_00494_, _00493_, _00488_);
  or (_00495_, _00494_, _00481_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _00495_, _00464_);
  and (_00496_, _00423_, _00431_);
  and (_00497_, _00432_, _00428_);
  or (_00498_, _00497_, _00496_);
  and (_00500_, _00429_, _00439_);
  and (_00502_, _00440_, _00435_);
  or (_00504_, _00502_, _00500_);
  or (_00506_, _00504_, _00498_);
  and (_00508_, _00455_, _00444_);
  and (_00510_, _00449_, _00453_);
  and (_00512_, _00437_, _00447_);
  or (_00513_, _00512_, _00510_);
  or (_00514_, _00513_, _00508_);
  or (_00515_, _00514_, _00506_);
  and (_00516_, _00371_, _00383_);
  and (_00517_, _00419_, _00421_);
  and (_00518_, _00389_, _00400_);
  and (_00520_, _00410_, _00412_);
  or (_00521_, _00520_, _00518_);
  or (_00523_, _00521_, _00517_);
  and (_00524_, _00445_, _00353_);
  and (_00525_, _00413_, _00417_);
  or (_00526_, _00525_, _00524_);
  and (_00527_, _00385_, _00373_);
  and (_00528_, _00381_, _00391_);
  and (_00529_, _00393_, _00388_);
  or (_00530_, _00529_, _00528_);
  or (_00531_, _00530_, _00527_);
  or (_00532_, _00531_, _00526_);
  or (_00533_, _00532_, _00523_);
  or (_00534_, _00533_, _00516_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _00534_, _00515_);
  and (_00535_, _00449_, _00353_);
  and (_00536_, _00445_, _00373_);
  and (_00537_, _00455_, _00383_);
  or (_00538_, _00537_, _00536_);
  and (_00539_, _00385_, _00388_);
  and (_00540_, _00371_, _00391_);
  or (_00541_, _00540_, _00539_);
  or (_00542_, _00541_, _00538_);
  and (_00543_, _00381_, _00400_);
  and (_00544_, _00393_, _00412_);
  or (_00545_, _00544_, _00543_);
  and (_00546_, _00410_, _00421_);
  and (_00547_, _00389_, _00417_);
  or (_00548_, _00547_, _00546_);
  or (_00549_, _00548_, _00545_);
  or (_00550_, _00549_, _00542_);
  and (_00552_, _00440_, _00453_);
  and (_00554_, _00437_, _00444_);
  and (_00556_, _00429_, _00447_);
  or (_00558_, _00556_, _00554_);
  or (_00560_, _00558_, _00552_);
  and (_00562_, _00423_, _00439_);
  and (_00564_, _00432_, _00435_);
  or (_00565_, _00564_, _00562_);
  and (_00566_, _00419_, _00428_);
  and (_00567_, _00413_, _00431_);
  or (_00568_, _00567_, _00566_);
  or (_00569_, _00568_, _00565_);
  or (_00570_, _00569_, _00560_);
  or (_00572_, _00570_, _00550_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _00572_, _00535_);
  not (_00574_, _27535_);
  and (_00575_, _00455_, _00574_);
  not (_00576_, _27371_);
  and (_00577_, _00381_, _00576_);
  not (_00578_, _27412_);
  and (_00579_, _00385_, _00578_);
  or (_00580_, _00579_, _00577_);
  not (_00581_, _27453_);
  and (_00582_, _00371_, _00581_);
  not (_00583_, _27494_);
  and (_00584_, _00445_, _00583_);
  or (_00585_, _00584_, _00582_);
  or (_00586_, _00585_, _00580_);
  not (_00587_, _27330_);
  and (_00588_, _00393_, _00587_);
  not (_00589_, _27289_);
  and (_00590_, _00389_, _00589_);
  or (_00591_, _00590_, _00588_);
  not (_00592_, _27248_);
  and (_00593_, _00410_, _00592_);
  not (_00594_, _27207_);
  and (_00595_, _00413_, _00594_);
  or (_00596_, _00595_, _00593_);
  or (_00597_, _00596_, _00591_);
  or (_00598_, _00597_, _00586_);
  not (_00599_, _27077_);
  and (_00600_, _00432_, _00599_);
  not (_00601_, _27028_);
  and (_00602_, _00429_, _00601_);
  or (_00604_, _00602_, _00600_);
  not (_00606_, _27166_);
  and (_00608_, _00419_, _00606_);
  not (_00610_, _27125_);
  and (_00612_, _00423_, _00610_);
  or (_00614_, _00612_, _00608_);
  or (_00616_, _00614_, _00604_);
  not (_00617_, _26905_);
  and (_00618_, _00449_, _00617_);
  not (_00619_, _26946_);
  and (_00620_, _00437_, _00619_);
  not (_00621_, _26987_);
  and (_00622_, _00440_, _00621_);
  or (_00624_, _00622_, _00620_);
  or (_00625_, _00624_, _00618_);
  or (_00627_, _00625_, _00616_);
  or (_00628_, _00627_, _00598_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _00628_, _00575_);
  not (_00629_, _27540_);
  and (_00630_, _00455_, _00629_);
  not (_00631_, _27376_);
  and (_00632_, _00381_, _00631_);
  not (_00633_, _27417_);
  and (_00634_, _00385_, _00633_);
  or (_00635_, _00634_, _00632_);
  not (_00636_, _27458_);
  and (_00637_, _00371_, _00636_);
  not (_00638_, _27499_);
  and (_00639_, _00445_, _00638_);
  or (_00640_, _00639_, _00637_);
  or (_00641_, _00640_, _00635_);
  not (_00642_, _27335_);
  and (_00643_, _00393_, _00642_);
  not (_00644_, _27294_);
  and (_00645_, _00389_, _00644_);
  or (_00646_, _00645_, _00643_);
  not (_00647_, _27253_);
  and (_00648_, _00410_, _00647_);
  not (_00649_, _27212_);
  and (_00650_, _00413_, _00649_);
  or (_00651_, _00650_, _00648_);
  or (_00652_, _00651_, _00646_);
  or (_00653_, _00652_, _00641_);
  not (_00654_, _27082_);
  and (_00656_, _00432_, _00654_);
  not (_00658_, _27033_);
  and (_00660_, _00429_, _00658_);
  or (_00662_, _00660_, _00656_);
  not (_00664_, _27171_);
  and (_00666_, _00419_, _00664_);
  not (_00668_, _27130_);
  and (_00669_, _00423_, _00668_);
  or (_00670_, _00669_, _00666_);
  or (_00671_, _00670_, _00662_);
  not (_00672_, _26910_);
  and (_00673_, _00449_, _00672_);
  not (_00674_, _26951_);
  and (_00676_, _00437_, _00674_);
  not (_00677_, _26992_);
  and (_00679_, _00440_, _00677_);
  or (_00680_, _00679_, _00676_);
  or (_00681_, _00680_, _00673_);
  or (_00682_, _00681_, _00671_);
  or (_00683_, _00682_, _00653_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _00683_, _00630_);
  not (_00684_, _27545_);
  and (_00685_, _00455_, _00684_);
  not (_00686_, _27422_);
  and (_00687_, _00385_, _00686_);
  not (_00688_, _27381_);
  and (_00689_, _00381_, _00688_);
  or (_00690_, _00689_, _00687_);
  not (_00691_, _27504_);
  and (_00692_, _00445_, _00691_);
  not (_00693_, _27463_);
  and (_00694_, _00371_, _00693_);
  or (_00695_, _00694_, _00692_);
  or (_00696_, _00695_, _00690_);
  not (_00697_, _27340_);
  and (_00698_, _00393_, _00697_);
  not (_00699_, _27299_);
  and (_00700_, _00389_, _00699_);
  or (_00701_, _00700_, _00698_);
  not (_00702_, _27258_);
  and (_00703_, _00410_, _00702_);
  not (_00704_, _27217_);
  and (_00705_, _00413_, _00704_);
  or (_00706_, _00705_, _00703_);
  or (_00708_, _00706_, _00701_);
  or (_00710_, _00708_, _00696_);
  not (_00712_, _27087_);
  and (_00714_, _00432_, _00712_);
  not (_00716_, _27038_);
  and (_00718_, _00429_, _00716_);
  or (_00720_, _00718_, _00714_);
  not (_00721_, _27176_);
  and (_00722_, _00419_, _00721_);
  not (_00723_, _27135_);
  and (_00724_, _00423_, _00723_);
  or (_00725_, _00724_, _00722_);
  or (_00726_, _00725_, _00720_);
  not (_00728_, _26915_);
  and (_00729_, _00449_, _00728_);
  not (_00731_, _26956_);
  and (_00732_, _00437_, _00731_);
  not (_00733_, _26997_);
  and (_00734_, _00440_, _00733_);
  or (_00735_, _00734_, _00732_);
  or (_00736_, _00735_, _00729_);
  or (_00737_, _00736_, _00726_);
  or (_00738_, _00737_, _00710_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _00738_, _00685_);
  not (_00739_, _27550_);
  and (_00740_, _00455_, _00739_);
  not (_00741_, _27345_);
  and (_00742_, _00393_, _00741_);
  not (_00743_, _27304_);
  and (_00744_, _00389_, _00743_);
  or (_00745_, _00744_, _00742_);
  not (_00746_, _27222_);
  and (_00747_, _00413_, _00746_);
  not (_00748_, _27263_);
  and (_00749_, _00410_, _00748_);
  or (_00750_, _00749_, _00747_);
  or (_00751_, _00750_, _00745_);
  not (_00752_, _27427_);
  and (_00753_, _00385_, _00752_);
  not (_00754_, _27386_);
  and (_00755_, _00381_, _00754_);
  or (_00756_, _00755_, _00753_);
  not (_00757_, _27509_);
  and (_00758_, _00445_, _00757_);
  not (_00760_, _27468_);
  and (_00762_, _00371_, _00760_);
  or (_00764_, _00762_, _00758_);
  or (_00766_, _00764_, _00756_);
  or (_00768_, _00766_, _00751_);
  not (_00770_, _27092_);
  and (_00772_, _00432_, _00770_);
  not (_00773_, _27043_);
  and (_00774_, _00429_, _00773_);
  or (_00775_, _00774_, _00772_);
  not (_00776_, _27181_);
  and (_00777_, _00419_, _00776_);
  not (_00778_, _27140_);
  and (_00780_, _00423_, _00778_);
  or (_00781_, _00780_, _00777_);
  or (_00783_, _00781_, _00775_);
  not (_00784_, _26920_);
  and (_00785_, _00449_, _00784_);
  not (_00786_, _26961_);
  and (_00787_, _00437_, _00786_);
  not (_00788_, _27002_);
  and (_00789_, _00440_, _00788_);
  or (_00790_, _00789_, _00787_);
  or (_00791_, _00790_, _00785_);
  or (_00792_, _00791_, _00783_);
  or (_00793_, _00792_, _00768_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _00793_, _00740_);
  not (_00794_, _27555_);
  and (_00795_, _00455_, _00794_);
  not (_00796_, _27432_);
  and (_00797_, _00385_, _00796_);
  not (_00798_, _27391_);
  and (_00799_, _00381_, _00798_);
  or (_00800_, _00799_, _00797_);
  not (_00801_, _27473_);
  and (_00802_, _00371_, _00801_);
  not (_00803_, _27514_);
  and (_00804_, _00445_, _00803_);
  or (_00805_, _00804_, _00802_);
  or (_00806_, _00805_, _00800_);
  not (_00807_, _27350_);
  and (_00808_, _00393_, _00807_);
  not (_00809_, _27309_);
  and (_00810_, _00389_, _00809_);
  or (_00812_, _00810_, _00808_);
  not (_00814_, _27227_);
  and (_00816_, _00413_, _00814_);
  not (_00818_, _27268_);
  and (_00820_, _00410_, _00818_);
  or (_00822_, _00820_, _00816_);
  or (_00824_, _00822_, _00812_);
  or (_00825_, _00824_, _00806_);
  not (_00826_, _27048_);
  and (_00827_, _00429_, _00826_);
  not (_00828_, _27097_);
  and (_00829_, _00432_, _00828_);
  or (_00830_, _00829_, _00827_);
  not (_00832_, _27186_);
  and (_00833_, _00419_, _00832_);
  not (_00835_, _27145_);
  and (_00836_, _00423_, _00835_);
  or (_00837_, _00836_, _00833_);
  or (_00838_, _00837_, _00830_);
  not (_00839_, _26925_);
  and (_00840_, _00449_, _00839_);
  not (_00841_, _26966_);
  and (_00842_, _00437_, _00841_);
  not (_00843_, _27007_);
  and (_00844_, _00440_, _00843_);
  or (_00845_, _00844_, _00842_);
  or (_00846_, _00845_, _00840_);
  or (_00847_, _00846_, _00838_);
  or (_00848_, _00847_, _00825_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _00848_, _00795_);
  not (_00849_, _27560_);
  and (_00850_, _00455_, _00849_);
  not (_00851_, _27355_);
  and (_00852_, _00393_, _00851_);
  not (_00853_, _27314_);
  and (_00854_, _00389_, _00853_);
  or (_00855_, _00854_, _00852_);
  not (_00856_, _27273_);
  and (_00857_, _00410_, _00856_);
  not (_00858_, _27232_);
  and (_00859_, _00413_, _00858_);
  or (_00860_, _00859_, _00857_);
  or (_00861_, _00860_, _00855_);
  not (_00862_, _27396_);
  and (_00864_, _00381_, _00862_);
  not (_00866_, _27437_);
  and (_00868_, _00385_, _00866_);
  or (_00870_, _00868_, _00864_);
  not (_00872_, _27519_);
  and (_00874_, _00445_, _00872_);
  not (_00876_, _27478_);
  and (_00877_, _00371_, _00876_);
  or (_00878_, _00877_, _00874_);
  or (_00879_, _00878_, _00870_);
  or (_00880_, _00879_, _00861_);
  not (_00881_, _27102_);
  and (_00882_, _00432_, _00881_);
  not (_00883_, _27054_);
  and (_00884_, _00429_, _00883_);
  or (_00885_, _00884_, _00882_);
  not (_00886_, _27191_);
  and (_00887_, _00419_, _00886_);
  not (_00888_, _27150_);
  and (_00889_, _00423_, _00888_);
  or (_00890_, _00889_, _00887_);
  or (_00891_, _00890_, _00885_);
  not (_00892_, _26930_);
  and (_00893_, _00449_, _00892_);
  not (_00894_, _26971_);
  and (_00895_, _00437_, _00894_);
  not (_00896_, _27012_);
  and (_00897_, _00440_, _00896_);
  or (_00898_, _00897_, _00895_);
  or (_00899_, _00898_, _00893_);
  or (_00900_, _00899_, _00891_);
  or (_00901_, _00900_, _00880_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _00901_, _00850_);
  not (_00902_, _27565_);
  and (_00903_, _00455_, _00902_);
  not (_00904_, _27360_);
  and (_00905_, _00393_, _00904_);
  not (_00907_, _27319_);
  and (_00908_, _00389_, _00907_);
  or (_00909_, _00908_, _00905_);
  not (_00911_, _27237_);
  and (_00912_, _00413_, _00911_);
  not (_00913_, _27278_);
  and (_00915_, _00410_, _00913_);
  or (_00916_, _00915_, _00912_);
  or (_00917_, _00916_, _00909_);
  not (_00918_, _27401_);
  and (_00919_, _00381_, _00918_);
  not (_00920_, _27442_);
  and (_00921_, _00385_, _00920_);
  or (_00922_, _00921_, _00919_);
  not (_00923_, _27524_);
  and (_00924_, _00445_, _00923_);
  not (_00925_, _27483_);
  and (_00926_, _00371_, _00925_);
  or (_00927_, _00926_, _00924_);
  or (_00928_, _00927_, _00922_);
  or (_00929_, _00928_, _00917_);
  not (_00930_, _26935_);
  and (_00931_, _00449_, _00930_);
  not (_00932_, _26976_);
  and (_00933_, _00437_, _00932_);
  not (_00934_, _27017_);
  and (_00935_, _00440_, _00934_);
  or (_00936_, _00935_, _00933_);
  or (_00937_, _00936_, _00931_);
  not (_00938_, _27062_);
  and (_00939_, _00429_, _00938_);
  not (_00940_, _27110_);
  and (_00941_, _00432_, _00940_);
  or (_00942_, _00941_, _00939_);
  not (_00943_, _27155_);
  and (_00944_, _00423_, _00943_);
  not (_00945_, _27196_);
  and (_00946_, _00419_, _00945_);
  or (_00947_, _00946_, _00944_);
  or (_00948_, _00947_, _00942_);
  or (_00949_, _00948_, _00937_);
  or (_00950_, _00949_, _00929_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _00950_, _00903_);
  and (_00951_, _00371_, _00574_);
  and (_00952_, _00385_, _00583_);
  and (_00953_, _00381_, _00581_);
  or (_00954_, _00953_, _00952_);
  and (_00955_, _00389_, _00576_);
  and (_00956_, _00393_, _00578_);
  or (_00957_, _00956_, _00955_);
  or (_00958_, _00957_, _00954_);
  and (_00959_, _00410_, _00587_);
  and (_00960_, _00413_, _00589_);
  or (_00961_, _00960_, _00959_);
  and (_00962_, _00419_, _00592_);
  and (_00963_, _00423_, _00594_);
  or (_00964_, _00963_, _00962_);
  or (_00965_, _00964_, _00961_);
  or (_00966_, _00965_, _00958_);
  and (_00967_, _00429_, _00610_);
  and (_00968_, _00432_, _00606_);
  or (_00969_, _00968_, _00967_);
  and (_00970_, _00437_, _00601_);
  and (_00971_, _00440_, _00599_);
  or (_00972_, _00971_, _00970_);
  or (_00973_, _00972_, _00969_);
  and (_00974_, _00445_, _00617_);
  and (_00975_, _00449_, _00621_);
  and (_00976_, _00455_, _00619_);
  or (_00977_, _00976_, _00975_);
  or (_00978_, _00977_, _00974_);
  or (_00979_, _00978_, _00973_);
  or (_00980_, _00979_, _00966_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _00980_, _00951_);
  and (_00981_, _00371_, _00629_);
  and (_00982_, _00381_, _00636_);
  and (_00983_, _00385_, _00638_);
  or (_00984_, _00983_, _00982_);
  and (_00985_, _00389_, _00631_);
  and (_00986_, _00393_, _00633_);
  or (_00987_, _00986_, _00985_);
  or (_00988_, _00987_, _00984_);
  and (_00989_, _00410_, _00642_);
  and (_00990_, _00413_, _00644_);
  or (_00991_, _00990_, _00989_);
  and (_00992_, _00419_, _00647_);
  and (_00993_, _00423_, _00649_);
  or (_00994_, _00993_, _00992_);
  or (_00995_, _00994_, _00991_);
  or (_00996_, _00995_, _00988_);
  and (_00997_, _00429_, _00668_);
  and (_00998_, _00432_, _00664_);
  or (_00999_, _00998_, _00997_);
  and (_01000_, _00437_, _00658_);
  and (_01001_, _00440_, _00654_);
  or (_01002_, _01001_, _01000_);
  or (_01003_, _01002_, _00999_);
  and (_01004_, _00445_, _00672_);
  and (_01005_, _00449_, _00677_);
  and (_01006_, _00455_, _00674_);
  or (_01007_, _01006_, _01005_);
  or (_01008_, _01007_, _01004_);
  or (_01009_, _01008_, _01003_);
  or (_01010_, _01009_, _00996_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _01010_, _00981_);
  and (_01011_, _00371_, _00684_);
  and (_01012_, _00381_, _00693_);
  and (_01013_, _00385_, _00691_);
  or (_01014_, _01013_, _01012_);
  and (_01015_, _00389_, _00688_);
  and (_01016_, _00393_, _00686_);
  or (_01017_, _01016_, _01015_);
  or (_01018_, _01017_, _01014_);
  and (_01019_, _00413_, _00699_);
  and (_01020_, _00410_, _00697_);
  or (_01021_, _01020_, _01019_);
  and (_01022_, _00419_, _00702_);
  and (_01023_, _00423_, _00704_);
  or (_01024_, _01023_, _01022_);
  or (_01025_, _01024_, _01021_);
  or (_01026_, _01025_, _01018_);
  and (_01027_, _00429_, _00723_);
  and (_01028_, _00432_, _00721_);
  or (_01029_, _01028_, _01027_);
  and (_01030_, _00437_, _00716_);
  and (_01031_, _00440_, _00712_);
  or (_01032_, _01031_, _01030_);
  or (_01033_, _01032_, _01029_);
  and (_01034_, _00445_, _00728_);
  and (_01035_, _00455_, _00731_);
  and (_01037_, _00449_, _00733_);
  or (_01038_, _01037_, _01035_);
  or (_01040_, _01038_, _01034_);
  or (_01041_, _01040_, _01033_);
  or (_01043_, _01041_, _01026_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _01043_, _01011_);
  and (_01045_, _00371_, _00739_);
  and (_01046_, _00432_, _00776_);
  and (_01048_, _00429_, _00778_);
  or (_01049_, _01048_, _01046_);
  and (_01051_, _00437_, _00773_);
  and (_01052_, _00440_, _00770_);
  or (_01054_, _01052_, _01051_);
  or (_01055_, _01054_, _01049_);
  and (_01057_, _00445_, _00784_);
  and (_01058_, _00449_, _00788_);
  and (_01060_, _00455_, _00786_);
  or (_01061_, _01060_, _01058_);
  or (_01063_, _01061_, _01057_);
  or (_01064_, _01063_, _01055_);
  and (_01066_, _00410_, _00741_);
  and (_01067_, _00413_, _00743_);
  or (_01069_, _01067_, _01066_);
  and (_01070_, _00419_, _00748_);
  or (_01072_, _01070_, _01069_);
  and (_01073_, _00393_, _00752_);
  and (_01075_, _00423_, _00746_);
  or (_01076_, _01075_, _01073_);
  and (_01078_, _00389_, _00754_);
  and (_01079_, _00381_, _00760_);
  and (_01081_, _00385_, _00757_);
  or (_01082_, _01081_, _01079_);
  or (_01084_, _01082_, _01078_);
  or (_01085_, _01084_, _01076_);
  or (_01087_, _01085_, _01072_);
  or (_01088_, _01087_, _01064_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _01088_, _01045_);
  and (_01090_, _00371_, _00794_);
  and (_01092_, _00381_, _00801_);
  and (_01093_, _00385_, _00803_);
  or (_01095_, _01093_, _01092_);
  and (_01096_, _00393_, _00796_);
  and (_01097_, _00389_, _00798_);
  or (_01098_, _01097_, _01096_);
  or (_01099_, _01098_, _01095_);
  and (_01100_, _00413_, _00809_);
  and (_01101_, _00410_, _00807_);
  or (_01102_, _01101_, _01100_);
  and (_01103_, _00423_, _00814_);
  and (_01104_, _00419_, _00818_);
  or (_01105_, _01104_, _01103_);
  or (_01106_, _01105_, _01102_);
  or (_01107_, _01106_, _01099_);
  and (_01108_, _00429_, _00835_);
  and (_01109_, _00432_, _00832_);
  or (_01110_, _01109_, _01108_);
  and (_01111_, _00437_, _00826_);
  and (_01112_, _00440_, _00828_);
  or (_01113_, _01112_, _01111_);
  or (_01114_, _01113_, _01110_);
  and (_01115_, _00445_, _00839_);
  and (_01116_, _00449_, _00843_);
  and (_01117_, _00455_, _00841_);
  or (_01118_, _01117_, _01116_);
  or (_01119_, _01118_, _01115_);
  or (_01120_, _01119_, _01114_);
  or (_01121_, _01120_, _01107_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _01121_, _01090_);
  and (_01122_, _00371_, _00849_);
  and (_01123_, _00381_, _00876_);
  and (_01124_, _00385_, _00872_);
  or (_01125_, _01124_, _01123_);
  and (_01126_, _00393_, _00866_);
  and (_01127_, _00389_, _00862_);
  or (_01128_, _01127_, _01126_);
  or (_01129_, _01128_, _01125_);
  and (_01130_, _00413_, _00853_);
  and (_01131_, _00410_, _00851_);
  or (_01132_, _01131_, _01130_);
  and (_01133_, _00423_, _00858_);
  and (_01134_, _00419_, _00856_);
  or (_01135_, _01134_, _01133_);
  or (_01136_, _01135_, _01132_);
  or (_01137_, _01136_, _01129_);
  and (_01138_, _00429_, _00888_);
  and (_01139_, _00432_, _00886_);
  or (_01140_, _01139_, _01138_);
  and (_01141_, _00437_, _00883_);
  and (_01142_, _00440_, _00881_);
  or (_01143_, _01142_, _01141_);
  or (_01144_, _01143_, _01140_);
  and (_01145_, _00445_, _00892_);
  and (_01146_, _00449_, _00896_);
  and (_01147_, _00455_, _00894_);
  or (_01148_, _01147_, _01146_);
  or (_01149_, _01148_, _01145_);
  or (_01150_, _01149_, _01144_);
  or (_01151_, _01150_, _01137_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _01151_, _01122_);
  and (_01152_, _00371_, _00902_);
  and (_01153_, _00385_, _00923_);
  and (_01154_, _00381_, _00925_);
  or (_01155_, _01154_, _01153_);
  and (_01156_, _00389_, _00918_);
  and (_01157_, _00393_, _00920_);
  or (_01158_, _01157_, _01156_);
  or (_01159_, _01158_, _01155_);
  and (_01160_, _00413_, _00907_);
  and (_01161_, _00410_, _00904_);
  or (_01162_, _01161_, _01160_);
  and (_01163_, _00423_, _00911_);
  and (_01164_, _00419_, _00913_);
  or (_01165_, _01164_, _01163_);
  or (_01166_, _01165_, _01162_);
  or (_01167_, _01166_, _01159_);
  and (_01168_, _00432_, _00945_);
  and (_01169_, _00429_, _00943_);
  or (_01170_, _01169_, _01168_);
  and (_01171_, _00437_, _00938_);
  and (_01172_, _00440_, _00940_);
  or (_01173_, _01172_, _01171_);
  or (_01174_, _01173_, _01170_);
  and (_01175_, _00445_, _00930_);
  and (_01176_, _00449_, _00934_);
  and (_01177_, _00455_, _00932_);
  or (_01178_, _01177_, _01176_);
  or (_01179_, _01178_, _01175_);
  or (_01180_, _01179_, _01174_);
  or (_01181_, _01180_, _01167_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _01181_, _01152_);
  and (_01182_, _00449_, _00574_);
  and (_01183_, _00445_, _00581_);
  and (_01184_, _00455_, _00583_);
  or (_01185_, _01184_, _01183_);
  and (_01186_, _00385_, _00576_);
  and (_01187_, _00371_, _00578_);
  or (_01188_, _01187_, _01186_);
  or (_01189_, _01188_, _01185_);
  and (_01190_, _00381_, _00587_);
  and (_01191_, _00393_, _00589_);
  or (_01192_, _01191_, _01190_);
  and (_01193_, _00389_, _00592_);
  and (_01194_, _00410_, _00594_);
  or (_01195_, _01194_, _01193_);
  or (_01196_, _01195_, _01192_);
  or (_01197_, _01196_, _01189_);
  and (_01198_, _00440_, _00619_);
  and (_01199_, _00437_, _00617_);
  and (_01200_, _00429_, _00621_);
  or (_01201_, _01200_, _01199_);
  or (_01202_, _01201_, _01198_);
  and (_01203_, _00423_, _00599_);
  and (_01204_, _00432_, _00601_);
  or (_01205_, _01204_, _01203_);
  and (_01206_, _00419_, _00610_);
  and (_01207_, _00413_, _00606_);
  or (_01208_, _01207_, _01206_);
  or (_01209_, _01208_, _01205_);
  or (_01210_, _01209_, _01202_);
  or (_01211_, _01210_, _01197_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _01211_, _01182_);
  and (_01212_, _00449_, _00629_);
  and (_01213_, _00440_, _00674_);
  and (_01214_, _00429_, _00677_);
  and (_01215_, _00437_, _00672_);
  or (_01216_, _01215_, _01214_);
  or (_01217_, _01216_, _01213_);
  and (_01218_, _00423_, _00654_);
  and (_01219_, _00432_, _00658_);
  or (_01220_, _01219_, _01218_);
  and (_01221_, _00419_, _00668_);
  and (_01222_, _00413_, _00664_);
  or (_01223_, _01222_, _01221_);
  or (_01224_, _01223_, _01220_);
  or (_01225_, _01224_, _01217_);
  and (_01226_, _00389_, _00647_);
  and (_01227_, _00410_, _00649_);
  and (_01228_, _00381_, _00642_);
  and (_01229_, _00393_, _00644_);
  or (_01230_, _01229_, _01228_);
  or (_01231_, _01230_, _01227_);
  or (_01232_, _01231_, _01226_);
  and (_01233_, _00455_, _00638_);
  and (_01234_, _00445_, _00636_);
  or (_01235_, _01234_, _01233_);
  and (_01236_, _00385_, _00631_);
  and (_01237_, _00371_, _00633_);
  or (_01238_, _01237_, _01236_);
  or (_01239_, _01238_, _01235_);
  or (_01240_, _01239_, _01232_);
  or (_01241_, _01240_, _01225_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _01241_, _01212_);
  and (_01242_, _00449_, _00684_);
  and (_01243_, _00445_, _00693_);
  and (_01244_, _00455_, _00691_);
  or (_01245_, _01244_, _01243_);
  and (_01246_, _00385_, _00688_);
  and (_01247_, _00371_, _00686_);
  or (_01248_, _01247_, _01246_);
  or (_01249_, _01248_, _01245_);
  and (_01250_, _00381_, _00697_);
  and (_01251_, _00393_, _00699_);
  or (_01252_, _01251_, _01250_);
  and (_01253_, _00410_, _00704_);
  and (_01254_, _00389_, _00702_);
  or (_01255_, _01254_, _01253_);
  or (_01256_, _01255_, _01252_);
  or (_01257_, _01256_, _01249_);
  and (_01258_, _00440_, _00731_);
  and (_01259_, _00437_, _00728_);
  and (_01260_, _00429_, _00733_);
  or (_01261_, _01260_, _01259_);
  or (_01262_, _01261_, _01258_);
  and (_01263_, _00423_, _00712_);
  and (_01264_, _00432_, _00716_);
  or (_01265_, _01264_, _01263_);
  and (_01266_, _00419_, _00723_);
  and (_01267_, _00413_, _00721_);
  or (_01268_, _01267_, _01266_);
  or (_01269_, _01268_, _01265_);
  or (_01270_, _01269_, _01262_);
  or (_01271_, _01270_, _01257_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _01271_, _01242_);
  and (_01272_, _00449_, _00739_);
  and (_01273_, _00440_, _00786_);
  and (_01274_, _00429_, _00788_);
  and (_01275_, _00437_, _00784_);
  or (_01276_, _01275_, _01274_);
  or (_01277_, _01276_, _01273_);
  and (_01278_, _00419_, _00778_);
  and (_01279_, _00413_, _00776_);
  or (_01280_, _01279_, _01278_);
  and (_01281_, _00432_, _00773_);
  and (_01282_, _00423_, _00770_);
  or (_01283_, _01282_, _01281_);
  or (_01284_, _01283_, _01280_);
  or (_01285_, _01284_, _01277_);
  and (_01286_, _00389_, _00748_);
  and (_01287_, _00410_, _00746_);
  and (_01288_, _00393_, _00743_);
  and (_01289_, _00381_, _00741_);
  or (_01290_, _01289_, _01288_);
  or (_01291_, _01290_, _01287_);
  or (_01292_, _01291_, _01286_);
  and (_01293_, _00455_, _00757_);
  and (_01294_, _00445_, _00760_);
  or (_01295_, _01294_, _01293_);
  and (_01296_, _00385_, _00754_);
  and (_01297_, _00371_, _00752_);
  or (_01298_, _01297_, _01296_);
  or (_01299_, _01298_, _01295_);
  or (_01300_, _01299_, _01292_);
  or (_01301_, _01300_, _01285_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _01301_, _01272_);
  and (_01302_, _00449_, _00794_);
  and (_01303_, _00440_, _00841_);
  and (_01304_, _00429_, _00843_);
  and (_01305_, _00437_, _00839_);
  or (_01306_, _01305_, _01304_);
  or (_01307_, _01306_, _01303_);
  and (_01308_, _00423_, _00828_);
  and (_01309_, _00432_, _00826_);
  or (_01310_, _01309_, _01308_);
  and (_01311_, _00419_, _00835_);
  and (_01312_, _00413_, _00832_);
  or (_01313_, _01312_, _01311_);
  or (_01314_, _01313_, _01310_);
  or (_01315_, _01314_, _01307_);
  and (_01316_, _00410_, _00814_);
  and (_01317_, _00381_, _00807_);
  and (_01318_, _00393_, _00809_);
  or (_01319_, _01318_, _01317_);
  and (_01320_, _00389_, _00818_);
  or (_01321_, _01320_, _01319_);
  or (_01322_, _01321_, _01316_);
  and (_01323_, _00445_, _00801_);
  and (_01324_, _00455_, _00803_);
  or (_01325_, _01324_, _01323_);
  and (_01326_, _00385_, _00798_);
  and (_01327_, _00371_, _00796_);
  or (_01328_, _01327_, _01326_);
  or (_01329_, _01328_, _01325_);
  or (_01330_, _01329_, _01322_);
  or (_01331_, _01330_, _01315_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _01331_, _01302_);
  and (_01332_, _00449_, _00849_);
  and (_01333_, _00455_, _00872_);
  and (_01334_, _00445_, _00876_);
  or (_01335_, _01334_, _01333_);
  and (_01336_, _00385_, _00862_);
  and (_01337_, _00371_, _00866_);
  or (_01338_, _01337_, _01336_);
  or (_01339_, _01338_, _01335_);
  and (_01340_, _00393_, _00853_);
  and (_01341_, _00381_, _00851_);
  or (_01342_, _01341_, _01340_);
  and (_01343_, _00410_, _00858_);
  and (_01344_, _00389_, _00856_);
  or (_01345_, _01344_, _01343_);
  or (_01346_, _01345_, _01342_);
  or (_01347_, _01346_, _01339_);
  and (_01348_, _00440_, _00894_);
  and (_01349_, _00437_, _00892_);
  and (_01350_, _00429_, _00896_);
  or (_01351_, _01350_, _01349_);
  or (_01352_, _01351_, _01348_);
  and (_01353_, _00423_, _00881_);
  and (_01354_, _00432_, _00883_);
  or (_01355_, _01354_, _01353_);
  and (_01356_, _00419_, _00888_);
  and (_01357_, _00413_, _00886_);
  or (_01358_, _01357_, _01356_);
  or (_01359_, _01358_, _01355_);
  or (_01360_, _01359_, _01352_);
  or (_01361_, _01360_, _01347_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _01361_, _01332_);
  and (_01362_, _00449_, _00902_);
  and (_01363_, _00445_, _00925_);
  and (_01364_, _00455_, _00923_);
  or (_01365_, _01364_, _01363_);
  and (_01366_, _00385_, _00918_);
  and (_01367_, _00371_, _00920_);
  or (_01368_, _01367_, _01366_);
  or (_01369_, _01368_, _01365_);
  and (_01370_, _00393_, _00907_);
  and (_01371_, _00381_, _00904_);
  or (_01372_, _01371_, _01370_);
  and (_01373_, _00389_, _00913_);
  and (_01374_, _00410_, _00911_);
  or (_01375_, _01374_, _01373_);
  or (_01376_, _01375_, _01372_);
  or (_01377_, _01376_, _01369_);
  and (_01378_, _00440_, _00932_);
  and (_01379_, _00437_, _00930_);
  and (_01380_, _00429_, _00934_);
  or (_01381_, _01380_, _01379_);
  or (_01382_, _01381_, _01378_);
  and (_01383_, _00423_, _00940_);
  and (_01384_, _00432_, _00938_);
  or (_01385_, _01384_, _01383_);
  and (_01386_, _00419_, _00943_);
  and (_01387_, _00413_, _00945_);
  or (_01388_, _01387_, _01386_);
  or (_01389_, _01388_, _01385_);
  or (_01390_, _01389_, _01382_);
  or (_01391_, _01390_, _01377_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _01391_, _01362_);
  and (_01392_, _00445_, _00574_);
  and (_01393_, _00381_, _00578_);
  and (_01394_, _00393_, _00576_);
  or (_01395_, _01394_, _01393_);
  and (_01396_, _00385_, _00581_);
  and (_01397_, _00371_, _00583_);
  or (_01398_, _01397_, _01396_);
  or (_01399_, _01398_, _01395_);
  and (_01400_, _00389_, _00587_);
  and (_01401_, _00410_, _00589_);
  or (_01402_, _01401_, _01400_);
  and (_01403_, _00419_, _00594_);
  and (_01404_, _00413_, _00592_);
  or (_01405_, _01404_, _01403_);
  or (_01406_, _01405_, _01402_);
  or (_01407_, _01406_, _01399_);
  and (_01408_, _00423_, _00606_);
  and (_01409_, _00432_, _00610_);
  or (_01410_, _01409_, _01408_);
  and (_01411_, _00429_, _00599_);
  and (_01412_, _00440_, _00601_);
  or (_01413_, _01412_, _01411_);
  or (_01414_, _01413_, _01410_);
  and (_01415_, _00455_, _00617_);
  and (_01416_, _00449_, _00619_);
  and (_01417_, _00437_, _00621_);
  or (_01418_, _01417_, _01416_);
  or (_01419_, _01418_, _01415_);
  or (_01420_, _01419_, _01414_);
  or (_01421_, _01420_, _01407_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _01421_, _01392_);
  and (_01422_, _00445_, _00629_);
  and (_01423_, _00423_, _00664_);
  and (_01424_, _00432_, _00668_);
  or (_01425_, _01424_, _01423_);
  and (_01426_, _00429_, _00654_);
  and (_01427_, _00440_, _00658_);
  or (_01428_, _01427_, _01426_);
  or (_01429_, _01428_, _01425_);
  and (_01430_, _00455_, _00672_);
  and (_01431_, _00449_, _00674_);
  and (_01432_, _00437_, _00677_);
  or (_01433_, _01432_, _01431_);
  or (_01434_, _01433_, _01430_);
  or (_01435_, _01434_, _01429_);
  and (_01436_, _00393_, _00631_);
  and (_01437_, _00381_, _00633_);
  or (_01438_, _01437_, _01436_);
  and (_01439_, _00385_, _00636_);
  and (_01440_, _00371_, _00638_);
  or (_01441_, _01440_, _01439_);
  or (_01442_, _01441_, _01438_);
  and (_01443_, _00389_, _00642_);
  and (_01444_, _00410_, _00644_);
  or (_01445_, _01444_, _01443_);
  and (_01446_, _00413_, _00647_);
  and (_01447_, _00419_, _00649_);
  or (_01448_, _01447_, _01446_);
  or (_01449_, _01448_, _01445_);
  or (_01450_, _01449_, _01442_);
  or (_01451_, _01450_, _01435_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _01451_, _01422_);
  and (_01452_, _00445_, _00684_);
  and (_01453_, _00423_, _00721_);
  and (_01454_, _00432_, _00723_);
  or (_01455_, _01454_, _01453_);
  and (_01456_, _00429_, _00712_);
  and (_01457_, _00440_, _00716_);
  or (_01458_, _01457_, _01456_);
  or (_01459_, _01458_, _01455_);
  and (_01460_, _00455_, _00728_);
  and (_01461_, _00449_, _00731_);
  and (_01462_, _00437_, _00733_);
  or (_01463_, _01462_, _01461_);
  or (_01464_, _01463_, _01460_);
  or (_01465_, _01464_, _01459_);
  and (_01466_, _00393_, _00688_);
  and (_01467_, _00381_, _00686_);
  or (_01468_, _01467_, _01466_);
  and (_01469_, _00385_, _00693_);
  and (_01470_, _00371_, _00691_);
  or (_01471_, _01470_, _01469_);
  or (_01472_, _01471_, _01468_);
  and (_01473_, _00389_, _00697_);
  and (_01474_, _00410_, _00699_);
  or (_01475_, _01474_, _01473_);
  and (_01476_, _00413_, _00702_);
  and (_01477_, _00419_, _00704_);
  or (_01478_, _01477_, _01476_);
  or (_01479_, _01478_, _01475_);
  or (_01480_, _01479_, _01472_);
  or (_01481_, _01480_, _01465_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _01481_, _01452_);
  and (_01482_, _00445_, _00739_);
  and (_01483_, _00381_, _00752_);
  and (_01484_, _00393_, _00754_);
  or (_01485_, _01484_, _01483_);
  and (_01486_, _00385_, _00760_);
  and (_01487_, _00371_, _00757_);
  or (_01488_, _01487_, _01486_);
  or (_01489_, _01488_, _01485_);
  and (_01490_, _00389_, _00741_);
  and (_01491_, _00410_, _00743_);
  or (_01492_, _01491_, _01490_);
  and (_01493_, _00419_, _00746_);
  and (_01494_, _00413_, _00748_);
  or (_01495_, _01494_, _01493_);
  or (_01496_, _01495_, _01492_);
  or (_01497_, _01496_, _01489_);
  and (_01498_, _00423_, _00776_);
  and (_01499_, _00432_, _00778_);
  or (_01500_, _01499_, _01498_);
  and (_01501_, _00429_, _00770_);
  and (_01502_, _00440_, _00773_);
  or (_01503_, _01502_, _01501_);
  or (_01504_, _01503_, _01500_);
  and (_01505_, _00455_, _00784_);
  and (_01507_, _00449_, _00786_);
  and (_01509_, _00437_, _00788_);
  or (_01511_, _01509_, _01507_);
  or (_01512_, _01511_, _01505_);
  or (_01514_, _01512_, _01504_);
  or (_01515_, _01514_, _01497_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _01515_, _01482_);
  and (_01516_, _00445_, _00794_);
  and (_01517_, _00381_, _00796_);
  and (_01518_, _00393_, _00798_);
  or (_01519_, _01518_, _01517_);
  and (_01520_, _00385_, _00801_);
  and (_01521_, _00371_, _00803_);
  or (_01522_, _01521_, _01520_);
  or (_01523_, _01522_, _01519_);
  and (_01524_, _00389_, _00807_);
  and (_01525_, _00410_, _00809_);
  or (_01526_, _01525_, _01524_);
  and (_01527_, _00413_, _00818_);
  and (_01528_, _00419_, _00814_);
  or (_01529_, _01528_, _01527_);
  or (_01530_, _01529_, _01526_);
  or (_01531_, _01530_, _01523_);
  and (_01532_, _00423_, _00832_);
  and (_01533_, _00432_, _00835_);
  or (_01534_, _01533_, _01532_);
  and (_01535_, _00429_, _00828_);
  and (_01536_, _00440_, _00826_);
  or (_01537_, _01536_, _01535_);
  or (_01538_, _01537_, _01534_);
  and (_01539_, _00455_, _00839_);
  and (_01540_, _00449_, _00841_);
  and (_01541_, _00437_, _00843_);
  or (_01542_, _01541_, _01540_);
  or (_01543_, _01542_, _01539_);
  or (_01544_, _01543_, _01538_);
  or (_01545_, _01544_, _01531_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _01545_, _01516_);
  and (_01546_, _00445_, _00849_);
  and (_01547_, _00393_, _00862_);
  and (_01548_, _00381_, _00866_);
  or (_01549_, _01548_, _01547_);
  and (_01550_, _00371_, _00872_);
  and (_01551_, _00385_, _00876_);
  or (_01552_, _01551_, _01550_);
  or (_01553_, _01552_, _01549_);
  and (_01554_, _00389_, _00851_);
  and (_01555_, _00410_, _00853_);
  or (_01556_, _01555_, _01554_);
  and (_01557_, _00419_, _00858_);
  and (_01558_, _00413_, _00856_);
  or (_01559_, _01558_, _01557_);
  or (_01560_, _01559_, _01556_);
  or (_01561_, _01560_, _01553_);
  and (_01562_, _00423_, _00886_);
  and (_01563_, _00432_, _00888_);
  or (_01564_, _01563_, _01562_);
  and (_01565_, _00429_, _00881_);
  and (_01566_, _00440_, _00883_);
  or (_01567_, _01566_, _01565_);
  or (_01568_, _01567_, _01564_);
  and (_01569_, _00455_, _00892_);
  and (_01570_, _00449_, _00894_);
  and (_01571_, _00437_, _00896_);
  or (_01572_, _01571_, _01570_);
  or (_01573_, _01572_, _01569_);
  or (_01574_, _01573_, _01568_);
  or (_01575_, _01574_, _01561_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _01575_, _01546_);
  and (_01576_, _00445_, _00902_);
  and (_01577_, _00423_, _00945_);
  and (_01578_, _00432_, _00943_);
  or (_01579_, _01578_, _01577_);
  and (_01580_, _00429_, _00940_);
  and (_01581_, _00440_, _00938_);
  or (_01582_, _01581_, _01580_);
  or (_01584_, _01582_, _01579_);
  and (_01585_, _00455_, _00930_);
  and (_01586_, _00449_, _00932_);
  and (_01587_, _00437_, _00934_);
  or (_01588_, _01587_, _01586_);
  or (_01589_, _01588_, _01585_);
  or (_01590_, _01589_, _01584_);
  and (_01591_, _00393_, _00918_);
  and (_01592_, _00381_, _00920_);
  or (_01593_, _01592_, _01591_);
  and (_01594_, _00385_, _00925_);
  and (_01595_, _00371_, _00923_);
  or (_01596_, _01595_, _01594_);
  or (_01597_, _01596_, _01593_);
  and (_01598_, _00389_, _00904_);
  and (_01599_, _00410_, _00907_);
  or (_01600_, _01599_, _01598_);
  and (_01601_, _00413_, _00913_);
  and (_01602_, _00419_, _00911_);
  or (_01603_, _01602_, _01601_);
  or (_01604_, _01603_, _01600_);
  or (_01605_, _01604_, _01597_);
  or (_01606_, _01605_, _01590_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _01606_, _01576_);
  and (_01607_, _27789_, \oc8051_golden_model_1.P3INREG [7]);
  or (_01608_, _01607_, _28182_);
  and (_26389_, _01608_, _27053_);
  and (_01609_, _27789_, \oc8051_golden_model_1.P2INREG [7]);
  or (_01610_, _01609_, _28034_);
  and (_26390_, _01610_, _27053_);
  and (_01611_, _27789_, \oc8051_golden_model_1.P1INREG [7]);
  or (_01612_, _01611_, _27829_);
  and (_26391_, _01612_, _27053_);
  and (_01613_, _27789_, \oc8051_golden_model_1.P0INREG [7]);
  or (_01614_, _01613_, _28148_);
  and (_26392_, _01614_, _27053_);
  nand (_01615_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_01616_, \oc8051_golden_model_1.PC [3]);
  or (_01617_, \oc8051_golden_model_1.PC [2], _01616_);
  or (_01618_, _01617_, _01615_);
  or (_01619_, _01618_, _27381_);
  not (_01620_, \oc8051_golden_model_1.PC [1]);
  or (_01621_, _01620_, \oc8051_golden_model_1.PC [0]);
  or (_01622_, _01621_, _01617_);
  or (_01623_, _01622_, _27340_);
  and (_01624_, _01623_, _01619_);
  not (_01625_, \oc8051_golden_model_1.PC [2]);
  or (_01626_, _01625_, \oc8051_golden_model_1.PC [3]);
  or (_01627_, _01626_, _01615_);
  or (_01628_, _01627_, _27217_);
  or (_01629_, _01626_, _01621_);
  or (_01630_, _01629_, _27176_);
  and (_01631_, _01630_, _01628_);
  and (_01632_, _01631_, _01624_);
  nand (_01633_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_01634_, _01633_, _01615_);
  or (_01635_, _01634_, _27545_);
  or (_01636_, _01633_, _01621_);
  or (_01637_, _01636_, _27504_);
  and (_01638_, _01637_, _01635_);
  or (_01639_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_01640_, _01639_, _01615_);
  or (_01641_, _01640_, _27038_);
  or (_01642_, _01639_, _01621_);
  or (_01643_, _01642_, _26997_);
  and (_01644_, _01643_, _01641_);
  and (_01645_, _01644_, _01638_);
  and (_01646_, _01645_, _01632_);
  not (_01647_, \oc8051_golden_model_1.PC [0]);
  or (_01648_, \oc8051_golden_model_1.PC [1], _01647_);
  or (_01649_, _01648_, _01633_);
  or (_01650_, _01649_, _27463_);
  or (_01651_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_01652_, _01651_, _01633_);
  or (_01653_, _01652_, _27422_);
  and (_01654_, _01653_, _01650_);
  or (_01655_, _01639_, _01651_);
  or (_01656_, _01655_, _26915_);
  or (_01657_, _01639_, _01648_);
  or (_01658_, _01657_, _26956_);
  and (_01659_, _01658_, _01656_);
  and (_01660_, _01659_, _01654_);
  or (_01661_, _01648_, _01617_);
  or (_01662_, _01661_, _27299_);
  or (_01663_, _01651_, _01617_);
  or (_01664_, _01663_, _27258_);
  and (_01665_, _01664_, _01662_);
  or (_01666_, _01648_, _01626_);
  or (_01667_, _01666_, _27135_);
  or (_01668_, _01651_, _01626_);
  or (_01669_, _01668_, _27087_);
  and (_01670_, _01669_, _01667_);
  and (_01671_, _01670_, _01665_);
  and (_01672_, _01671_, _01660_);
  nand (_01673_, _01672_, _01646_);
  or (_01674_, _01618_, _27386_);
  or (_01675_, _01622_, _27345_);
  and (_01676_, _01675_, _01674_);
  or (_01677_, _01627_, _27222_);
  or (_01678_, _01629_, _27181_);
  and (_01679_, _01678_, _01677_);
  and (_01680_, _01679_, _01676_);
  or (_01681_, _01634_, _27550_);
  or (_01682_, _01636_, _27509_);
  and (_01683_, _01682_, _01681_);
  or (_01684_, _01640_, _27043_);
  or (_01685_, _01642_, _27002_);
  and (_01686_, _01685_, _01684_);
  and (_01687_, _01686_, _01683_);
  and (_01688_, _01687_, _01680_);
  or (_01689_, _01649_, _27468_);
  or (_01690_, _01652_, _27427_);
  and (_01691_, _01690_, _01689_);
  or (_01692_, _01655_, _26920_);
  or (_01693_, _01657_, _26961_);
  and (_01694_, _01693_, _01692_);
  and (_01695_, _01694_, _01691_);
  or (_01696_, _01661_, _27304_);
  or (_01697_, _01663_, _27263_);
  and (_01698_, _01697_, _01696_);
  or (_01699_, _01666_, _27140_);
  or (_01700_, _01668_, _27092_);
  and (_01701_, _01700_, _01699_);
  and (_01702_, _01701_, _01698_);
  and (_01703_, _01702_, _01695_);
  nand (_01704_, _01703_, _01688_);
  or (_01705_, _01704_, _01673_);
  or (_01706_, _01618_, _27371_);
  or (_01707_, _01622_, _27330_);
  and (_01708_, _01707_, _01706_);
  or (_01709_, _01627_, _27207_);
  or (_01710_, _01629_, _27166_);
  and (_01711_, _01710_, _01709_);
  and (_01712_, _01711_, _01708_);
  or (_01713_, _01634_, _27535_);
  or (_01714_, _01636_, _27494_);
  and (_01715_, _01714_, _01713_);
  or (_01716_, _01640_, _27028_);
  or (_01717_, _01642_, _26987_);
  and (_01718_, _01717_, _01716_);
  and (_01719_, _01718_, _01715_);
  and (_01720_, _01719_, _01712_);
  or (_01721_, _01649_, _27453_);
  or (_01722_, _01652_, _27412_);
  and (_01723_, _01722_, _01721_);
  or (_01724_, _01655_, _26905_);
  or (_01725_, _01657_, _26946_);
  and (_01726_, _01725_, _01724_);
  and (_01727_, _01726_, _01723_);
  or (_01728_, _01661_, _27289_);
  or (_01729_, _01663_, _27248_);
  and (_01730_, _01729_, _01728_);
  or (_01731_, _01666_, _27125_);
  or (_01732_, _01668_, _27077_);
  and (_01733_, _01732_, _01731_);
  and (_01734_, _01733_, _01730_);
  and (_01735_, _01734_, _01727_);
  and (_01736_, _01735_, _01720_);
  or (_01737_, _01618_, _27376_);
  or (_01738_, _01622_, _27335_);
  and (_01739_, _01738_, _01737_);
  or (_01740_, _01627_, _27212_);
  or (_01741_, _01629_, _27171_);
  and (_01742_, _01741_, _01740_);
  and (_01743_, _01742_, _01739_);
  or (_01744_, _01634_, _27540_);
  or (_01745_, _01636_, _27499_);
  and (_01746_, _01745_, _01744_);
  or (_01747_, _01640_, _27033_);
  or (_01748_, _01642_, _26992_);
  and (_01749_, _01748_, _01747_);
  and (_01750_, _01749_, _01746_);
  and (_01751_, _01750_, _01743_);
  or (_01752_, _01649_, _27458_);
  or (_01753_, _01652_, _27417_);
  and (_01754_, _01753_, _01752_);
  or (_01755_, _01655_, _26910_);
  or (_01756_, _01657_, _26951_);
  and (_01757_, _01756_, _01755_);
  and (_01758_, _01757_, _01754_);
  or (_01759_, _01661_, _27294_);
  or (_01760_, _01663_, _27253_);
  and (_01761_, _01760_, _01759_);
  or (_01762_, _01666_, _27130_);
  or (_01763_, _01668_, _27082_);
  and (_01764_, _01763_, _01762_);
  and (_01765_, _01764_, _01761_);
  and (_01766_, _01765_, _01758_);
  nand (_01767_, _01766_, _01751_);
  or (_01768_, _01767_, _01736_);
  or (_01769_, _01768_, _01705_);
  not (_01770_, _01769_);
  or (_01771_, _01618_, _27401_);
  or (_01772_, _01622_, _27360_);
  and (_01773_, _01772_, _01771_);
  or (_01774_, _01627_, _27237_);
  or (_01775_, _01629_, _27196_);
  and (_01776_, _01775_, _01774_);
  and (_01777_, _01776_, _01773_);
  or (_01778_, _01634_, _27565_);
  or (_01779_, _01636_, _27524_);
  and (_01780_, _01779_, _01778_);
  or (_01781_, _01640_, _27062_);
  or (_01782_, _01642_, _27017_);
  and (_01783_, _01782_, _01781_);
  and (_01784_, _01783_, _01780_);
  and (_01785_, _01784_, _01777_);
  or (_01786_, _01649_, _27483_);
  or (_01787_, _01652_, _27442_);
  and (_01788_, _01787_, _01786_);
  or (_01789_, _01655_, _26935_);
  or (_01790_, _01657_, _26976_);
  and (_01791_, _01790_, _01789_);
  and (_01792_, _01791_, _01788_);
  or (_01793_, _01661_, _27319_);
  or (_01794_, _01663_, _27278_);
  and (_01795_, _01794_, _01793_);
  or (_01796_, _01666_, _27155_);
  or (_01797_, _01668_, _27110_);
  and (_01798_, _01797_, _01796_);
  and (_01799_, _01798_, _01795_);
  and (_01800_, _01799_, _01792_);
  and (_01801_, _01800_, _01785_);
  or (_01802_, _01618_, _27366_);
  or (_01803_, _01622_, _27325_);
  and (_01804_, _01803_, _01802_);
  or (_01805_, _01627_, _27202_);
  or (_01806_, _01629_, _27161_);
  and (_01807_, _01806_, _01805_);
  and (_01808_, _01807_, _01804_);
  or (_01809_, _01634_, _27530_);
  or (_01810_, _01636_, _27489_);
  and (_01811_, _01810_, _01809_);
  or (_01812_, _01640_, _27023_);
  or (_01813_, _01642_, _26982_);
  and (_01814_, _01813_, _01812_);
  and (_01815_, _01814_, _01811_);
  and (_01816_, _01815_, _01808_);
  or (_01817_, _01649_, _27448_);
  or (_01818_, _01652_, _27407_);
  and (_01819_, _01818_, _01817_);
  or (_01820_, _01655_, _26900_);
  or (_01821_, _01657_, _26941_);
  and (_01822_, _01821_, _01820_);
  and (_01823_, _01822_, _01819_);
  or (_01824_, _01661_, _27284_);
  or (_01825_, _01663_, _27243_);
  and (_01826_, _01825_, _01824_);
  or (_01827_, _01666_, _27120_);
  or (_01828_, _01668_, _27072_);
  and (_01829_, _01828_, _01827_);
  and (_01830_, _01829_, _01826_);
  and (_01831_, _01830_, _01823_);
  and (_01832_, _01831_, _01816_);
  and (_01833_, _01832_, _01801_);
  or (_01834_, _01618_, _27391_);
  or (_01835_, _01622_, _27350_);
  and (_01836_, _01835_, _01834_);
  or (_01837_, _01627_, _27227_);
  or (_01838_, _01629_, _27186_);
  and (_01839_, _01838_, _01837_);
  and (_01840_, _01839_, _01836_);
  or (_01841_, _01634_, _27555_);
  or (_01842_, _01636_, _27514_);
  and (_01843_, _01842_, _01841_);
  or (_01844_, _01640_, _27048_);
  or (_01845_, _01642_, _27007_);
  and (_01846_, _01845_, _01844_);
  and (_01847_, _01846_, _01843_);
  and (_01848_, _01847_, _01840_);
  or (_01849_, _01649_, _27473_);
  or (_01850_, _01652_, _27432_);
  and (_01851_, _01850_, _01849_);
  or (_01852_, _01655_, _26925_);
  or (_01853_, _01657_, _26966_);
  and (_01854_, _01853_, _01852_);
  and (_01855_, _01854_, _01851_);
  or (_01856_, _01661_, _27309_);
  or (_01857_, _01663_, _27268_);
  and (_01858_, _01857_, _01856_);
  or (_01859_, _01666_, _27145_);
  or (_01860_, _01668_, _27097_);
  and (_01861_, _01860_, _01859_);
  and (_01862_, _01861_, _01858_);
  and (_01863_, _01862_, _01855_);
  nand (_01864_, _01863_, _01848_);
  or (_01865_, _01618_, _27396_);
  or (_01866_, _01622_, _27355_);
  and (_01867_, _01866_, _01865_);
  or (_01868_, _01627_, _27232_);
  or (_01869_, _01629_, _27191_);
  and (_01870_, _01869_, _01868_);
  and (_01871_, _01870_, _01867_);
  or (_01872_, _01634_, _27560_);
  or (_01873_, _01636_, _27519_);
  and (_01874_, _01873_, _01872_);
  or (_01875_, _01640_, _27054_);
  or (_01876_, _01642_, _27012_);
  and (_01877_, _01876_, _01875_);
  and (_01878_, _01877_, _01874_);
  and (_01879_, _01878_, _01871_);
  or (_01880_, _01649_, _27478_);
  or (_01881_, _01652_, _27437_);
  and (_01882_, _01881_, _01880_);
  or (_01883_, _01655_, _26930_);
  or (_01884_, _01657_, _26971_);
  and (_01885_, _01884_, _01883_);
  and (_01886_, _01885_, _01882_);
  or (_01887_, _01661_, _27314_);
  or (_01888_, _01663_, _27273_);
  and (_01889_, _01888_, _01887_);
  or (_01890_, _01666_, _27150_);
  or (_01891_, _01668_, _27102_);
  and (_01892_, _01891_, _01890_);
  and (_01893_, _01892_, _01889_);
  and (_01894_, _01893_, _01886_);
  and (_01895_, _01894_, _01879_);
  or (_01896_, _01895_, _01864_);
  not (_01897_, _01896_);
  and (_01898_, _01897_, _01833_);
  and (_01899_, _01898_, _01770_);
  not (_01900_, _01634_);
  and (_01901_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_01902_, _01901_, _01900_);
  and (_01903_, _01902_, \oc8051_golden_model_1.PC [6]);
  and (_01904_, _01903_, \oc8051_golden_model_1.PC [7]);
  and (_01905_, _01904_, \oc8051_golden_model_1.PC [8]);
  and (_01906_, _01905_, \oc8051_golden_model_1.PC [9]);
  and (_01907_, _01906_, \oc8051_golden_model_1.PC [10]);
  and (_01908_, _01907_, \oc8051_golden_model_1.PC [11]);
  and (_01909_, _01908_, \oc8051_golden_model_1.PC [12]);
  and (_01910_, _01909_, \oc8051_golden_model_1.PC [13]);
  and (_01911_, _01910_, \oc8051_golden_model_1.PC [14]);
  or (_01912_, _01911_, \oc8051_golden_model_1.PC [15]);
  nand (_01913_, _01911_, \oc8051_golden_model_1.PC [15]);
  and (_01914_, _01913_, _01912_);
  not (_01915_, _01898_);
  not (_01916_, _01673_);
  and (_01917_, _01704_, _01916_);
  nand (_01918_, _01917_, _01767_);
  nor (_01919_, _01918_, _01915_);
  and (_01920_, _01704_, _01673_);
  and (_01921_, _01920_, _01898_);
  nor (_01922_, _01921_, _01919_);
  not (_01923_, _01922_);
  and (_01924_, _01767_, _01673_);
  nor (_01925_, _01924_, _01704_);
  not (_01926_, _01920_);
  nand (_01927_, _01926_, _01918_);
  nor (_01928_, _01927_, _01925_);
  and (_01929_, _01928_, _01898_);
  nor (_01930_, _01929_, _01923_);
  or (_01931_, _01930_, _01914_);
  and (_01932_, _01863_, _01848_);
  or (_01933_, _01895_, _01932_);
  not (_01934_, _01933_);
  and (_01935_, _01934_, _01833_);
  and (_01936_, _01935_, _01770_);
  nand (_01937_, _01894_, _01879_);
  or (_01938_, _01937_, _01864_);
  not (_01939_, _01938_);
  nand (_01940_, _01800_, _01785_);
  and (_01941_, _01832_, _01940_);
  and (_01942_, _01941_, _01939_);
  not (_01943_, _01942_);
  nor (_01944_, _01943_, _01925_);
  not (_01945_, _01944_);
  or (_01946_, _01945_, _01914_);
  nor (_01947_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_01948_, \oc8051_golden_model_1.ACC [6], \oc8051_golden_model_1.ACC [3]);
  and (_01949_, _01948_, _01947_);
  nor (_01950_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [7]);
  nor (_01951_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  and (_01952_, _01951_, _01950_);
  and (_01953_, _01952_, _01949_);
  and (_01954_, _01939_, _01833_);
  and (_01955_, _01954_, _01770_);
  not (_01956_, _01955_);
  and (_01957_, _01942_, _01770_);
  or (_01958_, _01832_, _01940_);
  nor (_01959_, _01958_, _01938_);
  and (_01960_, _01959_, _01770_);
  nor (_01961_, _01960_, _01957_);
  or (_01962_, _01937_, _01932_);
  not (_01963_, _01962_);
  and (_01964_, _01963_, _01941_);
  and (_01965_, _01964_, _01770_);
  and (_01966_, _01941_, _01934_);
  and (_01967_, _01966_, _01770_);
  nor (_01968_, _01967_, _01965_);
  and (_01969_, _01968_, _01961_);
  and (_01970_, _01963_, _01833_);
  and (_01971_, _01970_, _01770_);
  nor (_01972_, _01971_, _01899_);
  and (_01973_, _01941_, _01897_);
  and (_01974_, _01973_, _01770_);
  nor (_01975_, _01974_, _01936_);
  and (_01976_, _01975_, _01972_);
  and (_01977_, _01976_, _01969_);
  and (_01978_, _01977_, _01956_);
  or (_01979_, _01978_, _01620_);
  not (_01980_, _01767_);
  or (_01981_, _01980_, _01736_);
  or (_01982_, _01981_, _01705_);
  nor (_01983_, _01962_, _01958_);
  not (_01984_, _01983_);
  or (_01985_, _01984_, _01982_);
  or (_01986_, _01832_, _01801_);
  or (_01987_, _01986_, _01933_);
  or (_01988_, _01987_, _01769_);
  or (_01989_, _01986_, _01938_);
  or (_01990_, _01989_, _01769_);
  and (_01991_, _01990_, _01988_);
  or (_01992_, _01958_, _01896_);
  or (_01993_, _01992_, _01769_);
  or (_01994_, _01986_, _01962_);
  or (_01995_, _01994_, _01769_);
  and (_01996_, _01995_, _01993_);
  or (_01997_, _01986_, _01896_);
  or (_01998_, _01997_, _01769_);
  or (_01999_, _01958_, _01933_);
  or (_02000_, _01999_, _01769_);
  and (_02001_, _02000_, _01998_);
  and (_02002_, _02001_, _01996_);
  and (_02003_, _02002_, _01991_);
  or (_02004_, _02003_, \oc8051_golden_model_1.PC [1]);
  nand (_02005_, _02002_, _01991_);
  and (_02006_, _01651_, _01615_);
  not (_02007_, _02006_);
  or (_02008_, _02007_, _02005_);
  nand (_02009_, _02008_, _02004_);
  nand (_02010_, _02009_, _01985_);
  and (_02011_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  and (_02012_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_02013_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_02014_, _02013_, _02012_);
  and (_02015_, _02014_, _02011_);
  nor (_02016_, _02014_, _02011_);
  nor (_02017_, _02016_, _02015_);
  not (_02018_, _02017_);
  or (_02019_, _02018_, _01985_);
  not (_02020_, _01768_);
  not (_02021_, _01704_);
  and (_02022_, _02021_, _01673_);
  and (_02023_, _02022_, _02020_);
  and (_02024_, _02023_, _01959_);
  and (_02025_, _01983_, _01770_);
  nor (_02026_, _02025_, _02024_);
  and (_02027_, _02026_, _02019_);
  nand (_02028_, _02027_, _02010_);
  not (_02029_, _01959_);
  nor (_02030_, _01982_, _02029_);
  not (_02031_, _02030_);
  or (_02032_, _02026_, _01620_);
  and (_02033_, _02032_, _02031_);
  nand (_02034_, _02033_, _02028_);
  not (_02035_, _01978_);
  and (_02036_, \oc8051_golden_model_1.ACC [0], _01647_);
  and (_02037_, _02006_, \oc8051_golden_model_1.ACC [1]);
  nor (_02038_, _02006_, \oc8051_golden_model_1.ACC [1]);
  nor (_02039_, _02038_, _02037_);
  nor (_02040_, _02039_, _02036_);
  and (_02041_, _02039_, _02036_);
  nor (_02042_, _02041_, _02040_);
  and (_02043_, _02042_, _02030_);
  nor (_02044_, _02043_, _02035_);
  nand (_02045_, _02044_, _02034_);
  and (_02046_, _02045_, _01979_);
  not (_02047_, _01985_);
  nor (_02048_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_02049_, _02048_, _02011_);
  nand (_02050_, _02049_, _02047_);
  and (_02051_, _01985_, _01647_);
  nand (_02052_, _02051_, _02003_);
  nand (_02053_, _02052_, _02050_);
  nand (_02054_, _02053_, _02026_);
  and (_02055_, _02026_, _02003_);
  or (_02056_, _02055_, _01647_);
  nand (_02057_, _02056_, _02054_);
  nand (_02058_, _02057_, _02031_);
  not (_02059_, \oc8051_golden_model_1.ACC [0]);
  and (_02060_, _02059_, \oc8051_golden_model_1.PC [0]);
  or (_02061_, _02060_, _02031_);
  or (_02062_, _02061_, _02036_);
  and (_02063_, _02062_, _01978_);
  nand (_02064_, _02063_, _02058_);
  or (_02065_, _01978_, \oc8051_golden_model_1.PC [0]);
  nand (_02066_, _02065_, _02064_);
  or (_02067_, _02066_, _02046_);
  nor (_02068_, _02015_, _02012_);
  and (_02069_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_02070_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_02071_, _02070_, _02069_);
  not (_02072_, _02071_);
  nor (_02073_, _02072_, _02068_);
  and (_02074_, _02072_, _02068_);
  nor (_02075_, _02074_, _02073_);
  nand (_02076_, _02075_, _02047_);
  and (_02077_, _02076_, _02026_);
  nor (_02078_, _01615_, _01625_);
  and (_02079_, _01615_, _01625_);
  nor (_02080_, _02079_, _02078_);
  or (_02081_, _02080_, _02005_);
  nand (_02082_, _02081_, _01985_);
  nand (_02083_, _02082_, _02077_);
  and (_02084_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_02085_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_02086_, _02085_, _02084_);
  or (_02087_, _02086_, _02055_);
  and (_02088_, _02087_, _02031_);
  nand (_02089_, _02088_, _02083_);
  and (_02090_, _02086_, _01955_);
  nor (_02091_, _02041_, _02037_);
  and (_02092_, _02080_, \oc8051_golden_model_1.ACC [2]);
  nor (_02093_, _02080_, \oc8051_golden_model_1.ACC [2]);
  nor (_02094_, _02093_, _02092_);
  not (_02095_, _02094_);
  nor (_02096_, _02095_, _02091_);
  and (_02097_, _02095_, _02091_);
  nor (_02098_, _02097_, _02096_);
  and (_02099_, _02098_, _02030_);
  nor (_02100_, _02099_, _02090_);
  and (_02101_, _02100_, _01977_);
  nand (_02102_, _02101_, _02089_);
  or (_02103_, _02086_, _01978_);
  and (_02104_, _02103_, _02102_);
  and (_02105_, _02084_, \oc8051_golden_model_1.PC [3]);
  nor (_02106_, _02084_, \oc8051_golden_model_1.PC [3]);
  nor (_02107_, _02106_, _02105_);
  not (_02108_, _02107_);
  nand (_02109_, _02055_, _01978_);
  nand (_02110_, _02109_, _02108_);
  nor (_02111_, _02073_, _02069_);
  and (_02112_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_02113_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_02114_, _02113_, _02112_);
  not (_02115_, _02114_);
  nor (_02116_, _02115_, _02111_);
  and (_02117_, _02115_, _02111_);
  nor (_02118_, _02117_, _02116_);
  or (_02119_, _02118_, _01985_);
  not (_02120_, _01627_);
  nor (_02121_, _02078_, _01616_);
  nor (_02122_, _02121_, _02120_);
  and (_02123_, _01985_, _02122_);
  nand (_02124_, _02123_, _02003_);
  nand (_02125_, _02124_, _02119_);
  and (_02126_, _02031_, _02026_);
  and (_02127_, _02126_, _02125_);
  nor (_02128_, _02096_, _02092_);
  not (_02129_, \oc8051_golden_model_1.ACC [3]);
  nor (_02130_, _02122_, _02129_);
  and (_02131_, _02122_, _02129_);
  nor (_02132_, _02131_, _02130_);
  and (_02133_, _02132_, _02128_);
  nor (_02134_, _02132_, _02128_);
  nor (_02135_, _02134_, _02133_);
  and (_02136_, _02135_, _02030_);
  or (_02137_, _02136_, _02127_);
  nand (_02138_, _02137_, _01978_);
  nand (_02139_, _02138_, _02110_);
  or (_02140_, _02139_, _02104_);
  or (_02141_, _02140_, _02067_);
  or (_02142_, _02141_, _27284_);
  nand (_02143_, _02103_, _02102_);
  and (_02144_, _02138_, _02110_);
  or (_02145_, _02144_, _02143_);
  or (_02146_, _02145_, _02067_);
  or (_02147_, _02146_, _27120_);
  and (_02148_, _02147_, _02142_);
  or (_02149_, _02139_, _02143_);
  nand (_02150_, _02045_, _01979_);
  or (_02151_, _02066_, _02150_);
  or (_02152_, _02151_, _02149_);
  or (_02153_, _02152_, _27530_);
  or (_02154_, _02151_, _02145_);
  or (_02155_, _02154_, _27202_);
  and (_02156_, _02155_, _02153_);
  and (_02157_, _02156_, _02148_);
  and (_02158_, _02065_, _02064_);
  or (_02159_, _02158_, _02046_);
  or (_02160_, _02159_, _02140_);
  or (_02161_, _02160_, _27243_);
  or (_02162_, _02159_, _02145_);
  or (_02163_, _02162_, _27072_);
  and (_02164_, _02163_, _02161_);
  or (_02165_, _02144_, _02104_);
  or (_02166_, _02165_, _02159_);
  or (_02167_, _02166_, _26900_);
  or (_02168_, _02165_, _02067_);
  or (_02169_, _02168_, _26941_);
  and (_02170_, _02169_, _02167_);
  and (_02171_, _02170_, _02164_);
  and (_02172_, _02171_, _02157_);
  or (_02173_, _02159_, _02149_);
  or (_02174_, _02173_, _27407_);
  or (_02175_, _02158_, _02150_);
  or (_02176_, _02175_, _02140_);
  or (_02177_, _02176_, _27325_);
  and (_02178_, _02177_, _02174_);
  or (_02179_, _02175_, _02145_);
  or (_02180_, _02179_, _27161_);
  or (_02182_, _02165_, _02175_);
  or (_02184_, _02182_, _26982_);
  and (_02186_, _02184_, _02180_);
  and (_02188_, _02186_, _02178_);
  or (_02190_, _02149_, _02067_);
  or (_02192_, _02190_, _27448_);
  or (_02194_, _02151_, _02140_);
  or (_02195_, _02194_, _27366_);
  and (_02196_, _02195_, _02192_);
  or (_02197_, _02175_, _02149_);
  or (_02198_, _02197_, _27489_);
  or (_02199_, _02165_, _02151_);
  or (_02200_, _02199_, _27023_);
  and (_02201_, _02200_, _02198_);
  and (_02202_, _02201_, _02196_);
  and (_02203_, _02202_, _02188_);
  and (_02204_, _02203_, _02172_);
  and (_02205_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_02206_, _02205_, \oc8051_golden_model_1.PC [10]);
  and (_02207_, \oc8051_golden_model_1.PC [7], \oc8051_golden_model_1.PC [6]);
  and (_02208_, _02207_, _01901_);
  and (_02209_, _02105_, _02208_);
  and (_02210_, _02209_, _02206_);
  and (_02211_, _02210_, \oc8051_golden_model_1.PC [11]);
  and (_02212_, _02211_, \oc8051_golden_model_1.PC [12]);
  and (_02213_, _02212_, \oc8051_golden_model_1.PC [13]);
  nor (_02214_, _02213_, \oc8051_golden_model_1.PC [14]);
  and (_02215_, _02213_, \oc8051_golden_model_1.PC [14]);
  nor (_02216_, _02215_, _02214_);
  not (_02217_, _02216_);
  nor (_02218_, _02217_, _02204_);
  and (_02219_, _02217_, _02204_);
  nor (_02220_, _02219_, _02218_);
  not (_02221_, _02220_);
  not (_02222_, _02204_);
  and (_02223_, _02209_, \oc8051_golden_model_1.PC [8]);
  and (_02224_, _02223_, \oc8051_golden_model_1.PC [9]);
  and (_02225_, _02224_, \oc8051_golden_model_1.PC [10]);
  and (_02226_, _02225_, \oc8051_golden_model_1.PC [11]);
  and (_02227_, _02226_, \oc8051_golden_model_1.PC [12]);
  and (_02228_, _02227_, \oc8051_golden_model_1.PC [13]);
  nor (_02229_, _02227_, \oc8051_golden_model_1.PC [13]);
  nor (_02230_, _02229_, _02228_);
  and (_02231_, _02230_, _02222_);
  nor (_02232_, _02230_, _02222_);
  nor (_02233_, _02211_, \oc8051_golden_model_1.PC [12]);
  nor (_02234_, _02233_, _02212_);
  not (_02235_, _02234_);
  nor (_02236_, _02235_, _02204_);
  nor (_02237_, _02224_, \oc8051_golden_model_1.PC [10]);
  nor (_02238_, _02237_, _02210_);
  not (_02239_, _02238_);
  nor (_02240_, _02239_, _02204_);
  not (_02241_, _02240_);
  nor (_02242_, _02225_, \oc8051_golden_model_1.PC [11]);
  nor (_02243_, _02242_, _02226_);
  and (_02244_, _02243_, _02222_);
  nor (_02245_, _02243_, _02222_);
  nor (_02246_, _02245_, _02244_);
  and (_02247_, _02239_, _02204_);
  nor (_02248_, _02247_, _02240_);
  and (_02249_, _02248_, _02246_);
  nor (_02250_, _02223_, \oc8051_golden_model_1.PC [9]);
  nor (_02251_, _02250_, _02224_);
  not (_02252_, _02251_);
  nor (_02253_, _02252_, _02204_);
  and (_02254_, _02252_, _02204_);
  nor (_02255_, _02254_, _02253_);
  and (_02256_, _01901_, \oc8051_golden_model_1.PC [6]);
  and (_02257_, _02105_, _02256_);
  nor (_02258_, _02257_, \oc8051_golden_model_1.PC [7]);
  nor (_02259_, _02258_, _02209_);
  not (_02260_, _02259_);
  nor (_02261_, _02260_, _02204_);
  and (_02262_, _02260_, _02204_);
  nor (_02263_, _02262_, _02261_);
  not (_02264_, _02263_);
  nor (_02265_, _02152_, _27565_);
  nor (_02266_, _02194_, _27401_);
  nor (_02267_, _02266_, _02265_);
  nor (_02268_, _02179_, _27196_);
  nor (_02269_, _02168_, _26976_);
  nor (_02270_, _02269_, _02268_);
  and (_02271_, _02270_, _02267_);
  nor (_02272_, _02197_, _27524_);
  nor (_02273_, _02190_, _27483_);
  nor (_02274_, _02273_, _02272_);
  nor (_02275_, _02176_, _27360_);
  nor (_02276_, _02160_, _27278_);
  nor (_02277_, _02276_, _02275_);
  and (_02278_, _02277_, _02274_);
  and (_02279_, _02278_, _02271_);
  nor (_02280_, _02162_, _27110_);
  nor (_02281_, _02199_, _27062_);
  nor (_02282_, _02281_, _02280_);
  nor (_02283_, _02154_, _27237_);
  nor (_02284_, _02146_, _27155_);
  nor (_02285_, _02284_, _02283_);
  and (_02286_, _02285_, _02282_);
  nor (_02287_, _02173_, _27442_);
  nor (_02288_, _02141_, _27319_);
  nor (_02289_, _02288_, _02287_);
  nor (_02290_, _02166_, _26935_);
  nor (_02291_, _02182_, _27017_);
  nor (_02292_, _02291_, _02290_);
  and (_02293_, _02292_, _02289_);
  and (_02294_, _02293_, _02286_);
  and (_02295_, _02294_, _02279_);
  and (_02296_, _02105_, _01901_);
  nor (_02297_, _02296_, \oc8051_golden_model_1.PC [6]);
  nor (_02298_, _02297_, _02257_);
  not (_02299_, _02298_);
  nor (_02300_, _02299_, _02295_);
  and (_02301_, _02299_, _02295_);
  nor (_02302_, _02301_, _02300_);
  nor (_02303_, _02190_, _27478_);
  nor (_02304_, _02154_, _27232_);
  nor (_02305_, _02304_, _02303_);
  nor (_02306_, _02146_, _27150_);
  nor (_02307_, _02168_, _26971_);
  nor (_02308_, _02307_, _02306_);
  and (_02309_, _02308_, _02305_);
  nor (_02310_, _02141_, _27314_);
  nor (_02311_, _02176_, _27355_);
  nor (_02312_, _02311_, _02310_);
  nor (_02313_, _02194_, _27396_);
  nor (_02314_, _02199_, _27054_);
  nor (_02315_, _02314_, _02313_);
  and (_02316_, _02315_, _02312_);
  and (_02317_, _02316_, _02309_);
  nor (_02318_, _02179_, _27191_);
  nor (_02319_, _02162_, _27102_);
  nor (_02320_, _02319_, _02318_);
  nor (_02321_, _02197_, _27519_);
  nor (_02322_, _02166_, _26930_);
  nor (_02323_, _02322_, _02321_);
  and (_02324_, _02323_, _02320_);
  nor (_02325_, _02152_, _27560_);
  nor (_02326_, _02182_, _27012_);
  nor (_02327_, _02326_, _02325_);
  nor (_02328_, _02173_, _27437_);
  nor (_02329_, _02160_, _27273_);
  nor (_02330_, _02329_, _02328_);
  and (_02331_, _02330_, _02327_);
  and (_02332_, _02331_, _02324_);
  and (_02333_, _02332_, _02317_);
  and (_02334_, _02105_, \oc8051_golden_model_1.PC [4]);
  nor (_02335_, _02334_, \oc8051_golden_model_1.PC [5]);
  nor (_02336_, _02335_, _02296_);
  not (_02337_, _02336_);
  nor (_02338_, _02337_, _02333_);
  and (_02339_, _02337_, _02333_);
  nor (_02340_, _02154_, _27227_);
  nor (_02341_, _02199_, _27048_);
  nor (_02342_, _02341_, _02340_);
  nor (_02343_, _02197_, _27514_);
  nor (_02344_, _02160_, _27268_);
  nor (_02345_, _02344_, _02343_);
  and (_02346_, _02345_, _02342_);
  nor (_02347_, _02182_, _27007_);
  nor (_02348_, _02168_, _26966_);
  nor (_02349_, _02348_, _02347_);
  nor (_02350_, _02146_, _27145_);
  nor (_02351_, _02162_, _27097_);
  nor (_02352_, _02351_, _02350_);
  and (_02353_, _02352_, _02349_);
  and (_02354_, _02353_, _02346_);
  nor (_02355_, _02190_, _27473_);
  nor (_02356_, _02194_, _27391_);
  nor (_02357_, _02356_, _02355_);
  nor (_02358_, _02152_, _27555_);
  nor (_02359_, _02173_, _27432_);
  nor (_02360_, _02359_, _02358_);
  and (_02361_, _02360_, _02357_);
  nor (_02362_, _02176_, _27350_);
  nor (_02363_, _02141_, _27309_);
  nor (_02364_, _02363_, _02362_);
  nor (_02365_, _02179_, _27186_);
  nor (_02366_, _02166_, _26925_);
  nor (_02367_, _02366_, _02365_);
  and (_02368_, _02367_, _02364_);
  and (_02369_, _02368_, _02361_);
  and (_02370_, _02369_, _02354_);
  nor (_02371_, _02105_, \oc8051_golden_model_1.PC [4]);
  nor (_02372_, _02371_, _02334_);
  not (_02373_, _02372_);
  nor (_02374_, _02373_, _02370_);
  or (_02375_, _02152_, _27550_);
  or (_02376_, _02168_, _26961_);
  and (_02377_, _02376_, _02375_);
  or (_02378_, _02194_, _27386_);
  or (_02379_, _02166_, _26920_);
  and (_02380_, _02379_, _02378_);
  and (_02381_, _02380_, _02377_);
  or (_02382_, _02141_, _27304_);
  or (_02383_, _02182_, _27002_);
  and (_02384_, _02383_, _02382_);
  or (_02385_, _02154_, _27222_);
  or (_02386_, _02146_, _27140_);
  and (_02387_, _02386_, _02385_);
  and (_02388_, _02387_, _02384_);
  and (_02389_, _02388_, _02381_);
  or (_02390_, _02199_, _27043_);
  or (_02391_, _02162_, _27092_);
  and (_02392_, _02391_, _02390_);
  or (_02393_, _02197_, _27509_);
  or (_02394_, _02176_, _27345_);
  and (_02395_, _02394_, _02393_);
  and (_02396_, _02395_, _02392_);
  or (_02397_, _02190_, _27468_);
  or (_02398_, _02160_, _27263_);
  and (_02399_, _02398_, _02397_);
  or (_02400_, _02173_, _27427_);
  or (_02401_, _02179_, _27181_);
  and (_02402_, _02401_, _02400_);
  and (_02403_, _02402_, _02399_);
  and (_02404_, _02403_, _02396_);
  nand (_02405_, _02404_, _02389_);
  and (_02406_, _02405_, _02107_);
  nor (_02407_, _02405_, _02107_);
  not (_02408_, _02086_);
  nor (_02409_, _02154_, _27217_);
  nor (_02410_, _02168_, _26956_);
  nor (_02411_, _02410_, _02409_);
  nor (_02412_, _02160_, _27258_);
  nor (_02413_, _02182_, _26997_);
  nor (_02414_, _02413_, _02412_);
  and (_02415_, _02414_, _02411_);
  nor (_02416_, _02190_, _27463_);
  nor (_02417_, _02173_, _27422_);
  nor (_02418_, _02417_, _02416_);
  nor (_02419_, _02146_, _27135_);
  nor (_02420_, _02162_, _27087_);
  nor (_02421_, _02420_, _02419_);
  and (_02422_, _02421_, _02418_);
  and (_02423_, _02422_, _02415_);
  nor (_02424_, _02197_, _27504_);
  nor (_02425_, _02194_, _27381_);
  nor (_02426_, _02425_, _02424_);
  nor (_02427_, _02199_, _27038_);
  nor (_02428_, _02166_, _26915_);
  nor (_02429_, _02428_, _02427_);
  and (_02430_, _02429_, _02426_);
  nor (_02431_, _02176_, _27340_);
  nor (_02432_, _02141_, _27299_);
  nor (_02433_, _02432_, _02431_);
  nor (_02434_, _02152_, _27545_);
  nor (_02435_, _02179_, _27176_);
  nor (_02436_, _02435_, _02434_);
  and (_02437_, _02436_, _02433_);
  and (_02438_, _02437_, _02430_);
  and (_02439_, _02438_, _02423_);
  nor (_02440_, _02439_, _02408_);
  nor (_02441_, _02154_, _27212_);
  nor (_02442_, _02166_, _26910_);
  nor (_02443_, _02442_, _02441_);
  nor (_02444_, _02160_, _27253_);
  nor (_02445_, _02182_, _26992_);
  nor (_02446_, _02445_, _02444_);
  and (_02447_, _02446_, _02443_);
  nor (_02448_, _02179_, _27171_);
  nor (_02449_, _02146_, _27130_);
  nor (_02450_, _02449_, _02448_);
  nor (_02451_, _02190_, _27458_);
  nor (_02452_, _02173_, _27417_);
  nor (_02453_, _02452_, _02451_);
  and (_02454_, _02453_, _02450_);
  and (_02455_, _02454_, _02447_);
  nor (_02456_, _02197_, _27499_);
  nor (_02457_, _02194_, _27376_);
  nor (_02458_, _02457_, _02456_);
  nor (_02459_, _02199_, _27033_);
  nor (_02460_, _02168_, _26951_);
  nor (_02461_, _02460_, _02459_);
  and (_02462_, _02461_, _02458_);
  nor (_02463_, _02176_, _27335_);
  nor (_02464_, _02141_, _27294_);
  nor (_02465_, _02464_, _02463_);
  nor (_02466_, _02152_, _27540_);
  nor (_02467_, _02162_, _27082_);
  nor (_02468_, _02467_, _02466_);
  and (_02469_, _02468_, _02465_);
  and (_02470_, _02469_, _02462_);
  and (_02471_, _02470_, _02455_);
  nor (_02472_, _02471_, \oc8051_golden_model_1.PC [1]);
  or (_02473_, _02179_, _27166_);
  or (_02474_, _02146_, _27125_);
  and (_02475_, _02474_, _02473_);
  or (_02476_, _02199_, _27028_);
  or (_02477_, _02182_, _26987_);
  and (_02478_, _02477_, _02476_);
  and (_02479_, _02478_, _02475_);
  or (_02480_, _02173_, _27412_);
  or (_02481_, _02141_, _27289_);
  and (_02482_, _02481_, _02480_);
  or (_02483_, _02194_, _27371_);
  or (_02484_, _02160_, _27248_);
  and (_02485_, _02484_, _02483_);
  and (_02486_, _02485_, _02482_);
  and (_02487_, _02486_, _02479_);
  or (_02488_, _02166_, _26905_);
  or (_02489_, _02168_, _26946_);
  and (_02490_, _02489_, _02488_);
  or (_02491_, _02154_, _27207_);
  or (_02492_, _02162_, _27077_);
  and (_02493_, _02492_, _02491_);
  and (_02494_, _02493_, _02490_);
  or (_02495_, _02152_, _27535_);
  or (_02496_, _02197_, _27494_);
  and (_02497_, _02496_, _02495_);
  or (_02498_, _02190_, _27453_);
  or (_02499_, _02176_, _27330_);
  and (_02500_, _02499_, _02498_);
  and (_02501_, _02500_, _02497_);
  and (_02502_, _02501_, _02494_);
  and (_02503_, _02502_, _02487_);
  nor (_02504_, _02503_, _01647_);
  and (_02505_, _02471_, \oc8051_golden_model_1.PC [1]);
  nor (_02506_, _02505_, _02472_);
  and (_02507_, _02506_, _02504_);
  nor (_02508_, _02507_, _02472_);
  and (_02509_, _02439_, _02408_);
  nor (_02510_, _02509_, _02440_);
  not (_02511_, _02510_);
  nor (_02512_, _02511_, _02508_);
  nor (_02513_, _02512_, _02440_);
  nor (_02514_, _02513_, _02407_);
  nor (_02515_, _02514_, _02406_);
  and (_02516_, _02373_, _02370_);
  nor (_02517_, _02516_, _02374_);
  not (_02518_, _02517_);
  nor (_02519_, _02518_, _02515_);
  nor (_02520_, _02519_, _02374_);
  nor (_02521_, _02520_, _02339_);
  or (_02522_, _02521_, _02338_);
  and (_02523_, _02522_, _02302_);
  nor (_02524_, _02523_, _02300_);
  nor (_02525_, _02524_, _02264_);
  nor (_02526_, _02525_, _02261_);
  nor (_02527_, _02209_, \oc8051_golden_model_1.PC [8]);
  nor (_02528_, _02527_, _02223_);
  not (_02529_, _02528_);
  nor (_02530_, _02529_, _02204_);
  and (_02531_, _02529_, _02204_);
  nor (_02532_, _02531_, _02530_);
  not (_02533_, _02532_);
  nor (_02534_, _02533_, _02526_);
  and (_02535_, _02534_, _02255_);
  and (_02536_, _02535_, _02249_);
  nor (_02537_, _02530_, _02253_);
  not (_02538_, _02537_);
  and (_02539_, _02538_, _02249_);
  or (_02540_, _02539_, _02244_);
  nor (_02541_, _02540_, _02536_);
  and (_02542_, _02541_, _02241_);
  and (_02543_, _02235_, _02204_);
  nor (_02544_, _02543_, _02236_);
  not (_02545_, _02544_);
  nor (_02546_, _02545_, _02542_);
  nor (_02547_, _02546_, _02236_);
  nor (_02548_, _02547_, _02232_);
  nor (_02549_, _02548_, _02231_);
  nor (_02550_, _02549_, _02221_);
  nor (_02551_, _02550_, _02218_);
  nor (_02552_, _02215_, \oc8051_golden_model_1.PC [15]);
  and (_02553_, _02228_, \oc8051_golden_model_1.PC [14]);
  and (_02554_, _02553_, \oc8051_golden_model_1.PC [15]);
  nor (_02555_, _02554_, _02552_);
  not (_02556_, _02555_);
  and (_02557_, _02556_, _02204_);
  nor (_02558_, _02556_, _02204_);
  nor (_02559_, _02558_, _02557_);
  nor (_02560_, _02559_, _02551_);
  and (_02561_, _02559_, _02551_);
  or (_02562_, _02561_, _02560_);
  or (_02563_, _02562_, _01953_);
  not (_02564_, _01705_);
  and (_02565_, _01980_, _01736_);
  and (_02566_, _02565_, _02564_);
  and (_02567_, _02566_, _01966_);
  not (_02568_, _01953_);
  or (_02569_, _02555_, _02568_);
  and (_02570_, _02569_, _02567_);
  and (_02571_, _02570_, _02563_);
  not (_02572_, _01982_);
  and (_02573_, _02572_, _01966_);
  not (_02574_, _02573_);
  and (_02575_, _02023_, _01966_);
  not (_02576_, _01966_);
  nor (_02577_, _02576_, _01925_);
  nand (_02578_, _02577_, _02556_);
  and (_02579_, _01651_, \oc8051_golden_model_1.PC [2]);
  and (_02580_, _02579_, \oc8051_golden_model_1.PC [3]);
  and (_02581_, _02580_, _02208_);
  and (_02582_, _02581_, _02206_);
  and (_02583_, _02582_, \oc8051_golden_model_1.PC [11]);
  and (_02584_, _02583_, \oc8051_golden_model_1.PC [12]);
  and (_02585_, _02584_, \oc8051_golden_model_1.PC [13]);
  and (_02586_, _02585_, \oc8051_golden_model_1.PC [14]);
  nor (_02587_, _02586_, \oc8051_golden_model_1.PC [15]);
  and (_02588_, _02581_, \oc8051_golden_model_1.PC [8]);
  and (_02589_, _02588_, \oc8051_golden_model_1.PC [9]);
  and (_02590_, _02589_, \oc8051_golden_model_1.PC [10]);
  and (_02591_, _02590_, \oc8051_golden_model_1.PC [11]);
  and (_02592_, _02591_, \oc8051_golden_model_1.PC [12]);
  and (_02593_, _02592_, \oc8051_golden_model_1.PC [13]);
  and (_02594_, _02593_, \oc8051_golden_model_1.PC [14]);
  and (_02595_, _02594_, \oc8051_golden_model_1.PC [15]);
  nor (_02596_, _02595_, _02587_);
  and (_02597_, _02596_, _02024_);
  nor (_02598_, _01999_, _01982_);
  not (_02599_, _02598_);
  nor (_02600_, _02439_, \oc8051_golden_model_1.ACC [2]);
  and (_02601_, _02439_, \oc8051_golden_model_1.ACC [2]);
  nor (_02602_, _02601_, _02600_);
  and (_02603_, _02405_, _02129_);
  nor (_02604_, _02405_, _02129_);
  nor (_02605_, _02604_, _02603_);
  and (_02606_, _02605_, _02602_);
  nor (_02607_, _02471_, \oc8051_golden_model_1.ACC [1]);
  and (_02608_, _02471_, \oc8051_golden_model_1.ACC [1]);
  nor (_02609_, _02608_, _02607_);
  nor (_02610_, _02503_, \oc8051_golden_model_1.ACC [0]);
  and (_02611_, _02503_, \oc8051_golden_model_1.ACC [0]);
  nor (_02612_, _02611_, _02610_);
  and (_02613_, _02612_, _02609_);
  and (_02614_, _02613_, _02606_);
  nor (_02615_, _02204_, \oc8051_golden_model_1.ACC [7]);
  and (_02616_, _02204_, \oc8051_golden_model_1.ACC [7]);
  nor (_02617_, _02616_, _02615_);
  nor (_02618_, _02295_, \oc8051_golden_model_1.ACC [6]);
  and (_02619_, _02295_, \oc8051_golden_model_1.ACC [6]);
  nor (_02620_, _02619_, _02618_);
  and (_02621_, _02620_, _02617_);
  nor (_02622_, _02370_, \oc8051_golden_model_1.ACC [4]);
  and (_02623_, _02370_, \oc8051_golden_model_1.ACC [4]);
  nor (_02624_, _02623_, _02622_);
  nor (_02625_, _02333_, \oc8051_golden_model_1.ACC [5]);
  and (_02626_, _02333_, \oc8051_golden_model_1.ACC [5]);
  nor (_02627_, _02626_, _02625_);
  and (_02628_, _02627_, _02624_);
  and (_02629_, _02628_, _02621_);
  and (_02630_, _02629_, _02614_);
  and (_02631_, _01767_, _01736_);
  and (_02632_, _01917_, _02631_);
  and (_02633_, _01917_, _02020_);
  nor (_02634_, _02633_, _02632_);
  not (_02635_, _01981_);
  and (_02636_, _02635_, _01917_);
  and (_02637_, _01920_, _02631_);
  nor (_02638_, _02637_, _02636_);
  nor (_02639_, _01926_, _01981_);
  and (_02640_, _02565_, _01917_);
  nor (_02641_, _02640_, _02639_);
  and (_02642_, _02641_, _02638_);
  and (_02643_, _02642_, _02634_);
  or (_02644_, _02643_, _01999_);
  and (_02645_, _02631_, _02564_);
  and (_02646_, _02645_, _01970_);
  and (_02647_, _02566_, _01898_);
  nor (_02648_, _02647_, _02646_);
  and (_02649_, _02645_, _01954_);
  and (_02650_, _02566_, _01970_);
  nor (_02651_, _02650_, _02649_);
  and (_02652_, _02651_, _02648_);
  and (_02653_, _02566_, _01935_);
  and (_02654_, _02572_, _01942_);
  nor (_02655_, _02654_, _02653_);
  and (_02656_, _02572_, _01973_);
  nor (_02657_, _02656_, _02575_);
  and (_02658_, _02657_, _02655_);
  and (_02659_, _02658_, _02652_);
  not (_02660_, _01994_);
  and (_02661_, _02023_, _02660_);
  not (_02662_, _02661_);
  not (_02663_, _01999_);
  and (_02664_, _02023_, _02663_);
  and (_02665_, _01920_, _01980_);
  and (_02666_, _02663_, _02665_);
  nor (_02667_, _02666_, _02664_);
  and (_02668_, _02667_, _02662_);
  and (_02669_, _02572_, _01964_);
  and (_02670_, _02566_, _01983_);
  nor (_02671_, _02670_, _02669_);
  and (_02672_, _02022_, _02565_);
  and (_02673_, _02672_, _02663_);
  and (_02674_, _01924_, _02021_);
  and (_02675_, _02663_, _02674_);
  nor (_02676_, _02675_, _02673_);
  and (_02677_, _02676_, _02671_);
  and (_02678_, _02677_, _02668_);
  and (_02679_, _02678_, _02659_);
  and (_02680_, _02679_, _02644_);
  nor (_02681_, _02680_, _02086_);
  not (_02682_, _02080_);
  and (_02683_, _02680_, _02682_);
  nor (_02684_, _02683_, _02681_);
  nor (_02685_, _02680_, _02108_);
  not (_02686_, _02122_);
  and (_02687_, _02680_, _02686_);
  nor (_02688_, _02687_, _02685_);
  not (_02689_, _02688_);
  and (_02690_, _02689_, _02684_);
  nor (_02691_, _02680_, _01647_);
  and (_02692_, _02680_, _01647_);
  nor (_02693_, _02692_, _02691_);
  nor (_02694_, _02680_, \oc8051_golden_model_1.PC [1]);
  and (_02695_, _02680_, _02006_);
  nor (_02696_, _02695_, _02694_);
  nor (_02697_, _02696_, _02693_);
  and (_02698_, _02697_, _02690_);
  and (_02699_, _02698_, _00353_);
  nor (_02700_, _02688_, _02684_);
  and (_02701_, _02700_, _02697_);
  and (_02702_, _02701_, _00388_);
  nor (_02703_, _02702_, _02699_);
  not (_02704_, _02693_);
  and (_02705_, _02696_, _02704_);
  and (_02706_, _02688_, _02684_);
  and (_02707_, _02706_, _02705_);
  and (_02708_, _02707_, _00428_);
  and (_02709_, _02693_, \oc8051_golden_model_1.PC [1]);
  and (_02710_, _02706_, _02709_);
  and (_02711_, _02710_, _00439_);
  nor (_02712_, _02711_, _02708_);
  and (_02713_, _02712_, _02703_);
  and (_02714_, _02693_, _01620_);
  and (_02715_, _02700_, _02714_);
  and (_02716_, _02715_, _00400_);
  and (_02717_, _02700_, _02705_);
  and (_02718_, _02717_, _00412_);
  nor (_02719_, _02718_, _02716_);
  and (_02720_, _02714_, _02690_);
  and (_02721_, _02720_, _00383_);
  and (_02722_, _02709_, _02690_);
  and (_02723_, _02722_, _00391_);
  nor (_02724_, _02723_, _02721_);
  and (_02725_, _02724_, _02719_);
  and (_02726_, _02725_, _02713_);
  and (_02727_, _02706_, _02697_);
  and (_02728_, _02727_, _00421_);
  and (_02729_, _02706_, _02714_);
  and (_02730_, _02729_, _00431_);
  nor (_02731_, _02730_, _02728_);
  nor (_02732_, _02689_, _02684_);
  and (_02733_, _02732_, _02709_);
  and (_02734_, _02733_, _00444_);
  and (_02735_, _02732_, _02714_);
  and (_02736_, _02735_, _00447_);
  nor (_02737_, _02736_, _02734_);
  and (_02738_, _02737_, _02731_);
  and (_02739_, _02705_, _02690_);
  and (_02740_, _02739_, _00373_);
  and (_02741_, _02709_, _02700_);
  and (_02742_, _02741_, _00417_);
  nor (_02743_, _02742_, _02740_);
  and (_02744_, _02732_, _02697_);
  and (_02745_, _02744_, _00435_);
  and (_02746_, _02732_, _02705_);
  and (_02747_, _02746_, _00453_);
  nor (_02748_, _02747_, _02745_);
  and (_02750_, _02748_, _02743_);
  and (_02751_, _02750_, _02738_);
  and (_02752_, _02751_, _02726_);
  nor (_02754_, _02585_, \oc8051_golden_model_1.PC [14]);
  nor (_02755_, _02754_, _02586_);
  not (_02756_, _02755_);
  nor (_02757_, _02756_, _02752_);
  and (_02758_, _02756_, _02752_);
  nor (_02759_, _02758_, _02757_);
  not (_02760_, _02759_);
  not (_02761_, \oc8051_golden_model_1.PC [13]);
  and (_02762_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_02763_, _02762_, _02205_);
  and (_02764_, _02581_, _02763_);
  and (_02765_, _02764_, \oc8051_golden_model_1.PC [12]);
  nor (_02766_, _02765_, _02761_);
  and (_02767_, _02765_, _02761_);
  or (_02768_, _02767_, _02766_);
  not (_02769_, _02768_);
  nor (_02770_, _02769_, _02752_);
  and (_02771_, _02769_, _02752_);
  nor (_02772_, _02583_, \oc8051_golden_model_1.PC [12]);
  nor (_02773_, _02772_, _02584_);
  not (_02774_, _02773_);
  nor (_02775_, _02774_, _02752_);
  nor (_02776_, _02589_, \oc8051_golden_model_1.PC [10]);
  nor (_02777_, _02776_, _02582_);
  not (_02778_, _02777_);
  nor (_02779_, _02778_, _02752_);
  not (_02780_, _02779_);
  not (_02781_, \oc8051_golden_model_1.PC [11]);
  nor (_02782_, _02582_, _02781_);
  and (_02783_, _02582_, _02781_);
  or (_02784_, _02783_, _02782_);
  not (_02785_, _02784_);
  nor (_02786_, _02785_, _02752_);
  and (_02787_, _02785_, _02752_);
  nor (_02788_, _02787_, _02786_);
  and (_02789_, _02778_, _02752_);
  nor (_02790_, _02789_, _02779_);
  and (_02791_, _02790_, _02788_);
  nor (_02792_, _02588_, \oc8051_golden_model_1.PC [9]);
  nor (_02793_, _02792_, _02589_);
  not (_02794_, _02793_);
  nor (_02795_, _02794_, _02752_);
  and (_02796_, _02794_, _02752_);
  nor (_02797_, _02796_, _02795_);
  and (_02798_, _02580_, _02256_);
  nor (_02799_, _02798_, \oc8051_golden_model_1.PC [7]);
  nor (_02800_, _02799_, _02581_);
  not (_02801_, _02800_);
  nor (_02802_, _02801_, _02752_);
  and (_02803_, _02801_, _02752_);
  and (_02804_, _02701_, _00918_);
  and (_02805_, _02727_, _00911_);
  nor (_02806_, _02805_, _02804_);
  and (_02807_, _02729_, _00945_);
  and (_02808_, _02733_, _00930_);
  nor (_02809_, _02808_, _02807_);
  and (_02810_, _02809_, _02806_);
  and (_02811_, _02698_, _00902_);
  and (_02812_, _02744_, _00938_);
  nor (_02813_, _02812_, _02811_);
  and (_02814_, _02720_, _00923_);
  and (_02815_, _02741_, _00913_);
  nor (_02816_, _02815_, _02814_);
  and (_02817_, _02816_, _02813_);
  and (_02818_, _02817_, _02810_);
  and (_02819_, _02707_, _00943_);
  and (_02820_, _02710_, _00940_);
  nor (_02821_, _02820_, _02819_);
  and (_02822_, _02715_, _00904_);
  and (_02823_, _02746_, _00932_);
  nor (_02824_, _02823_, _02822_);
  and (_02825_, _02824_, _02821_);
  and (_02826_, _02722_, _00920_);
  and (_02827_, _02735_, _00934_);
  nor (_02828_, _02827_, _02826_);
  and (_02829_, _02739_, _00925_);
  and (_02830_, _02717_, _00907_);
  nor (_02831_, _02830_, _02829_);
  and (_02832_, _02831_, _02828_);
  and (_02833_, _02832_, _02825_);
  and (_02834_, _02833_, _02818_);
  and (_02835_, _02580_, _01901_);
  nor (_02836_, _02835_, \oc8051_golden_model_1.PC [6]);
  nor (_02837_, _02836_, _02798_);
  not (_02838_, _02837_);
  nor (_02839_, _02838_, _02834_);
  and (_02840_, _02838_, _02834_);
  nor (_02841_, _02840_, _02839_);
  not (_02842_, _02841_);
  and (_02843_, _02701_, _00862_);
  and (_02844_, _02727_, _00858_);
  nor (_02845_, _02844_, _02843_);
  and (_02846_, _02729_, _00886_);
  and (_02847_, _02733_, _00892_);
  nor (_02848_, _02847_, _02846_);
  and (_02849_, _02848_, _02845_);
  and (_02850_, _02698_, _00849_);
  and (_02851_, _02744_, _00883_);
  nor (_02852_, _02851_, _02850_);
  and (_02853_, _02720_, _00872_);
  and (_02854_, _02717_, _00853_);
  nor (_02855_, _02854_, _02853_);
  and (_02856_, _02855_, _02852_);
  and (_02857_, _02856_, _02849_);
  and (_02858_, _02707_, _00888_);
  and (_02859_, _02710_, _00881_);
  nor (_02860_, _02859_, _02858_);
  and (_02861_, _02739_, _00876_);
  and (_02862_, _02746_, _00894_);
  nor (_02863_, _02862_, _02861_);
  and (_02864_, _02863_, _02860_);
  and (_02865_, _02715_, _00851_);
  and (_02866_, _02735_, _00896_);
  nor (_02867_, _02866_, _02865_);
  and (_02868_, _02722_, _00866_);
  and (_02869_, _02741_, _00856_);
  nor (_02870_, _02869_, _02868_);
  and (_02871_, _02870_, _02867_);
  and (_02872_, _02871_, _02864_);
  and (_02873_, _02872_, _02857_);
  and (_02874_, _02580_, \oc8051_golden_model_1.PC [4]);
  nor (_02875_, _02874_, \oc8051_golden_model_1.PC [5]);
  nor (_02876_, _02875_, _02835_);
  not (_02877_, _02876_);
  nor (_02878_, _02877_, _02873_);
  and (_02879_, _02877_, _02873_);
  and (_02880_, _02701_, _00798_);
  and (_02881_, _02746_, _00841_);
  nor (_02882_, _02881_, _02880_);
  and (_02883_, _02698_, _00794_);
  and (_02884_, _02710_, _00828_);
  nor (_02885_, _02884_, _02883_);
  and (_02886_, _02885_, _02882_);
  and (_02887_, _02715_, _00807_);
  and (_02888_, _02717_, _00809_);
  nor (_02889_, _02888_, _02887_);
  and (_02890_, _02720_, _00803_);
  and (_02891_, _02735_, _00843_);
  nor (_02892_, _02891_, _02890_);
  and (_02893_, _02892_, _02889_);
  and (_02894_, _02893_, _02886_);
  and (_02895_, _02727_, _00814_);
  and (_02896_, _02729_, _00832_);
  nor (_02897_, _02896_, _02895_);
  and (_02898_, _02707_, _00835_);
  and (_02899_, _02733_, _00839_);
  nor (_02900_, _02899_, _02898_);
  and (_02901_, _02900_, _02897_);
  and (_02902_, _02741_, _00818_);
  and (_02903_, _02744_, _00826_);
  nor (_02904_, _02903_, _02902_);
  and (_02905_, _02739_, _00801_);
  and (_02906_, _02722_, _00796_);
  nor (_02907_, _02906_, _02905_);
  and (_02908_, _02907_, _02904_);
  and (_02909_, _02908_, _02901_);
  and (_02910_, _02909_, _02894_);
  nor (_02911_, _02580_, \oc8051_golden_model_1.PC [4]);
  nor (_02912_, _02911_, _02874_);
  not (_02913_, _02912_);
  nor (_02914_, _02913_, _02910_);
  and (_02915_, _02727_, _00746_);
  and (_02916_, _02733_, _00784_);
  nor (_02917_, _02916_, _02915_);
  and (_02918_, _02741_, _00748_);
  and (_02919_, _02744_, _00773_);
  nor (_02920_, _02919_, _02918_);
  and (_02921_, _02920_, _02917_);
  and (_02922_, _02739_, _00760_);
  and (_02923_, _02722_, _00752_);
  nor (_02924_, _02923_, _02922_);
  and (_02925_, _02707_, _00778_);
  and (_02926_, _02710_, _00770_);
  nor (_02927_, _02926_, _02925_);
  and (_02928_, _02927_, _02924_);
  and (_02929_, _02928_, _02921_);
  and (_02930_, _02735_, _00788_);
  and (_02931_, _02746_, _00786_);
  nor (_02932_, _02931_, _02930_);
  and (_02933_, _02720_, _00757_);
  and (_02934_, _02701_, _00754_);
  nor (_02935_, _02934_, _02933_);
  and (_02936_, _02935_, _02932_);
  and (_02937_, _02715_, _00741_);
  and (_02938_, _02717_, _00743_);
  nor (_02939_, _02938_, _02937_);
  and (_02940_, _02698_, _00739_);
  and (_02941_, _02729_, _00776_);
  nor (_02942_, _02941_, _02940_);
  and (_02943_, _02942_, _02939_);
  and (_02944_, _02943_, _02936_);
  and (_02945_, _02944_, _02929_);
  nor (_02946_, _02579_, \oc8051_golden_model_1.PC [3]);
  nor (_02947_, _02946_, _02580_);
  not (_02948_, _02947_);
  nor (_02949_, _02948_, _02945_);
  and (_02950_, _02948_, _02945_);
  and (_02951_, _02698_, _00684_);
  and (_02952_, _02733_, _00728_);
  nor (_02953_, _02952_, _02951_);
  and (_02954_, _02701_, _00688_);
  and (_02955_, _02746_, _00731_);
  nor (_02956_, _02955_, _02954_);
  and (_02957_, _02956_, _02953_);
  and (_02958_, _02717_, _00699_);
  and (_02959_, _02735_, _00733_);
  nor (_02960_, _02959_, _02958_);
  and (_02961_, _02727_, _00704_);
  and (_02962_, _02707_, _00723_);
  nor (_02963_, _02962_, _02961_);
  and (_02964_, _02963_, _02960_);
  and (_02965_, _02964_, _02957_);
  and (_02966_, _02744_, _00716_);
  and (_02967_, _02710_, _00712_);
  nor (_02968_, _02967_, _02966_);
  and (_02969_, _02720_, _00691_);
  and (_02970_, _02715_, _00697_);
  nor (_02971_, _02970_, _02969_);
  and (_02972_, _02971_, _02968_);
  and (_02973_, _02739_, _00693_);
  and (_02974_, _02741_, _00702_);
  nor (_02975_, _02974_, _02973_);
  and (_02976_, _02722_, _00686_);
  and (_02977_, _02729_, _00721_);
  nor (_02978_, _02977_, _02976_);
  and (_02979_, _02978_, _02975_);
  and (_02980_, _02979_, _02972_);
  and (_02981_, _02980_, _02965_);
  nor (_02982_, _01651_, \oc8051_golden_model_1.PC [2]);
  nor (_02983_, _02982_, _02579_);
  not (_02984_, _02983_);
  nor (_02985_, _02984_, _02981_);
  and (_02986_, _02727_, _00649_);
  and (_02987_, _02746_, _00674_);
  nor (_02988_, _02987_, _02986_);
  and (_02989_, _02717_, _00644_);
  and (_02990_, _02735_, _00677_);
  nor (_02991_, _02990_, _02989_);
  and (_02992_, _02991_, _02988_);
  and (_02993_, _02701_, _00631_);
  and (_02994_, _02733_, _00672_);
  nor (_02995_, _02994_, _02993_);
  and (_02996_, _02739_, _00636_);
  and (_02997_, _02722_, _00633_);
  nor (_02998_, _02997_, _02996_);
  and (_02999_, _02998_, _02995_);
  and (_03000_, _02999_, _02992_);
  and (_03001_, _02720_, _00638_);
  and (_03002_, _02744_, _00658_);
  nor (_03003_, _03002_, _03001_);
  and (_03004_, _02741_, _00647_);
  and (_03005_, _02729_, _00664_);
  nor (_03006_, _03005_, _03004_);
  and (_03007_, _03006_, _03003_);
  and (_03008_, _02715_, _00642_);
  and (_03009_, _02710_, _00654_);
  nor (_03010_, _03009_, _03008_);
  and (_03011_, _02698_, _00629_);
  and (_03012_, _02707_, _00668_);
  nor (_03013_, _03012_, _03011_);
  and (_03014_, _03013_, _03010_);
  and (_03015_, _03014_, _03007_);
  and (_03016_, _03015_, _03000_);
  nor (_03017_, _03016_, _02006_);
  and (_03018_, _02698_, _00574_);
  and (_03019_, _02701_, _00576_);
  nor (_03020_, _03019_, _03018_);
  and (_03021_, _02727_, _00594_);
  and (_03022_, _02746_, _00619_);
  nor (_03023_, _03022_, _03021_);
  and (_03024_, _03023_, _03020_);
  and (_03025_, _02715_, _00587_);
  and (_03026_, _02717_, _00589_);
  nor (_03027_, _03026_, _03025_);
  and (_03028_, _02739_, _00581_);
  and (_03029_, _02722_, _00578_);
  nor (_03030_, _03029_, _03028_);
  and (_03031_, _03030_, _03027_);
  and (_03032_, _03031_, _03024_);
  and (_03033_, _02707_, _00610_);
  and (_03034_, _02744_, _00601_);
  nor (_03035_, _03034_, _03033_);
  and (_03036_, _02729_, _00606_);
  and (_03037_, _02710_, _00599_);
  nor (_03038_, _03037_, _03036_);
  and (_03039_, _03038_, _03035_);
  and (_03040_, _02720_, _00583_);
  and (_03041_, _02741_, _00592_);
  nor (_03042_, _03041_, _03040_);
  and (_03043_, _02733_, _00617_);
  and (_03044_, _02735_, _00621_);
  nor (_03045_, _03044_, _03043_);
  and (_03046_, _03045_, _03042_);
  and (_03047_, _03046_, _03039_);
  and (_03048_, _03047_, _03032_);
  nor (_03049_, _03048_, \oc8051_golden_model_1.PC [0]);
  and (_03050_, _03016_, _02006_);
  nor (_03051_, _03050_, _03017_);
  and (_03052_, _03051_, _03049_);
  nor (_03053_, _03052_, _03017_);
  and (_03054_, _02984_, _02981_);
  nor (_03055_, _03054_, _02985_);
  not (_03056_, _03055_);
  nor (_03057_, _03056_, _03053_);
  nor (_03058_, _03057_, _02985_);
  nor (_03059_, _03058_, _02950_);
  nor (_03060_, _03059_, _02949_);
  and (_03061_, _02913_, _02910_);
  nor (_03062_, _03061_, _02914_);
  not (_03063_, _03062_);
  nor (_03064_, _03063_, _03060_);
  nor (_03065_, _03064_, _02914_);
  nor (_03066_, _03065_, _02879_);
  nor (_03067_, _03066_, _02878_);
  nor (_03068_, _03067_, _02842_);
  nor (_03069_, _03068_, _02839_);
  nor (_03070_, _03069_, _02803_);
  or (_03071_, _03070_, _02802_);
  nor (_03072_, _02581_, \oc8051_golden_model_1.PC [8]);
  nor (_03073_, _03072_, _02588_);
  not (_03074_, _03073_);
  nor (_03075_, _03074_, _02752_);
  and (_03076_, _03074_, _02752_);
  nor (_03077_, _03076_, _03075_);
  and (_03078_, _03077_, _03071_);
  and (_03079_, _03078_, _02797_);
  and (_03080_, _03079_, _02791_);
  nor (_03081_, _03075_, _02795_);
  not (_03082_, _03081_);
  and (_03083_, _03082_, _02791_);
  or (_03084_, _03083_, _02786_);
  nor (_03085_, _03084_, _03080_);
  and (_03086_, _03085_, _02780_);
  and (_03087_, _02774_, _02752_);
  nor (_03088_, _03087_, _02775_);
  not (_03089_, _03088_);
  nor (_03090_, _03089_, _03086_);
  nor (_03091_, _03090_, _02775_);
  nor (_03092_, _03091_, _02771_);
  nor (_03093_, _03092_, _02770_);
  nor (_03094_, _03093_, _02760_);
  nor (_03095_, _03094_, _02757_);
  not (_03096_, _02596_);
  and (_03097_, _02752_, _03096_);
  nor (_03098_, _02752_, _03096_);
  nor (_03099_, _03098_, _03097_);
  and (_03100_, _03099_, _03095_);
  nor (_03101_, _03099_, _03095_);
  or (_03102_, _03101_, _03100_);
  or (_03103_, _03102_, _02630_);
  nand (_03104_, _02630_, _03096_);
  and (_03105_, _03104_, _02673_);
  and (_03106_, _03105_, _03103_);
  not (_03107_, _02675_);
  and (_03108_, _02645_, _01898_);
  and (_03109_, _02645_, _01935_);
  nor (_03110_, _03109_, _03108_);
  not (_03111_, \oc8051_golden_model_1.SP [2]);
  nor (_03112_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_03113_, _03112_, _03111_);
  nor (_03114_, _03112_, _03111_);
  nor (_03115_, _03114_, _03113_);
  nor (_03116_, _03115_, _03110_);
  not (_03117_, _03116_);
  not (_03118_, _01992_);
  and (_03119_, _03118_, _02674_);
  not (_03120_, _03119_);
  and (_03121_, _02023_, _01954_);
  not (_03122_, _02650_);
  and (_03123_, _02023_, _01970_);
  not (_03124_, _03123_);
  not (_03125_, _02647_);
  not (_03126_, _03108_);
  not (_03127_, _02405_);
  and (_03128_, _02023_, _01898_);
  and (_03129_, _03128_, _03127_);
  nor (_03130_, _02405_, _02204_);
  and (_03132_, _02295_, _02204_);
  nor (_03133_, _03132_, _03130_);
  and (_03134_, _02645_, _01966_);
  and (_03135_, _02645_, _01959_);
  nor (_03136_, _03135_, _03134_);
  nor (_03137_, _03136_, _03133_);
  not (_03139_, _02024_);
  and (_03140_, _02645_, _01983_);
  not (_03141_, _03140_);
  and (_03143_, _02566_, _02663_);
  and (_03144_, _02645_, _02663_);
  nor (_03146_, _03144_, _03143_);
  not (_03147_, _03146_);
  and (_03149_, _03147_, _03133_);
  and (_03150_, _02645_, _02660_);
  and (_03152_, _03150_, _03133_);
  not (_03153_, _01997_);
  and (_03154_, _02023_, _03153_);
  nor (_03156_, _03154_, _02661_);
  or (_03157_, _03156_, _02405_);
  not (_03159_, \oc8051_golden_model_1.PSW [3]);
  nand (_03160_, _03156_, _03159_);
  and (_03162_, _02566_, _02660_);
  nor (_03163_, _03162_, _03150_);
  and (_03165_, _03163_, _03160_);
  and (_03166_, _03165_, _03157_);
  not (_03167_, _01989_);
  and (_03168_, _02023_, _03167_);
  and (_03170_, _03162_, \oc8051_golden_model_1.SP [3]);
  or (_03171_, _03170_, _03168_);
  or (_03173_, _03171_, _03166_);
  or (_03174_, _03173_, _03152_);
  and (_03176_, _02645_, _03167_);
  not (_03177_, _03176_);
  not (_03179_, _03168_);
  or (_03181_, _03179_, _02405_);
  and (_03183_, _03181_, _03177_);
  and (_03184_, _03183_, _03174_);
  nand (_03186_, _03176_, _03133_);
  and (_03187_, _02566_, _03167_);
  nor (_03189_, _03187_, _02664_);
  nand (_03191_, _03189_, _03186_);
  or (_03192_, _03191_, _03184_);
  or (_03194_, _03189_, _02405_);
  and (_03195_, _03194_, _03146_);
  and (_03197_, _03195_, _03192_);
  nor (_03198_, _03197_, _03149_);
  nor (_03200_, _01992_, _02021_);
  nor (_03201_, _03200_, _03198_);
  and (_03203_, _02566_, _03118_);
  and (_03205_, _02645_, _03118_);
  nor (_03207_, _03205_, _03203_);
  not (_03209_, _03207_);
  and (_03211_, _03200_, _02405_);
  nor (_03213_, _03211_, _03209_);
  not (_03215_, _03213_);
  nor (_03217_, _03215_, _03201_);
  and (_03219_, _02023_, _01983_);
  nor (_03221_, _03207_, _03133_);
  nor (_03223_, _03221_, _03219_);
  not (_03224_, _03223_);
  nor (_03225_, _03224_, _03217_);
  and (_03226_, _03219_, _02405_);
  or (_03227_, _03226_, _03225_);
  and (_03228_, _03227_, _03141_);
  and (_03229_, _03140_, _03133_);
  or (_03230_, _03229_, _03228_);
  and (_03231_, _03230_, _03139_);
  not (_03232_, _03136_);
  nor (_03233_, _02945_, _03139_);
  nor (_03234_, _03233_, _03232_);
  not (_03235_, _03234_);
  nor (_03236_, _03235_, _03231_);
  nor (_03237_, _03236_, _03137_);
  and (_03238_, _02023_, _01942_);
  and (_03239_, _02645_, _01942_);
  nor (_03240_, _03239_, _02654_);
  not (_03241_, _03240_);
  nor (_03242_, _03241_, _03238_);
  and (_03243_, _02645_, _01964_);
  not (_03244_, _03243_);
  and (_03245_, _02023_, _01964_);
  nor (_03246_, _03245_, _02669_);
  and (_03247_, _03246_, _03244_);
  and (_03248_, _03247_, _03242_);
  and (_03249_, _02023_, _01935_);
  not (_03250_, _03249_);
  and (_03251_, _02645_, _01973_);
  not (_03252_, _03251_);
  and (_03253_, _02023_, _01973_);
  nor (_03254_, _03253_, _02656_);
  and (_03255_, _03254_, _03252_);
  and (_03256_, _03255_, _03250_);
  and (_03257_, _03256_, _03248_);
  not (_03258_, _03257_);
  nor (_03259_, _03258_, _03237_);
  nor (_03260_, _03257_, _02405_);
  nor (_03261_, _03260_, _03109_);
  not (_03262_, _03261_);
  nor (_03263_, _03262_, _03259_);
  and (_03264_, _03109_, \oc8051_golden_model_1.SP [3]);
  or (_03265_, _03264_, _02653_);
  or (_03266_, _03265_, _03263_);
  not (_03267_, _02653_);
  or (_03268_, _03133_, _03267_);
  and (_03269_, _03268_, _03266_);
  nor (_03270_, _03269_, _03128_);
  nor (_03271_, _03270_, _03129_);
  and (_03272_, _03271_, _03126_);
  and (_03273_, _03108_, \oc8051_golden_model_1.SP [3]);
  or (_03274_, _03273_, _03272_);
  and (_03275_, _03274_, _03125_);
  and (_03276_, _03133_, _02647_);
  or (_03277_, _03276_, _03275_);
  and (_03278_, _03277_, _03124_);
  and (_03279_, _03123_, _02405_);
  or (_03280_, _03279_, _03278_);
  and (_03281_, _03280_, _03122_);
  and (_03282_, _03133_, _02650_);
  nor (_03283_, _03282_, _03281_);
  nor (_03284_, _03283_, _03121_);
  and (_03285_, _03121_, _02405_);
  nor (_03286_, _03285_, _03284_);
  and (_03287_, _02650_, _02204_);
  and (_03288_, _03150_, _02204_);
  nor (_03289_, _03288_, _03287_);
  and (_03290_, _03207_, _03136_);
  and (_03291_, _03290_, _03146_);
  nor (_03292_, _03176_, _02647_);
  and (_03293_, _03292_, _03291_);
  nor (_03294_, _03293_, _02222_);
  not (_03295_, _03294_);
  and (_03296_, _03295_, _03289_);
  nor (_03297_, _03296_, _02333_);
  not (_03298_, _03297_);
  not (_03299_, _02333_);
  and (_03300_, _03140_, _02204_);
  and (_03301_, _03300_, _03299_);
  not (_03302_, _03301_);
  nor (_03303_, _02333_, _02222_);
  and (_03304_, _03303_, _02653_);
  not (_03305_, _03304_);
  and (_03306_, _03189_, _03156_);
  nor (_03307_, _03219_, _03200_);
  and (_03308_, _03307_, _03179_);
  and (_03309_, _03308_, _03306_);
  nor (_03310_, _03249_, _03121_);
  nor (_03311_, _03123_, _03128_);
  and (_03312_, _03311_, _03310_);
  and (_03313_, _03312_, _03255_);
  and (_03314_, _03313_, _03248_);
  and (_03315_, _03314_, _03309_);
  nor (_03316_, _03315_, _02439_);
  not (_03317_, _03316_);
  nor (_03318_, _02981_, _03139_);
  and (_03319_, _01920_, _02020_);
  not (_03320_, _03319_);
  nor (_03321_, _01970_, _01959_);
  and (_03322_, _03321_, _01984_);
  nor (_03323_, _03322_, _03320_);
  not (_03324_, _03323_);
  and (_03325_, _03153_, _02639_);
  and (_03326_, _01920_, _01981_);
  and (_03327_, _03326_, _03153_);
  nor (_03328_, _03327_, _03325_);
  and (_03329_, _01924_, _01704_);
  not (_03330_, _03329_);
  nor (_03331_, _01933_, _01940_);
  not (_03332_, _03331_);
  and (_03333_, _01989_, _01984_);
  and (_03334_, _03333_, _03332_);
  nor (_03335_, _03334_, _03330_);
  not (_03336_, _03335_);
  and (_03337_, _03336_, _03328_);
  and (_03338_, _03337_, _03324_);
  or (_03339_, _03329_, _03319_);
  and (_03340_, _03339_, _01898_);
  not (_03341_, _03340_);
  nor (_03342_, _01994_, _01926_);
  and (_03343_, _01954_, _03329_);
  nor (_03344_, _03343_, _03342_);
  and (_03345_, _03344_, _03341_);
  and (_03346_, _01970_, _03329_);
  nor (_03347_, _03346_, _02666_);
  and (_03348_, _01942_, _03329_);
  and (_03349_, _02565_, _01920_);
  and (_03350_, _01970_, _03349_);
  nor (_03351_, _03350_, _03348_);
  and (_03352_, _03351_, _03347_);
  and (_03353_, _03352_, _03345_);
  not (_03354_, _03349_);
  nor (_03355_, _01959_, _01898_);
  and (_03356_, _03355_, _01984_);
  nor (_03357_, _03356_, _03354_);
  not (_03358_, _02665_);
  not (_03359_, _01964_);
  nor (_03360_, _01954_, _01935_);
  and (_03361_, _03360_, _03359_);
  nor (_03362_, _03361_, _03358_);
  nor (_03363_, _03362_, _03357_);
  and (_03364_, _03363_, _03353_);
  not (_03365_, _03162_);
  and (_03366_, _03365_, _03110_);
  nor (_03367_, _03366_, _03111_);
  not (_03368_, _03367_);
  nor (_03369_, _01964_, _01959_);
  nor (_03370_, _03369_, _03330_);
  not (_03371_, _03370_);
  nor (_03372_, _03167_, _01942_);
  nor (_03373_, _03372_, _03358_);
  and (_03374_, _01973_, _01920_);
  nor (_03375_, _03374_, _03373_);
  and (_03376_, _03375_, _03371_);
  and (_03377_, _03376_, _03368_);
  and (_03378_, _03377_, _03364_);
  and (_03379_, _03378_, _03338_);
  not (_03380_, _03379_);
  nor (_03381_, _03380_, _03318_);
  and (_03382_, _03381_, _03317_);
  and (_03383_, _03382_, _03305_);
  and (_03384_, _03383_, _03302_);
  and (_03385_, _03384_, _03298_);
  not (_03386_, \oc8051_golden_model_1.IRAM[0] [2]);
  not (_03387_, _02664_);
  nor (_03388_, _03387_, _02503_);
  or (_03389_, _03179_, _02503_);
  not (_03390_, _03150_);
  and (_03391_, _02405_, _02204_);
  or (_03392_, _03391_, _03390_);
  nor (_03393_, _03156_, _02503_);
  not (_03394_, _01987_);
  and (_03395_, _02022_, _02631_);
  or (_03396_, _03395_, _02645_);
  and (_03397_, _03396_, _03394_);
  not (_03398_, _03397_);
  not (_03399_, _01736_);
  nor (_03400_, _01925_, _03399_);
  and (_03401_, _03400_, _03153_);
  nor (_03402_, _03401_, _03154_);
  and (_03403_, _03402_, _03398_);
  and (_03404_, _02660_, _02640_);
  or (_03405_, _01767_, _01673_);
  nor (_03406_, _01994_, _02021_);
  and (_03407_, _03406_, _01736_);
  and (_03408_, _03407_, _03405_);
  and (_03409_, _03395_, _02660_);
  and (_03410_, _02645_, _03153_);
  or (_03411_, _03410_, _02661_);
  or (_03412_, _03411_, _03409_);
  or (_03413_, _03412_, _03408_);
  nor (_03414_, _03413_, _03404_);
  and (_03415_, _03414_, _03403_);
  or (_03416_, _03415_, _03393_);
  not (_03417_, \oc8051_golden_model_1.SP [0]);
  and (_03418_, _03162_, _03417_);
  nor (_03419_, _03418_, _03168_);
  and (_03420_, _03395_, _03167_);
  and (_03421_, _01736_, _01704_);
  and (_03422_, _03167_, _03421_);
  nor (_03423_, _03422_, _03420_);
  and (_03424_, _03423_, _03419_);
  and (_03425_, _03424_, _03416_);
  nand (_03426_, _03425_, _03392_);
  nand (_03427_, _03426_, _03389_);
  nor (_03428_, _03187_, _03176_);
  nand (_03429_, _03428_, _03427_);
  not (_03430_, _03187_);
  or (_03431_, _03430_, _02503_);
  nand (_03432_, _03391_, _03176_);
  and (_03433_, _03432_, _03431_);
  and (_03434_, _03433_, _03429_);
  nor (_03435_, _03400_, _02023_);
  nor (_03436_, _03435_, _01999_);
  nor (_03437_, _03436_, _03434_);
  or (_03438_, _03437_, _03388_);
  and (_03439_, _03438_, _03146_);
  and (_03440_, _03391_, _03147_);
  or (_03441_, _03440_, _03439_);
  and (_03442_, _03200_, _02503_);
  and (_03443_, _03395_, _03118_);
  nor (_03444_, _03443_, _03209_);
  not (_03445_, _03444_);
  nor (_03446_, _03445_, _03442_);
  and (_03447_, _03446_, _03441_);
  and (_03448_, _03391_, _03209_);
  nor (_03449_, _03448_, _03447_);
  nor (_03450_, _03435_, _01984_);
  nor (_03451_, _03450_, _03449_);
  not (_03452_, _02503_);
  and (_03453_, _03219_, _03452_);
  or (_03454_, _03453_, _03451_);
  and (_03455_, _03454_, _03141_);
  and (_03456_, _03391_, _03140_);
  nor (_03457_, _03456_, _03455_);
  nor (_03458_, _03435_, _02029_);
  nor (_03459_, _03458_, _03457_);
  nor (_03460_, _03048_, _03139_);
  or (_03461_, _03460_, _03459_);
  not (_03462_, _03135_);
  nor (_03463_, _03391_, _03462_);
  and (_03464_, _03396_, _01966_);
  nor (_03465_, _03464_, _03463_);
  and (_03466_, _03465_, _03461_);
  and (_03467_, _03391_, _03134_);
  or (_03468_, _03467_, _03466_);
  and (_03469_, _03395_, _01973_);
  and (_03470_, _01973_, _03421_);
  nor (_03471_, _03470_, _03469_);
  and (_03472_, _03471_, _03468_);
  nor (_03473_, _03255_, _03452_);
  and (_03474_, _03400_, _01964_);
  nor (_03475_, _03474_, _03473_);
  and (_03476_, _03475_, _03472_);
  nor (_03477_, _03247_, _03452_);
  and (_03478_, _03400_, _01942_);
  nor (_03479_, _03478_, _03477_);
  and (_03480_, _03479_, _03476_);
  nor (_03481_, _03242_, _03452_);
  not (_03482_, _01935_);
  nor (_03483_, _03435_, _03482_);
  nor (_03484_, _03483_, _03481_);
  and (_03485_, _03484_, _03480_);
  nor (_03486_, _03250_, _02503_);
  or (_03487_, _03486_, _03485_);
  and (_03488_, _03109_, _03417_);
  nor (_03489_, _03488_, _02653_);
  and (_03490_, _03489_, _03487_);
  and (_03491_, _03391_, _02653_);
  nor (_03492_, _03491_, _03490_);
  nor (_03493_, _03435_, _01915_);
  nor (_03494_, _03493_, _03492_);
  and (_03495_, _03128_, _03452_);
  or (_03496_, _03495_, _03494_);
  and (_03497_, _03108_, _03417_);
  nor (_03498_, _03497_, _02647_);
  and (_03499_, _03498_, _03496_);
  and (_03500_, _03391_, _02647_);
  nor (_03501_, _03500_, _03499_);
  not (_03502_, _01970_);
  nor (_03503_, _03435_, _03502_);
  nor (_03504_, _03503_, _03501_);
  nor (_03505_, _03124_, _02503_);
  or (_03506_, _03505_, _03504_);
  and (_03507_, _03506_, _03122_);
  and (_03508_, _03391_, _02650_);
  nor (_03509_, _03508_, _03507_);
  not (_03510_, _01954_);
  nor (_03511_, _03435_, _03510_);
  or (_03512_, _03511_, _03509_);
  not (_03513_, _03121_);
  nor (_03514_, _03513_, _02503_);
  not (_03515_, _03514_);
  nand (_03516_, _03515_, _03512_);
  or (_03517_, _03516_, _03386_);
  not (_03518_, _02370_);
  and (_03519_, _03300_, _03518_);
  not (_03520_, _03519_);
  nor (_03521_, _02370_, _02222_);
  nor (_03522_, _02647_, _02650_);
  nor (_03523_, _03176_, _02653_);
  and (_03524_, _03523_, _03390_);
  and (_03525_, _03524_, _03522_);
  and (_03526_, _03525_, _03291_);
  not (_03527_, _03526_);
  and (_03528_, _03527_, _03521_);
  not (_03529_, _03528_);
  nor (_03530_, _03315_, _02471_);
  not (_03531_, _03530_);
  nor (_03532_, _03016_, _03139_);
  not (_03533_, _01918_);
  or (_03534_, _01983_, _01964_);
  nand (_03535_, _01999_, _01989_);
  or (_03536_, _03535_, _03534_);
  and (_03537_, _03536_, _03533_);
  nor (_03538_, _02029_, _01918_);
  or (_03539_, _03538_, _01919_);
  or (_03540_, _03539_, _03537_);
  and (_03541_, _01935_, _02632_);
  and (_03542_, _01767_, _01704_);
  or (_03543_, _02660_, _01973_);
  and (_03544_, _03543_, _03542_);
  or (_03545_, _03544_, _03541_);
  and (_03546_, _01970_, _02632_);
  and (_03547_, _01970_, _01917_);
  and (_03548_, _03547_, _02635_);
  or (_03549_, _03548_, _03546_);
  or (_03550_, _03549_, _03545_);
  nor (_03551_, _01943_, _01918_);
  and (_03552_, _03542_, _03153_);
  and (_03553_, _01954_, _03533_);
  or (_03554_, _03553_, _03552_);
  or (_03555_, _03554_, _03551_);
  or (_03556_, _03346_, _03348_);
  and (_03557_, _01935_, _02636_);
  or (_03558_, _03557_, _03343_);
  or (_03559_, _03558_, _03556_);
  or (_03560_, _03559_, _03555_);
  or (_03561_, _03560_, _03550_);
  and (_03562_, _03369_, _01915_);
  nand (_03563_, _03562_, _03334_);
  and (_03564_, _03563_, _03329_);
  not (_03565_, \oc8051_golden_model_1.SP [1]);
  nor (_03566_, _03366_, _03565_);
  or (_03567_, _03566_, _03564_);
  or (_03568_, _03567_, _03561_);
  nor (_03569_, _03568_, _03540_);
  not (_03570_, _03569_);
  nor (_03571_, _03570_, _03532_);
  and (_03572_, _03571_, _03531_);
  and (_03573_, _03572_, _03529_);
  and (_03574_, _03573_, _03520_);
  not (_03575_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_03576_, _03515_, _03512_);
  or (_03577_, _03576_, _03575_);
  and (_03578_, _03577_, _03574_);
  nand (_03579_, _03578_, _03517_);
  not (_03580_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_03581_, _03576_, _03580_);
  not (_03582_, _03574_);
  not (_03583_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_03584_, _03516_, _03583_);
  and (_03585_, _03584_, _03582_);
  nand (_03586_, _03585_, _03581_);
  nand (_03587_, _03586_, _03579_);
  nand (_03588_, _03587_, _03385_);
  not (_03589_, _03385_);
  not (_03590_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_03591_, _03576_, _03590_);
  not (_03592_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_03593_, _03516_, _03592_);
  and (_03594_, _03593_, _03582_);
  nand (_03595_, _03594_, _03591_);
  not (_03596_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_03597_, _03516_, _03596_);
  not (_03598_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_03599_, _03576_, _03598_);
  and (_03600_, _03599_, _03574_);
  nand (_03601_, _03600_, _03597_);
  nand (_03602_, _03601_, _03595_);
  nand (_03603_, _03602_, _03589_);
  nand (_03605_, _03603_, _03588_);
  nand (_03607_, _03605_, _03286_);
  not (_03609_, _03286_);
  nand (_03611_, _03516_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_03613_, _03576_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_03615_, _03613_, _03582_);
  nand (_03617_, _03615_, _03611_);
  nand (_03619_, _03576_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_03621_, _03516_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_03623_, _03621_, _03574_);
  nand (_03625_, _03623_, _03619_);
  nand (_03627_, _03625_, _03617_);
  nand (_03629_, _03627_, _03385_);
  nand (_03631_, _03516_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_03633_, _03576_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_03634_, _03633_, _03582_);
  nand (_03635_, _03634_, _03631_);
  nand (_03636_, _03576_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_03637_, _03516_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_03638_, _03637_, _03574_);
  nand (_03639_, _03638_, _03636_);
  nand (_03640_, _03639_, _03635_);
  nand (_03641_, _03640_, _03589_);
  nand (_03642_, _03641_, _03629_);
  nand (_03643_, _03642_, _03609_);
  nand (_03644_, _03643_, _03607_);
  nand (_03645_, _03644_, _03120_);
  not (_03646_, _03110_);
  and (_03647_, _03119_, _02439_);
  nor (_03648_, _03647_, _03646_);
  nand (_03649_, _03648_, _03645_);
  and (_03650_, _03649_, _03117_);
  nand (_03651_, _03385_, \oc8051_golden_model_1.IRAM[3] [0]);
  nand (_03652_, _03589_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_03653_, _03652_, _03651_);
  or (_03654_, _03653_, _03576_);
  nand (_03655_, _03385_, \oc8051_golden_model_1.IRAM[2] [0]);
  nand (_03656_, _03589_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_03657_, _03656_, _03655_);
  or (_03658_, _03657_, _03516_);
  and (_03659_, _03658_, _03582_);
  and (_03660_, _03659_, _03654_);
  nand (_03661_, _03385_, \oc8051_golden_model_1.IRAM[1] [0]);
  nand (_03662_, _03589_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_03663_, _03662_, _03661_);
  or (_03665_, _03663_, _03576_);
  nand (_03667_, _03385_, \oc8051_golden_model_1.IRAM[0] [0]);
  nand (_03669_, _03589_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_03671_, _03669_, _03667_);
  or (_03673_, _03671_, _03516_);
  and (_03675_, _03673_, _03574_);
  and (_03677_, _03675_, _03665_);
  or (_03679_, _03677_, _03660_);
  nand (_03681_, _03679_, _03286_);
  not (_03683_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_03685_, _03516_, _03683_);
  not (_03687_, \oc8051_golden_model_1.IRAM[9] [0]);
  or (_03689_, _03576_, _03687_);
  and (_03691_, _03689_, _03574_);
  nand (_03693_, _03691_, _03685_);
  not (_03694_, \oc8051_golden_model_1.IRAM[11] [0]);
  or (_03695_, _03576_, _03694_);
  nand (_03696_, _03576_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_03697_, _03696_, _03582_);
  nand (_03698_, _03697_, _03695_);
  nand (_03699_, _03698_, _03693_);
  nand (_03700_, _03699_, _03385_);
  not (_03701_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_03702_, _03576_, _03701_);
  nand (_03703_, _03576_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_03704_, _03703_, _03582_);
  nand (_03705_, _03704_, _03702_);
  not (_03706_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_03707_, _03516_, _03706_);
  not (_03708_, \oc8051_golden_model_1.IRAM[13] [0]);
  or (_03709_, _03576_, _03708_);
  and (_03710_, _03709_, _03574_);
  nand (_03711_, _03710_, _03707_);
  nand (_03712_, _03711_, _03705_);
  nand (_03713_, _03712_, _03589_);
  nand (_03714_, _03713_, _03700_);
  nand (_03715_, _03714_, _03609_);
  and (_03716_, _03715_, _03681_);
  or (_03717_, _03716_, _03119_);
  and (_03718_, _03119_, _02503_);
  nor (_03719_, _03718_, _03646_);
  nand (_03720_, _03719_, _03717_);
  nor (_03721_, _03110_, \oc8051_golden_model_1.SP [0]);
  not (_03722_, _03721_);
  and (_03723_, _03722_, _03720_);
  nand (_03724_, _03723_, \oc8051_golden_model_1.IRAM[0] [5]);
  not (_03725_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_03726_, _03516_, _03725_);
  not (_03727_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_03728_, _03576_, _03727_);
  and (_03729_, _03728_, _03574_);
  nand (_03730_, _03729_, _03726_);
  not (_03731_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_03732_, _03576_, _03731_);
  not (_03733_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_03734_, _03516_, _03733_);
  and (_03735_, _03734_, _03582_);
  nand (_03736_, _03735_, _03732_);
  nand (_03737_, _03736_, _03730_);
  nand (_03738_, _03737_, _03385_);
  not (_03739_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_03740_, _03576_, _03739_);
  not (_03741_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_03742_, _03516_, _03741_);
  and (_03743_, _03742_, _03582_);
  nand (_03744_, _03743_, _03740_);
  not (_03745_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_03746_, _03516_, _03745_);
  not (_03747_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_03748_, _03576_, _03747_);
  and (_03749_, _03748_, _03574_);
  nand (_03750_, _03749_, _03746_);
  nand (_03751_, _03750_, _03744_);
  nand (_03752_, _03751_, _03589_);
  nand (_03753_, _03752_, _03738_);
  nand (_03754_, _03753_, _03286_);
  nand (_03755_, _03516_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_03756_, _03576_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_03757_, _03756_, _03582_);
  nand (_03758_, _03757_, _03755_);
  nand (_03759_, _03576_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand (_03760_, _03516_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_03761_, _03760_, _03574_);
  nand (_03762_, _03761_, _03759_);
  nand (_03763_, _03762_, _03758_);
  nand (_03764_, _03763_, _03385_);
  nand (_03765_, _03516_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_03766_, _03576_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_03767_, _03766_, _03582_);
  nand (_03768_, _03767_, _03765_);
  nand (_03769_, _03576_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand (_03770_, _03516_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_03771_, _03770_, _03574_);
  nand (_03772_, _03771_, _03769_);
  nand (_03773_, _03772_, _03768_);
  nand (_03774_, _03773_, _03589_);
  nand (_03775_, _03774_, _03764_);
  nand (_03776_, _03775_, _03609_);
  nand (_03777_, _03776_, _03754_);
  or (_03778_, _03777_, _03119_);
  nor (_03779_, _03120_, _02471_);
  nor (_03780_, _03779_, _03646_);
  nand (_03781_, _03780_, _03778_);
  and (_03782_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  nor (_03783_, _03782_, _03112_);
  not (_03784_, _03783_);
  nor (_03785_, _03784_, _03110_);
  not (_03786_, _03785_);
  and (_03787_, _03786_, _03781_);
  not (_03788_, _03787_);
  not (_03789_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_03790_, _03723_, _03789_);
  and (_03791_, _03790_, _03788_);
  nand (_03792_, _03791_, _03724_);
  nand (_03793_, _03723_, \oc8051_golden_model_1.IRAM[2] [5]);
  not (_03794_, \oc8051_golden_model_1.IRAM[3] [5]);
  or (_03795_, _03723_, _03794_);
  and (_03796_, _03795_, _03787_);
  nand (_03797_, _03796_, _03793_);
  nand (_03798_, _03797_, _03792_);
  nand (_03799_, _03798_, _03650_);
  not (_03800_, \oc8051_golden_model_1.SP [3]);
  nor (_03801_, _03113_, _03800_);
  nor (_03802_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_03803_, _03802_, _03800_);
  and (_03804_, _03803_, _03417_);
  nor (_03805_, _03804_, _03801_);
  nor (_03806_, _03805_, _03110_);
  not (_03807_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_03808_, _03516_, _03807_);
  not (_03809_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_03810_, _03576_, _03809_);
  and (_03811_, _03810_, _03574_);
  nand (_03812_, _03811_, _03808_);
  not (_03813_, \oc8051_golden_model_1.IRAM[3] [3]);
  or (_03814_, _03576_, _03813_);
  not (_03815_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_03816_, _03516_, _03815_);
  and (_03817_, _03816_, _03582_);
  nand (_03818_, _03817_, _03814_);
  nand (_03819_, _03818_, _03812_);
  nand (_03820_, _03819_, _03385_);
  not (_03821_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_03822_, _03576_, _03821_);
  not (_03823_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_03824_, _03516_, _03823_);
  and (_03825_, _03824_, _03582_);
  nand (_03826_, _03825_, _03822_);
  not (_03827_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_03828_, _03516_, _03827_);
  not (_03829_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_03830_, _03576_, _03829_);
  and (_03831_, _03830_, _03574_);
  nand (_03832_, _03831_, _03828_);
  nand (_03833_, _03832_, _03826_);
  nand (_03834_, _03833_, _03589_);
  nand (_03835_, _03834_, _03820_);
  nand (_03836_, _03835_, _03286_);
  nand (_03837_, _03516_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_03838_, _03576_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_03839_, _03838_, _03582_);
  nand (_03840_, _03839_, _03837_);
  nand (_03841_, _03576_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_03842_, _03516_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_03843_, _03842_, _03574_);
  nand (_03844_, _03843_, _03841_);
  nand (_03845_, _03844_, _03840_);
  nand (_03846_, _03845_, _03385_);
  nand (_03847_, _03516_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_03848_, _03576_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_03849_, _03848_, _03582_);
  nand (_03850_, _03849_, _03847_);
  nand (_03851_, _03576_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand (_03852_, _03516_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_03853_, _03852_, _03574_);
  nand (_03854_, _03853_, _03851_);
  nand (_03855_, _03854_, _03850_);
  nand (_03856_, _03855_, _03589_);
  nand (_03857_, _03856_, _03846_);
  nand (_03858_, _03857_, _03609_);
  nand (_03859_, _03858_, _03836_);
  and (_03860_, _03859_, _03120_);
  nor (_03861_, _03120_, _02405_);
  or (_03862_, _03861_, _03646_);
  nor (_03863_, _03862_, _03860_);
  nor (_03864_, _03863_, _03806_);
  not (_03865_, _03650_);
  nand (_03866_, _03723_, \oc8051_golden_model_1.IRAM[4] [5]);
  not (_03867_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_03868_, _03723_, _03867_);
  and (_03869_, _03868_, _03788_);
  nand (_03870_, _03869_, _03866_);
  nand (_03871_, _03723_, \oc8051_golden_model_1.IRAM[6] [5]);
  not (_03872_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_03873_, _03723_, _03872_);
  and (_03874_, _03873_, _03787_);
  nand (_03875_, _03874_, _03871_);
  nand (_03876_, _03875_, _03870_);
  nand (_03877_, _03876_, _03865_);
  and (_03878_, _03877_, _03864_);
  and (_03879_, _03878_, _03799_);
  not (_03880_, _03723_);
  or (_03881_, _03880_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_03882_, _03723_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_03883_, _03882_, _03881_);
  nand (_03884_, _03883_, _03787_);
  or (_03885_, _03880_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_03886_, _03723_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand (_03887_, _03886_, _03885_);
  nand (_03888_, _03887_, _03788_);
  nand (_03889_, _03888_, _03884_);
  nand (_03890_, _03889_, _03650_);
  not (_03891_, _03864_);
  or (_03892_, _03880_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_03893_, _03723_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_03894_, _03893_, _03892_);
  nand (_03895_, _03894_, _03787_);
  or (_03896_, _03880_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_03897_, _03723_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand (_03898_, _03897_, _03896_);
  nand (_03899_, _03898_, _03788_);
  nand (_03900_, _03899_, _03895_);
  nand (_03901_, _03900_, _03865_);
  and (_03902_, _03901_, _03891_);
  and (_03903_, _03902_, _03890_);
  or (_03904_, _03903_, _03879_);
  or (_03905_, _03904_, _02333_);
  nor (_03906_, _03903_, _03879_);
  or (_03907_, _03906_, _03299_);
  and (_03908_, _03907_, _03905_);
  not (_03909_, _02295_);
  nand (_03910_, _03723_, \oc8051_golden_model_1.IRAM[0] [6]);
  not (_03911_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_03912_, _03723_, _03911_);
  and (_03913_, _03912_, _03788_);
  nand (_03914_, _03913_, _03910_);
  nand (_03915_, _03723_, \oc8051_golden_model_1.IRAM[2] [6]);
  not (_03916_, \oc8051_golden_model_1.IRAM[3] [6]);
  or (_03917_, _03723_, _03916_);
  and (_03918_, _03917_, _03787_);
  nand (_03919_, _03918_, _03915_);
  nand (_03920_, _03919_, _03914_);
  nand (_03921_, _03920_, _03650_);
  nand (_03922_, _03723_, \oc8051_golden_model_1.IRAM[4] [6]);
  not (_03923_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_03924_, _03723_, _03923_);
  and (_03925_, _03924_, _03788_);
  nand (_03926_, _03925_, _03922_);
  nand (_03927_, _03723_, \oc8051_golden_model_1.IRAM[6] [6]);
  not (_03928_, \oc8051_golden_model_1.IRAM[7] [6]);
  or (_03929_, _03723_, _03928_);
  and (_03930_, _03929_, _03787_);
  nand (_03931_, _03930_, _03927_);
  nand (_03932_, _03931_, _03926_);
  nand (_03933_, _03932_, _03865_);
  and (_03934_, _03933_, _03864_);
  and (_03935_, _03934_, _03921_);
  or (_03936_, _03880_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_03937_, _03723_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_03938_, _03937_, _03936_);
  nand (_03939_, _03938_, _03787_);
  or (_03940_, _03880_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_03941_, _03723_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand (_03942_, _03941_, _03940_);
  nand (_03943_, _03942_, _03788_);
  nand (_03944_, _03943_, _03939_);
  nand (_03945_, _03944_, _03650_);
  or (_03946_, _03880_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_03947_, _03723_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_03948_, _03947_, _03946_);
  nand (_03949_, _03948_, _03787_);
  or (_03950_, _03880_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_03951_, _03723_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand (_03952_, _03951_, _03950_);
  nand (_03953_, _03952_, _03788_);
  nand (_03954_, _03953_, _03949_);
  nand (_03955_, _03954_, _03865_);
  and (_03956_, _03955_, _03891_);
  and (_03957_, _03956_, _03945_);
  nor (_03958_, _03957_, _03935_);
  or (_03959_, _03958_, _03909_);
  or (_03960_, _03957_, _03935_);
  or (_03961_, _03960_, _02295_);
  and (_03962_, _03961_, _03959_);
  and (_03963_, _03962_, _03908_);
  nand (_03964_, _03723_, \oc8051_golden_model_1.IRAM[0] [4]);
  not (_03965_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_03966_, _03723_, _03965_);
  and (_03967_, _03966_, _03788_);
  nand (_03968_, _03967_, _03964_);
  nand (_03969_, _03723_, \oc8051_golden_model_1.IRAM[2] [4]);
  not (_03970_, \oc8051_golden_model_1.IRAM[3] [4]);
  or (_03971_, _03723_, _03970_);
  and (_03972_, _03971_, _03787_);
  nand (_03973_, _03972_, _03969_);
  nand (_03974_, _03973_, _03968_);
  nand (_03975_, _03974_, _03650_);
  nand (_03976_, _03723_, \oc8051_golden_model_1.IRAM[4] [4]);
  not (_03977_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_03978_, _03723_, _03977_);
  and (_03979_, _03978_, _03788_);
  nand (_03980_, _03979_, _03976_);
  nand (_03981_, _03723_, \oc8051_golden_model_1.IRAM[6] [4]);
  not (_03982_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_03983_, _03723_, _03982_);
  and (_03984_, _03983_, _03787_);
  nand (_03985_, _03984_, _03981_);
  nand (_03986_, _03985_, _03980_);
  nand (_03987_, _03986_, _03865_);
  and (_03988_, _03987_, _03864_);
  and (_03989_, _03988_, _03975_);
  or (_03990_, _03880_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_03991_, _03723_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_03992_, _03991_, _03990_);
  nand (_03993_, _03992_, _03787_);
  or (_03994_, _03880_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_03995_, _03723_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand (_03996_, _03995_, _03994_);
  nand (_03997_, _03996_, _03788_);
  nand (_03998_, _03997_, _03993_);
  nand (_03999_, _03998_, _03650_);
  or (_04000_, _03880_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_04001_, _03723_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_04002_, _04001_, _04000_);
  nand (_04003_, _04002_, _03787_);
  or (_04004_, _03880_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_04005_, _03723_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand (_04006_, _04005_, _04004_);
  nand (_04007_, _04006_, _03788_);
  nand (_04008_, _04007_, _04003_);
  nand (_04009_, _04008_, _03865_);
  and (_04010_, _04009_, _03891_);
  and (_04011_, _04010_, _03999_);
  or (_04012_, _04011_, _03989_);
  or (_04013_, _04012_, _02370_);
  nor (_04014_, _04011_, _03989_);
  or (_04015_, _04014_, _03518_);
  and (_04016_, _04015_, _04013_);
  nand (_04017_, _03723_, \oc8051_golden_model_1.IRAM[0] [7]);
  not (_04018_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_04019_, _03723_, _04018_);
  and (_04020_, _04019_, _03788_);
  nand (_04021_, _04020_, _04017_);
  nand (_04022_, _03723_, \oc8051_golden_model_1.IRAM[2] [7]);
  not (_04023_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_04024_, _03723_, _04023_);
  and (_04025_, _04024_, _03787_);
  nand (_04026_, _04025_, _04022_);
  nand (_04027_, _04026_, _04021_);
  nand (_04028_, _04027_, _03650_);
  nand (_04029_, _03723_, \oc8051_golden_model_1.IRAM[4] [7]);
  not (_04030_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_04031_, _03723_, _04030_);
  and (_04032_, _04031_, _03788_);
  nand (_04033_, _04032_, _04029_);
  nand (_04034_, _03723_, \oc8051_golden_model_1.IRAM[6] [7]);
  not (_04035_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_04036_, _03723_, _04035_);
  and (_04037_, _04036_, _03787_);
  nand (_04038_, _04037_, _04034_);
  nand (_04039_, _04038_, _04033_);
  nand (_04040_, _04039_, _03865_);
  and (_04041_, _04040_, _03864_);
  and (_04042_, _04041_, _04028_);
  or (_04043_, _03880_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_04044_, _03723_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand (_04045_, _04044_, _04043_);
  nand (_04046_, _04045_, _03787_);
  nand (_04047_, _03723_, \oc8051_golden_model_1.IRAM[8] [7]);
  not (_04048_, \oc8051_golden_model_1.IRAM[9] [7]);
  or (_04049_, _03723_, _04048_);
  and (_04050_, _04049_, _04047_);
  nand (_04051_, _04050_, _03788_);
  nand (_04052_, _04051_, _04046_);
  nand (_04053_, _04052_, _03650_);
  not (_04054_, \oc8051_golden_model_1.IRAM[14] [7]);
  nand (_04055_, _03723_, _04054_);
  or (_04056_, _03723_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand (_04057_, _04056_, _04055_);
  nand (_04058_, _04057_, _03787_);
  or (_04059_, _03880_, \oc8051_golden_model_1.IRAM[12] [7]);
  or (_04060_, _03723_, \oc8051_golden_model_1.IRAM[13] [7]);
  nand (_04061_, _04060_, _04059_);
  nand (_04062_, _04061_, _03788_);
  nand (_04063_, _04062_, _04058_);
  nand (_04064_, _04063_, _03865_);
  and (_04065_, _04064_, _03891_);
  and (_04066_, _04065_, _04053_);
  or (_04067_, _04066_, _04042_);
  or (_04068_, _04067_, _02204_);
  nor (_04069_, _04066_, _04042_);
  or (_04070_, _04069_, _02222_);
  and (_04071_, _04070_, _04068_);
  and (_04072_, _04071_, _04016_);
  and (_04073_, _04072_, _03963_);
  nand (_04074_, _03723_, \oc8051_golden_model_1.IRAM[0] [3]);
  or (_04075_, _03723_, _03809_);
  and (_04076_, _04075_, _03788_);
  nand (_04077_, _04076_, _04074_);
  nand (_04078_, _03723_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_04079_, _03723_, _03813_);
  and (_04080_, _04079_, _03787_);
  nand (_04081_, _04080_, _04078_);
  nand (_04082_, _04081_, _04077_);
  nand (_04083_, _04082_, _03650_);
  nand (_04084_, _03723_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_04085_, _03723_, _03829_);
  and (_04086_, _04085_, _03788_);
  nand (_04087_, _04086_, _04084_);
  nand (_04088_, _03723_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_04089_, _03723_, _03821_);
  and (_04090_, _04089_, _03787_);
  nand (_04091_, _04090_, _04088_);
  nand (_04092_, _04091_, _04087_);
  nand (_04093_, _04092_, _03865_);
  and (_04094_, _04093_, _03864_);
  and (_04095_, _04094_, _04083_);
  or (_04096_, _03880_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_04097_, _03723_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_04098_, _04097_, _04096_);
  nand (_04099_, _04098_, _03787_);
  or (_04100_, _03880_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_04101_, _03723_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_04102_, _04101_, _04100_);
  nand (_04103_, _04102_, _03788_);
  nand (_04104_, _04103_, _04099_);
  nand (_04105_, _04104_, _03650_);
  or (_04106_, _03880_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_04107_, _03723_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_04108_, _04107_, _04106_);
  nand (_04109_, _04108_, _03787_);
  or (_04110_, _03880_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_04111_, _03723_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand (_04112_, _04111_, _04110_);
  nand (_04113_, _04112_, _03788_);
  nand (_04114_, _04113_, _04109_);
  nand (_04115_, _04114_, _03865_);
  and (_04116_, _04115_, _03891_);
  and (_04117_, _04116_, _04105_);
  nor (_04118_, _04117_, _04095_);
  and (_04119_, _04118_, _02405_);
  or (_04120_, _04117_, _04095_);
  and (_04121_, _04120_, _03127_);
  nor (_04122_, _04121_, _04119_);
  not (_04123_, _02439_);
  nand (_04124_, _03723_, \oc8051_golden_model_1.IRAM[0] [2]);
  or (_04125_, _03723_, _03575_);
  and (_04126_, _04125_, _03788_);
  nand (_04127_, _04126_, _04124_);
  nand (_04128_, _03723_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_04129_, _03723_, _03580_);
  and (_04130_, _04129_, _03787_);
  nand (_04131_, _04130_, _04128_);
  nand (_04132_, _04131_, _04127_);
  nand (_04133_, _04132_, _03650_);
  nand (_04134_, _03723_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_04135_, _03723_, _03598_);
  and (_04136_, _04135_, _03788_);
  nand (_04137_, _04136_, _04134_);
  nand (_04138_, _03723_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_04139_, _03723_, _03590_);
  and (_04140_, _04139_, _03787_);
  nand (_04141_, _04140_, _04138_);
  nand (_04142_, _04141_, _04137_);
  nand (_04143_, _04142_, _03865_);
  and (_04144_, _04143_, _03864_);
  and (_04145_, _04144_, _04133_);
  or (_04146_, _03880_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_04147_, _03723_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_04148_, _04147_, _04146_);
  nand (_04149_, _04148_, _03787_);
  or (_04150_, _03880_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_04151_, _03723_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_04152_, _04151_, _04150_);
  nand (_04153_, _04152_, _03788_);
  nand (_04154_, _04153_, _04149_);
  nand (_04155_, _04154_, _03650_);
  or (_04156_, _03880_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_04157_, _03723_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_04158_, _04157_, _04156_);
  nand (_04159_, _04158_, _03787_);
  or (_04160_, _03880_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_04161_, _03723_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_04162_, _04161_, _04160_);
  nand (_04163_, _04162_, _03788_);
  nand (_04164_, _04163_, _04159_);
  nand (_04165_, _04164_, _03865_);
  and (_04166_, _04165_, _03891_);
  and (_04167_, _04166_, _04155_);
  nor (_04168_, _04167_, _04145_);
  or (_04169_, _04168_, _04123_);
  or (_04170_, _04167_, _04145_);
  or (_04171_, _04170_, _02439_);
  and (_04172_, _04171_, _04169_);
  and (_04173_, _04172_, _04122_);
  nand (_04174_, _03723_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_04175_, _03723_, _03727_);
  and (_04176_, _04175_, _03788_);
  nand (_04177_, _04176_, _04174_);
  nand (_04178_, _03723_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_04179_, _03723_, _03731_);
  and (_04180_, _04179_, _03787_);
  nand (_04181_, _04180_, _04178_);
  nand (_04182_, _04181_, _04177_);
  nand (_04183_, _04182_, _03650_);
  nand (_04184_, _03723_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_04185_, _03723_, _03747_);
  and (_04186_, _04185_, _03788_);
  nand (_04187_, _04186_, _04184_);
  nand (_04188_, _03723_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_04189_, _03723_, _03739_);
  and (_04190_, _04189_, _03787_);
  nand (_04191_, _04190_, _04188_);
  nand (_04192_, _04191_, _04187_);
  nand (_04193_, _04192_, _03865_);
  and (_04194_, _04193_, _03864_);
  and (_04195_, _04194_, _04183_);
  or (_04196_, _03880_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_04197_, _03723_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_04198_, _04197_, _04196_);
  nand (_04199_, _04198_, _03787_);
  or (_04200_, _03880_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_04201_, _03723_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_04202_, _04201_, _04200_);
  nand (_04203_, _04202_, _03788_);
  nand (_04204_, _04203_, _04199_);
  nand (_04205_, _04204_, _03650_);
  or (_04206_, _03880_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_04207_, _03723_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_04208_, _04207_, _04206_);
  nand (_04209_, _04208_, _03787_);
  or (_04210_, _03880_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_04211_, _03723_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_04212_, _04211_, _04210_);
  nand (_04213_, _04212_, _03788_);
  nand (_04214_, _04213_, _04209_);
  nand (_04215_, _04214_, _03865_);
  and (_04216_, _04215_, _03891_);
  and (_04217_, _04216_, _04205_);
  or (_04218_, _04217_, _04195_);
  and (_04219_, _04218_, _02471_);
  not (_04220_, _02471_);
  nor (_04221_, _04217_, _04195_);
  and (_04222_, _04221_, _04220_);
  nor (_04223_, _04222_, _04219_);
  nand (_04224_, _03723_, \oc8051_golden_model_1.IRAM[0] [0]);
  nand (_04225_, _03880_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_04226_, _04225_, _03788_);
  nand (_04227_, _04226_, _04224_);
  nand (_04228_, _03723_, \oc8051_golden_model_1.IRAM[2] [0]);
  nand (_04229_, _03880_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_04230_, _04229_, _03787_);
  nand (_04231_, _04230_, _04228_);
  nand (_04232_, _04231_, _04227_);
  nand (_04233_, _04232_, _03650_);
  nand (_04234_, _03723_, \oc8051_golden_model_1.IRAM[4] [0]);
  nand (_04235_, _03880_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_04236_, _04235_, _03788_);
  nand (_04237_, _04236_, _04234_);
  nand (_04238_, _03723_, \oc8051_golden_model_1.IRAM[6] [0]);
  nand (_04239_, _03880_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_04240_, _04239_, _03787_);
  nand (_04241_, _04240_, _04238_);
  nand (_04242_, _04241_, _04237_);
  nand (_04243_, _04242_, _03865_);
  and (_04244_, _04243_, _03864_);
  and (_04245_, _04244_, _04233_);
  nand (_04246_, _03723_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_04247_, _03723_, _03694_);
  and (_04248_, _04247_, _04246_);
  nand (_04249_, _04248_, _03787_);
  nand (_04250_, _03723_, _03683_);
  or (_04251_, _03723_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_04252_, _04251_, _04250_);
  nand (_04253_, _04252_, _03788_);
  nand (_04254_, _04253_, _04249_);
  nand (_04255_, _04254_, _03650_);
  nand (_04256_, _03723_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_04257_, _03723_, _03701_);
  and (_04258_, _04257_, _04256_);
  nand (_04259_, _04258_, _03787_);
  nand (_04260_, _03723_, _03706_);
  or (_04261_, _03723_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand (_04262_, _04261_, _04260_);
  nand (_04263_, _04262_, _03788_);
  nand (_04264_, _04263_, _04259_);
  nand (_04265_, _04264_, _03865_);
  and (_04266_, _04265_, _03891_);
  and (_04267_, _04266_, _04255_);
  or (_04268_, _04267_, _04245_);
  or (_04269_, _04268_, _02503_);
  nor (_04270_, _04267_, _04245_);
  or (_04271_, _04270_, _03452_);
  and (_04272_, _04271_, _04269_);
  and (_04273_, _04272_, _04223_);
  and (_04274_, _04273_, _04173_);
  and (_04275_, _04274_, _04073_);
  and (_04276_, _04275_, _02596_);
  nand (_04277_, _04274_, _04073_);
  and (_04278_, _04277_, _03102_);
  or (_04279_, _04278_, _04276_);
  or (_04280_, _04279_, _03107_);
  nand (_04281_, _03576_, \oc8051_golden_model_1.IRAM[0] [4]);
  or (_04282_, _03576_, _03965_);
  and (_04283_, _04282_, _03574_);
  nand (_04284_, _04283_, _04281_);
  or (_04285_, _03576_, _03970_);
  nand (_04286_, _03576_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_04287_, _04286_, _03582_);
  nand (_04288_, _04287_, _04285_);
  nand (_04289_, _04288_, _04284_);
  nand (_04290_, _04289_, _03385_);
  or (_04291_, _03576_, _03982_);
  nand (_04292_, _03576_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_04293_, _04292_, _03582_);
  nand (_04294_, _04293_, _04291_);
  nand (_04295_, _03576_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_04296_, _03576_, _03977_);
  and (_04297_, _04296_, _03574_);
  nand (_04298_, _04297_, _04295_);
  nand (_04299_, _04298_, _04294_);
  nand (_04300_, _04299_, _03589_);
  nand (_04301_, _04300_, _04290_);
  nand (_04302_, _04301_, _03286_);
  nand (_04303_, _03516_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_04304_, _03576_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_04305_, _04304_, _03582_);
  nand (_04306_, _04305_, _04303_);
  nand (_04307_, _03576_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand (_04308_, _03516_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_04309_, _04308_, _03574_);
  nand (_04310_, _04309_, _04307_);
  nand (_04311_, _04310_, _04306_);
  nand (_04312_, _04311_, _03385_);
  nand (_04313_, _03516_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_04314_, _03576_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_04315_, _04314_, _03582_);
  nand (_04316_, _04315_, _04313_);
  nand (_04317_, _03576_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand (_04318_, _03516_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_04319_, _04318_, _03574_);
  nand (_04320_, _04319_, _04317_);
  nand (_04321_, _04320_, _04316_);
  nand (_04322_, _04321_, _03589_);
  nand (_04323_, _04322_, _04312_);
  nand (_04324_, _04323_, _03609_);
  nand (_04325_, _04324_, _04302_);
  and (_04326_, _04325_, _02370_);
  nor (_04327_, _04325_, _02370_);
  nor (_04328_, _04327_, _04326_);
  nand (_04329_, _03576_, \oc8051_golden_model_1.IRAM[0] [6]);
  or (_04330_, _03576_, _03911_);
  and (_04331_, _04330_, _03574_);
  nand (_04332_, _04331_, _04329_);
  or (_04333_, _03576_, _03916_);
  nand (_04334_, _03576_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_04335_, _04334_, _03582_);
  nand (_04336_, _04335_, _04333_);
  nand (_04337_, _04336_, _04332_);
  nand (_04338_, _04337_, _03385_);
  or (_04339_, _03576_, _03928_);
  nand (_04340_, _03576_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_04341_, _04340_, _03582_);
  nand (_04342_, _04341_, _04339_);
  nand (_04343_, _03576_, \oc8051_golden_model_1.IRAM[4] [6]);
  or (_04344_, _03576_, _03923_);
  and (_04345_, _04344_, _03574_);
  nand (_04346_, _04345_, _04343_);
  nand (_04347_, _04346_, _04342_);
  nand (_04348_, _04347_, _03589_);
  nand (_04349_, _04348_, _04338_);
  nand (_04350_, _04349_, _03286_);
  nand (_04351_, _03516_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_04352_, _03576_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_04353_, _04352_, _03582_);
  nand (_04354_, _04353_, _04351_);
  nand (_04355_, _03576_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_04356_, _03516_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_04357_, _04356_, _03574_);
  nand (_04358_, _04357_, _04355_);
  nand (_04359_, _04358_, _04354_);
  nand (_04360_, _04359_, _03385_);
  nand (_04361_, _03516_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_04362_, _03576_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_04363_, _04362_, _03582_);
  nand (_04364_, _04363_, _04361_);
  nand (_04365_, _03576_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_04366_, _03516_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_04367_, _04366_, _03574_);
  nand (_04368_, _04367_, _04365_);
  nand (_04369_, _04368_, _04364_);
  nand (_04370_, _04369_, _03589_);
  nand (_04371_, _04370_, _04360_);
  nand (_04372_, _04371_, _03609_);
  nand (_04373_, _04372_, _04350_);
  and (_04374_, _04373_, _02295_);
  nor (_04375_, _04373_, _02295_);
  nor (_04376_, _04375_, _04374_);
  nor (_04377_, _04376_, _04328_);
  and (_04378_, _03644_, _02439_);
  nor (_04379_, _03644_, _02439_);
  nor (_04380_, _04379_, _04378_);
  not (_04381_, _04380_);
  nand (_04382_, _03576_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_04383_, _03576_, _04018_);
  and (_04384_, _04383_, _03574_);
  nand (_04385_, _04384_, _04382_);
  or (_04386_, _03576_, _04023_);
  nand (_04387_, _03576_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_04388_, _04387_, _03582_);
  nand (_04389_, _04388_, _04386_);
  nand (_04390_, _04389_, _04385_);
  nand (_04391_, _04390_, _03385_);
  or (_04392_, _03576_, _04035_);
  nand (_04393_, _03576_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_04394_, _04393_, _03582_);
  nand (_04395_, _04394_, _04392_);
  nand (_04396_, _03576_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_04397_, _03576_, _04030_);
  and (_04398_, _04397_, _03574_);
  nand (_04399_, _04398_, _04396_);
  nand (_04400_, _04399_, _04395_);
  nand (_04401_, _04400_, _03589_);
  nand (_04402_, _04401_, _04391_);
  nand (_04403_, _04402_, _03286_);
  nand (_04404_, _03516_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand (_04405_, _03576_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_04406_, _04405_, _03582_);
  nand (_04407_, _04406_, _04404_);
  nand (_04408_, _03576_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_04409_, _03576_, _04048_);
  and (_04410_, _04409_, _03574_);
  nand (_04411_, _04410_, _04408_);
  nand (_04412_, _04411_, _04407_);
  nand (_04413_, _04412_, _03385_);
  nand (_04414_, _03516_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_04415_, _03516_, _04054_);
  and (_04416_, _04415_, _03582_);
  nand (_04417_, _04416_, _04414_);
  nand (_04418_, _03576_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand (_04419_, _03516_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_04420_, _04419_, _03574_);
  nand (_04421_, _04420_, _04418_);
  nand (_04422_, _04421_, _04417_);
  nand (_04423_, _04422_, _03589_);
  nand (_04424_, _04423_, _04413_);
  nand (_04425_, _04424_, _03609_);
  nand (_04426_, _04425_, _04403_);
  or (_04427_, _04426_, _02222_);
  not (_04428_, _04427_);
  nor (_04429_, _03777_, _04220_);
  nor (_04430_, _04429_, _04428_);
  and (_04431_, _04430_, _04381_);
  and (_04432_, _04431_, _04377_);
  and (_04433_, _03859_, _02405_);
  nor (_04434_, _03859_, _02405_);
  nor (_04435_, _04434_, _04433_);
  nand (_04436_, _03576_, \oc8051_golden_model_1.IRAM[0] [5]);
  or (_04437_, _03576_, _03789_);
  and (_04438_, _04437_, _03574_);
  nand (_04439_, _04438_, _04436_);
  or (_04440_, _03576_, _03794_);
  nand (_04441_, _03576_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_04442_, _04441_, _03582_);
  nand (_04443_, _04442_, _04440_);
  nand (_04444_, _04443_, _04439_);
  nand (_04445_, _04444_, _03385_);
  or (_04446_, _03576_, _03872_);
  nand (_04447_, _03576_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_04448_, _04447_, _03582_);
  nand (_04449_, _04448_, _04446_);
  nand (_04450_, _03576_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_04451_, _03576_, _03867_);
  and (_04452_, _04451_, _03574_);
  nand (_04453_, _04452_, _04450_);
  nand (_04454_, _04453_, _04449_);
  nand (_04455_, _04454_, _03589_);
  nand (_04456_, _04455_, _04445_);
  nand (_04457_, _04456_, _03286_);
  nand (_04458_, _03516_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_04459_, _03576_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_04460_, _04459_, _03582_);
  nand (_04461_, _04460_, _04458_);
  nand (_04462_, _03576_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand (_04463_, _03516_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_04464_, _04463_, _03574_);
  nand (_04465_, _04464_, _04462_);
  nand (_04466_, _04465_, _04461_);
  nand (_04467_, _04466_, _03385_);
  nand (_04468_, _03516_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_04469_, _03576_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_04470_, _04469_, _03582_);
  nand (_04471_, _04470_, _04468_);
  nand (_04472_, _03576_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand (_04473_, _03516_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_04474_, _04473_, _03574_);
  nand (_04475_, _04474_, _04472_);
  nand (_04476_, _04475_, _04471_);
  nand (_04477_, _04476_, _03589_);
  nand (_04478_, _04477_, _04467_);
  nand (_04479_, _04478_, _03609_);
  nand (_04480_, _04479_, _04457_);
  and (_04481_, _04480_, _03299_);
  nor (_04482_, _04480_, _03299_);
  nor (_04483_, _04482_, _04481_);
  and (_04484_, _04483_, _04435_);
  nand (_04485_, _03715_, _03681_);
  and (_04486_, _04485_, _03452_);
  and (_04487_, _03716_, _02503_);
  nor (_04488_, _04487_, _04486_);
  and (_04489_, _03777_, _04220_);
  and (_04490_, _04426_, _02222_);
  nor (_04491_, _04490_, _04489_);
  and (_04492_, _04491_, _04488_);
  and (_04493_, _04492_, _04484_);
  and (_04494_, _04493_, _04432_);
  or (_04495_, _04494_, _03102_);
  nand (_04496_, _04494_, _03096_);
  and (_04497_, _04496_, _04495_);
  nor (_04498_, _01999_, _02021_);
  not (_04499_, _04498_);
  or (_04500_, _04499_, _04497_);
  and (_04501_, _03168_, _02555_);
  and (_04502_, _02672_, _03153_);
  not (_04503_, _03154_);
  not (_04504_, _01988_);
  and (_04505_, _02023_, _03394_);
  nor (_04506_, _04505_, _04504_);
  and (_04507_, _04506_, _04503_);
  or (_04508_, _04507_, _02555_);
  or (_04509_, _04504_, \oc8051_golden_model_1.PC [15]);
  nor (_04510_, _01997_, _01925_);
  or (_04511_, _04510_, _03154_);
  nor (_04512_, _01987_, _01925_);
  and (_04513_, _02022_, _01980_);
  and (_04514_, _04513_, _03394_);
  or (_04515_, _04514_, _04512_);
  or (_04516_, _04515_, _04511_);
  or (_04517_, _04516_, _04509_);
  and (_04518_, _04517_, _04508_);
  or (_04519_, _04518_, _04502_);
  and (_04520_, _02672_, _03394_);
  nor (_04521_, _04520_, _04512_);
  nor (_04522_, _04510_, _04502_);
  and (_04523_, _04522_, _04521_);
  or (_04524_, _04523_, _01914_);
  and (_04525_, _04524_, _01998_);
  and (_04526_, _04525_, _04519_);
  not (_04527_, _01998_);
  and (_04528_, _02555_, _04527_);
  or (_04529_, _04528_, _03406_);
  or (_04530_, _04529_, _04526_);
  and (_04531_, _04480_, _04325_);
  and (_04532_, _04426_, _04373_);
  and (_04533_, _04532_, _04531_);
  and (_04534_, _03777_, _03716_);
  and (_04535_, _03859_, _03644_);
  and (_04536_, _04535_, _04534_);
  nand (_04537_, _04536_, _04533_);
  and (_04538_, _04537_, _02562_);
  not (_04539_, _03406_);
  and (_04540_, _04536_, _04533_);
  and (_04541_, _04540_, _02555_);
  or (_04542_, _04541_, _04539_);
  or (_04543_, _04542_, _04538_);
  and (_04544_, _04543_, _04530_);
  and (_04545_, _02660_, _02674_);
  or (_04546_, _04545_, _04544_);
  and (_04547_, _04546_, _02662_);
  or (_04548_, _03859_, _02222_);
  and (_04549_, _02295_, _02222_);
  and (_04550_, _02370_, _02333_);
  and (_04551_, _04550_, _04549_);
  and (_04552_, _04551_, _03127_);
  nor (_04553_, _03452_, _02471_);
  and (_04554_, _04553_, _02439_);
  and (_04555_, _04554_, _04552_);
  and (_04556_, _04555_, \oc8051_golden_model_1.DPL [3]);
  not (_04557_, _04556_);
  nor (_04558_, _02503_, _02471_);
  and (_04559_, _04558_, _02439_);
  and (_04560_, _04559_, _04552_);
  and (_04561_, _04560_, \oc8051_golden_model_1.DPH [3]);
  and (_04562_, _03452_, _02471_);
  and (_04563_, _04562_, _02439_);
  and (_04564_, _04563_, _04552_);
  and (_04565_, _04564_, \oc8051_golden_model_1.SP [3]);
  nor (_04566_, _04565_, _04561_);
  and (_04567_, _04566_, _04557_);
  and (_04568_, _02503_, _02471_);
  and (_04569_, _02439_, _03127_);
  and (_04570_, _04569_, _04568_);
  and (_04571_, _03518_, _02333_);
  nor (_04572_, _02295_, _02204_);
  and (_04573_, _04572_, _04571_);
  and (_04574_, _04573_, _04570_);
  and (_04575_, _04574_, \oc8051_golden_model_1.PSW [3]);
  not (_04576_, _04575_);
  and (_04577_, _02439_, _02405_);
  and (_04578_, _04577_, _04568_);
  nor (_04579_, _02370_, _02333_);
  and (_04580_, _04579_, _04549_);
  and (_04581_, _04580_, _04578_);
  and (_04582_, _04581_, \oc8051_golden_model_1.IP [3]);
  and (_04583_, _02370_, _03299_);
  and (_04584_, _04583_, _04572_);
  and (_04585_, _04584_, _04570_);
  and (_04586_, _04585_, \oc8051_golden_model_1.ACC [3]);
  nor (_04587_, _04586_, _04582_);
  and (_04588_, _04587_, _04576_);
  and (_04589_, _04577_, _04558_);
  and (_04590_, _04589_, _04551_);
  and (_04591_, _04590_, \oc8051_golden_model_1.TL1 [3]);
  nor (_04592_, _02439_, _03127_);
  and (_04593_, _04592_, _04562_);
  and (_04594_, _04593_, _04551_);
  and (_04595_, _04594_, \oc8051_golden_model_1.TH1 [3]);
  nor (_04596_, _04595_, _04591_);
  and (_04597_, _04578_, _04551_);
  and (_04598_, _04597_, \oc8051_golden_model_1.TCON [3]);
  and (_04599_, _04579_, _04572_);
  and (_04600_, _04599_, _04570_);
  and (_04601_, _04600_, \oc8051_golden_model_1.B [3]);
  nor (_04602_, _04601_, _04598_);
  and (_04603_, _04602_, _04596_);
  and (_04604_, _04577_, _04562_);
  and (_04605_, _04604_, _04551_);
  and (_04606_, _04605_, \oc8051_golden_model_1.TMOD [3]);
  and (_04607_, _04577_, _04553_);
  and (_04608_, _04607_, _04551_);
  and (_04609_, _04608_, \oc8051_golden_model_1.TL0 [3]);
  nor (_04610_, _04609_, _04606_);
  and (_04611_, _04592_, _04568_);
  and (_04612_, _04611_, _04551_);
  and (_04613_, _04612_, \oc8051_golden_model_1.TH0 [3]);
  and (_04614_, _04571_, _04549_);
  and (_04615_, _04614_, _04578_);
  and (_04616_, _04615_, \oc8051_golden_model_1.SCON [3]);
  nor (_04617_, _04616_, _04613_);
  and (_04618_, _04617_, _04610_);
  and (_04619_, _04618_, _04603_);
  and (_04620_, _04619_, _04588_);
  and (_04621_, _04620_, _04567_);
  and (_04622_, _04558_, _04123_);
  and (_04623_, _04622_, _04552_);
  and (_04624_, _04623_, \oc8051_golden_model_1.PCON [3]);
  not (_04625_, _04624_);
  and (_04626_, _04614_, _04604_);
  and (_04627_, _04626_, \oc8051_golden_model_1.SBUF [3]);
  and (_04628_, _04583_, _04549_);
  and (_04629_, _04628_, _04578_);
  and (_04630_, _04629_, \oc8051_golden_model_1.IE [3]);
  nor (_04631_, _04630_, _04627_);
  and (_04632_, _04631_, _04625_);
  and (_04633_, _04568_, _02439_);
  and (_04634_, _04633_, _04552_);
  and (_04635_, _04634_, \oc8051_golden_model_1.P0 [3]);
  not (_04636_, _04635_);
  and (_04637_, _04614_, _04570_);
  and (_04638_, _04637_, \oc8051_golden_model_1.P1 [3]);
  not (_04639_, _04638_);
  and (_04640_, _04628_, _04570_);
  and (_04641_, _04640_, \oc8051_golden_model_1.P2 [3]);
  and (_04642_, _04580_, _04570_);
  and (_04643_, _04642_, \oc8051_golden_model_1.P3 [3]);
  nor (_04644_, _04643_, _04641_);
  and (_04645_, _04644_, _04639_);
  and (_04646_, _04645_, _04636_);
  and (_04647_, _04646_, _04632_);
  and (_04648_, _04647_, _04621_);
  and (_04649_, _04648_, _04548_);
  or (_04650_, _03644_, _02222_);
  and (_04651_, _04560_, \oc8051_golden_model_1.DPH [2]);
  not (_04652_, _04651_);
  and (_04653_, _04555_, \oc8051_golden_model_1.DPL [2]);
  and (_04654_, _04564_, \oc8051_golden_model_1.SP [2]);
  nor (_04655_, _04654_, _04653_);
  and (_04656_, _04655_, _04652_);
  and (_04657_, _04597_, \oc8051_golden_model_1.TCON [2]);
  not (_04658_, _04657_);
  and (_04659_, _04612_, \oc8051_golden_model_1.TH0 [2]);
  and (_04660_, _04615_, \oc8051_golden_model_1.SCON [2]);
  nor (_04661_, _04660_, _04659_);
  and (_04662_, _04661_, _04658_);
  and (_04663_, _04605_, \oc8051_golden_model_1.TMOD [2]);
  and (_04664_, _04594_, \oc8051_golden_model_1.TH1 [2]);
  nor (_04665_, _04664_, _04663_);
  and (_04666_, _04608_, \oc8051_golden_model_1.TL0 [2]);
  and (_04667_, _04590_, \oc8051_golden_model_1.TL1 [2]);
  nor (_04668_, _04667_, _04666_);
  and (_04669_, _04668_, _04665_);
  and (_04670_, _04669_, _04662_);
  and (_04671_, _04670_, _04656_);
  and (_04672_, _04574_, \oc8051_golden_model_1.PSW [2]);
  and (_04673_, _04585_, \oc8051_golden_model_1.ACC [2]);
  nor (_04674_, _04673_, _04672_);
  and (_04675_, _04581_, \oc8051_golden_model_1.IP [2]);
  and (_04676_, _04600_, \oc8051_golden_model_1.B [2]);
  nor (_04677_, _04676_, _04675_);
  and (_04678_, _04677_, _04674_);
  and (_04679_, _04623_, \oc8051_golden_model_1.PCON [2]);
  not (_04680_, _04679_);
  and (_04681_, _04626_, \oc8051_golden_model_1.SBUF [2]);
  and (_04682_, _04629_, \oc8051_golden_model_1.IE [2]);
  nor (_04683_, _04682_, _04681_);
  and (_04684_, _04683_, _04680_);
  and (_04685_, _04684_, _04678_);
  nand (_04686_, _04634_, \oc8051_golden_model_1.P0 [2]);
  and (_04687_, _04640_, \oc8051_golden_model_1.P2 [2]);
  and (_04688_, _04637_, \oc8051_golden_model_1.P1 [2]);
  and (_04689_, _04642_, \oc8051_golden_model_1.P3 [2]);
  or (_04690_, _04689_, _04688_);
  nor (_04691_, _04690_, _04687_);
  and (_04692_, _04691_, _04686_);
  and (_04693_, _04692_, _04685_);
  and (_04694_, _04693_, _04671_);
  and (_04695_, _04694_, _04650_);
  and (_04696_, _04695_, _04649_);
  or (_04697_, _04325_, _02222_);
  and (_04698_, _04615_, \oc8051_golden_model_1.SCON [4]);
  and (_04699_, _04626_, \oc8051_golden_model_1.SBUF [4]);
  nor (_04700_, _04699_, _04698_);
  and (_04701_, _04605_, \oc8051_golden_model_1.TMOD [4]);
  and (_04702_, _04629_, \oc8051_golden_model_1.IE [4]);
  nor (_04703_, _04702_, _04701_);
  and (_04704_, _04703_, _04700_);
  and (_04705_, _04564_, \oc8051_golden_model_1.SP [4]);
  not (_04706_, _04705_);
  and (_04707_, _04608_, \oc8051_golden_model_1.TL0 [4]);
  and (_04708_, _04594_, \oc8051_golden_model_1.TH1 [4]);
  nor (_04709_, _04708_, _04707_);
  and (_04710_, _04709_, _04706_);
  and (_04711_, _04560_, \oc8051_golden_model_1.DPH [4]);
  and (_04712_, _04555_, \oc8051_golden_model_1.DPL [4]);
  nor (_04713_, _04712_, _04711_);
  and (_04714_, _04713_, _04710_);
  and (_04715_, _04714_, _04704_);
  and (_04716_, _04581_, \oc8051_golden_model_1.IP [4]);
  and (_04717_, _04585_, \oc8051_golden_model_1.ACC [4]);
  nor (_04718_, _04717_, _04716_);
  and (_04719_, _04574_, \oc8051_golden_model_1.PSW [4]);
  and (_04720_, _04600_, \oc8051_golden_model_1.B [4]);
  nor (_04721_, _04720_, _04719_);
  and (_04722_, _04721_, _04718_);
  and (_04723_, _04597_, \oc8051_golden_model_1.TCON [4]);
  not (_04724_, _04723_);
  and (_04725_, _04612_, \oc8051_golden_model_1.TH0 [4]);
  and (_04726_, _04590_, \oc8051_golden_model_1.TL1 [4]);
  nor (_04727_, _04726_, _04725_);
  and (_04728_, _04727_, _04724_);
  and (_04729_, _04728_, _04722_);
  and (_04730_, _04637_, \oc8051_golden_model_1.P1 [4]);
  and (_04731_, _04640_, \oc8051_golden_model_1.P2 [4]);
  and (_04732_, _04642_, \oc8051_golden_model_1.P3 [4]);
  or (_04733_, _04732_, _04731_);
  nor (_04734_, _04733_, _04730_);
  and (_04735_, _04623_, \oc8051_golden_model_1.PCON [4]);
  and (_04736_, _04634_, \oc8051_golden_model_1.P0 [4]);
  nor (_04737_, _04736_, _04735_);
  and (_04738_, _04737_, _04734_);
  and (_04739_, _04738_, _04729_);
  and (_04740_, _04739_, _04715_);
  and (_04741_, _04740_, _04697_);
  or (_04742_, _04480_, _02222_);
  and (_04743_, _04560_, \oc8051_golden_model_1.DPH [5]);
  not (_04744_, _04743_);
  and (_04745_, _04555_, \oc8051_golden_model_1.DPL [5]);
  and (_04746_, _04564_, \oc8051_golden_model_1.SP [5]);
  nor (_04747_, _04746_, _04745_);
  and (_04748_, _04747_, _04744_);
  and (_04749_, _04597_, \oc8051_golden_model_1.TCON [5]);
  not (_04750_, _04749_);
  and (_04751_, _04612_, \oc8051_golden_model_1.TH0 [5]);
  and (_04752_, _04615_, \oc8051_golden_model_1.SCON [5]);
  nor (_04753_, _04752_, _04751_);
  and (_04754_, _04753_, _04750_);
  and (_04755_, _04605_, \oc8051_golden_model_1.TMOD [5]);
  and (_04756_, _04594_, \oc8051_golden_model_1.TH1 [5]);
  nor (_04757_, _04756_, _04755_);
  and (_04758_, _04608_, \oc8051_golden_model_1.TL0 [5]);
  and (_04759_, _04590_, \oc8051_golden_model_1.TL1 [5]);
  nor (_04760_, _04759_, _04758_);
  and (_04761_, _04760_, _04757_);
  and (_04762_, _04761_, _04754_);
  and (_04763_, _04762_, _04748_);
  and (_04764_, _04574_, \oc8051_golden_model_1.PSW [5]);
  and (_04765_, _04600_, \oc8051_golden_model_1.B [5]);
  nor (_04766_, _04765_, _04764_);
  and (_04767_, _04581_, \oc8051_golden_model_1.IP [5]);
  and (_04768_, _04585_, \oc8051_golden_model_1.ACC [5]);
  nor (_04769_, _04768_, _04767_);
  and (_04770_, _04769_, _04766_);
  and (_04771_, _04623_, \oc8051_golden_model_1.PCON [5]);
  not (_04772_, _04771_);
  and (_04773_, _04626_, \oc8051_golden_model_1.SBUF [5]);
  and (_04774_, _04629_, \oc8051_golden_model_1.IE [5]);
  nor (_04775_, _04774_, _04773_);
  and (_04776_, _04775_, _04772_);
  and (_04777_, _04776_, _04770_);
  nand (_04778_, _04634_, \oc8051_golden_model_1.P0 [5]);
  and (_04779_, _04640_, \oc8051_golden_model_1.P2 [5]);
  and (_04780_, _04637_, \oc8051_golden_model_1.P1 [5]);
  and (_04781_, _04642_, \oc8051_golden_model_1.P3 [5]);
  or (_04782_, _04781_, _04780_);
  nor (_04783_, _04782_, _04779_);
  and (_04784_, _04783_, _04778_);
  and (_04785_, _04784_, _04777_);
  and (_04786_, _04785_, _04763_);
  and (_04787_, _04786_, _04742_);
  and (_04788_, _04787_, _04741_);
  and (_04789_, _04788_, _04696_);
  or (_04790_, _03777_, _02222_);
  and (_04791_, _04608_, \oc8051_golden_model_1.TL0 [1]);
  and (_04792_, _04594_, \oc8051_golden_model_1.TH1 [1]);
  nor (_04793_, _04792_, _04791_);
  and (_04794_, _04605_, \oc8051_golden_model_1.TMOD [1]);
  and (_04795_, _04626_, \oc8051_golden_model_1.SBUF [1]);
  nor (_04796_, _04795_, _04794_);
  and (_04797_, _04796_, _04793_);
  and (_04798_, _04564_, \oc8051_golden_model_1.SP [1]);
  not (_04799_, _04798_);
  and (_04800_, _04615_, \oc8051_golden_model_1.SCON [1]);
  and (_04801_, _04629_, \oc8051_golden_model_1.IE [1]);
  nor (_04802_, _04801_, _04800_);
  and (_04803_, _04802_, _04799_);
  and (_04804_, _04555_, \oc8051_golden_model_1.DPL [1]);
  and (_04805_, _04560_, \oc8051_golden_model_1.DPH [1]);
  nor (_04806_, _04805_, _04804_);
  and (_04807_, _04806_, _04803_);
  and (_04808_, _04807_, _04797_);
  and (_04809_, _04581_, \oc8051_golden_model_1.IP [1]);
  and (_04810_, _04585_, \oc8051_golden_model_1.ACC [1]);
  nor (_04811_, _04810_, _04809_);
  and (_04812_, _04574_, \oc8051_golden_model_1.PSW [1]);
  and (_04813_, _04600_, \oc8051_golden_model_1.B [1]);
  nor (_04814_, _04813_, _04812_);
  and (_04815_, _04814_, _04811_);
  and (_04816_, _04612_, \oc8051_golden_model_1.TH0 [1]);
  not (_04817_, _04816_);
  and (_04818_, _04597_, \oc8051_golden_model_1.TCON [1]);
  and (_04819_, _04590_, \oc8051_golden_model_1.TL1 [1]);
  nor (_04820_, _04819_, _04818_);
  and (_04821_, _04820_, _04817_);
  and (_04822_, _04821_, _04815_);
  and (_04823_, _04642_, \oc8051_golden_model_1.P3 [1]);
  not (_04824_, _04823_);
  and (_04825_, _04637_, \oc8051_golden_model_1.P1 [1]);
  and (_04826_, _04640_, \oc8051_golden_model_1.P2 [1]);
  nor (_04827_, _04826_, _04825_);
  and (_04828_, _04827_, _04824_);
  and (_04829_, _04623_, \oc8051_golden_model_1.PCON [1]);
  and (_04830_, _04634_, \oc8051_golden_model_1.P0 [1]);
  nor (_04831_, _04830_, _04829_);
  and (_04832_, _04831_, _04828_);
  and (_04833_, _04832_, _04822_);
  and (_04834_, _04833_, _04808_);
  and (_04835_, _04834_, _04790_);
  or (_04836_, _04485_, _02222_);
  and (_04837_, _04623_, \oc8051_golden_model_1.PCON [0]);
  not (_04838_, _04837_);
  and (_04839_, _04629_, \oc8051_golden_model_1.IE [0]);
  and (_04840_, _04626_, \oc8051_golden_model_1.SBUF [0]);
  nor (_04841_, _04840_, _04839_);
  and (_04842_, _04841_, _04838_);
  and (_04843_, _04640_, \oc8051_golden_model_1.P2 [0]);
  and (_04844_, _04642_, \oc8051_golden_model_1.P3 [0]);
  nor (_04845_, _04844_, _04843_);
  and (_04846_, _04845_, _04842_);
  and (_04847_, _04581_, \oc8051_golden_model_1.IP [0]);
  and (_04848_, _04585_, \oc8051_golden_model_1.ACC [0]);
  nor (_04849_, _04848_, _04847_);
  and (_04850_, _04574_, \oc8051_golden_model_1.PSW [0]);
  and (_04851_, _04600_, \oc8051_golden_model_1.B [0]);
  nor (_04852_, _04851_, _04850_);
  and (_04853_, _04852_, _04849_);
  and (_04854_, _04612_, \oc8051_golden_model_1.TH0 [0]);
  and (_04855_, _04597_, \oc8051_golden_model_1.TCON [0]);
  nor (_04856_, _04855_, _04854_);
  and (_04857_, _04590_, \oc8051_golden_model_1.TL1 [0]);
  and (_04858_, _04637_, \oc8051_golden_model_1.P1 [0]);
  nor (_04859_, _04858_, _04857_);
  and (_04860_, _04859_, _04856_);
  and (_04861_, _04605_, \oc8051_golden_model_1.TMOD [0]);
  and (_04862_, _04608_, \oc8051_golden_model_1.TL0 [0]);
  nor (_04863_, _04862_, _04861_);
  and (_04864_, _04594_, \oc8051_golden_model_1.TH1 [0]);
  and (_04865_, _04615_, \oc8051_golden_model_1.SCON [0]);
  nor (_04866_, _04865_, _04864_);
  and (_04867_, _04866_, _04863_);
  and (_04868_, _04867_, _04860_);
  and (_04869_, _04868_, _04853_);
  and (_04870_, _04869_, _04846_);
  and (_04871_, _04570_, _04551_);
  and (_04872_, _04871_, \oc8051_golden_model_1.P0 [0]);
  not (_04873_, _04872_);
  and (_04874_, _04569_, _04558_);
  and (_04875_, _04874_, _04551_);
  and (_04876_, _04875_, \oc8051_golden_model_1.DPH [0]);
  not (_04877_, _04876_);
  and (_04878_, _04569_, _04562_);
  and (_04879_, _04878_, _04551_);
  and (_04880_, _04879_, \oc8051_golden_model_1.SP [0]);
  and (_04881_, _04569_, _04553_);
  and (_04882_, _04881_, _04551_);
  and (_04883_, _04882_, \oc8051_golden_model_1.DPL [0]);
  nor (_04884_, _04883_, _04880_);
  and (_04885_, _04884_, _04877_);
  and (_04886_, _04885_, _04873_);
  and (_04887_, _04886_, _04870_);
  nand (_04888_, _04887_, _04836_);
  and (_04889_, _04888_, _04835_);
  or (_04890_, _04373_, _02222_);
  and (_04891_, _04555_, \oc8051_golden_model_1.DPL [6]);
  not (_04892_, _04891_);
  and (_04893_, _04560_, \oc8051_golden_model_1.DPH [6]);
  and (_04894_, _04564_, \oc8051_golden_model_1.SP [6]);
  nor (_04895_, _04894_, _04893_);
  and (_04896_, _04895_, _04892_);
  and (_04897_, _04615_, \oc8051_golden_model_1.SCON [6]);
  not (_04898_, _04897_);
  and (_04899_, _04605_, \oc8051_golden_model_1.TMOD [6]);
  and (_04900_, _04594_, \oc8051_golden_model_1.TH1 [6]);
  nor (_04901_, _04900_, _04899_);
  and (_04902_, _04901_, _04898_);
  and (_04903_, _04612_, \oc8051_golden_model_1.TH0 [6]);
  and (_04904_, _04590_, \oc8051_golden_model_1.TL1 [6]);
  nor (_04905_, _04904_, _04903_);
  and (_04906_, _04597_, \oc8051_golden_model_1.TCON [6]);
  and (_04907_, _04608_, \oc8051_golden_model_1.TL0 [6]);
  nor (_04908_, _04907_, _04906_);
  and (_04909_, _04908_, _04905_);
  and (_04910_, _04909_, _04902_);
  and (_04911_, _04910_, _04896_);
  and (_04912_, _04623_, \oc8051_golden_model_1.PCON [6]);
  not (_04913_, _04912_);
  and (_04914_, _04626_, \oc8051_golden_model_1.SBUF [6]);
  and (_04915_, _04629_, \oc8051_golden_model_1.IE [6]);
  nor (_04916_, _04915_, _04914_);
  and (_04917_, _04916_, _04913_);
  and (_04918_, _04581_, \oc8051_golden_model_1.IP [6]);
  and (_04919_, _04600_, \oc8051_golden_model_1.B [6]);
  nor (_04920_, _04919_, _04918_);
  and (_04921_, _04574_, \oc8051_golden_model_1.PSW [6]);
  and (_04922_, _04585_, \oc8051_golden_model_1.ACC [6]);
  nor (_04923_, _04922_, _04921_);
  and (_04924_, _04923_, _04920_);
  and (_04925_, _04924_, _04917_);
  and (_04926_, _04634_, \oc8051_golden_model_1.P0 [6]);
  not (_04927_, _04926_);
  and (_04928_, _04640_, \oc8051_golden_model_1.P2 [6]);
  not (_04929_, _04928_);
  and (_04930_, _04637_, \oc8051_golden_model_1.P1 [6]);
  and (_04931_, _04642_, \oc8051_golden_model_1.P3 [6]);
  nor (_04932_, _04931_, _04930_);
  and (_04933_, _04932_, _04929_);
  and (_04934_, _04933_, _04927_);
  and (_04935_, _04934_, _04925_);
  and (_04936_, _04935_, _04911_);
  and (_04937_, _04936_, _04890_);
  and (_04938_, _04581_, \oc8051_golden_model_1.IP [7]);
  not (_04939_, _04938_);
  and (_04940_, _04574_, \oc8051_golden_model_1.PSW [7]);
  not (_04941_, _04940_);
  and (_04942_, _04600_, \oc8051_golden_model_1.B [7]);
  and (_04943_, _04585_, \oc8051_golden_model_1.ACC [7]);
  nor (_04944_, _04943_, _04942_);
  and (_04945_, _04944_, _04941_);
  and (_04946_, _04945_, _04939_);
  and (_04947_, _04871_, \oc8051_golden_model_1.P0 [7]);
  and (_04948_, _04875_, \oc8051_golden_model_1.DPH [7]);
  nor (_04949_, _04948_, _04947_);
  and (_04950_, _04626_, \oc8051_golden_model_1.SBUF [7]);
  and (_04951_, _04629_, \oc8051_golden_model_1.IE [7]);
  nor (_04952_, _04951_, _04950_);
  and (_04953_, _04642_, \oc8051_golden_model_1.P3 [7]);
  not (_04954_, _04953_);
  and (_04955_, _04640_, \oc8051_golden_model_1.P2 [7]);
  and (_04956_, _04623_, \oc8051_golden_model_1.PCON [7]);
  nor (_04957_, _04956_, _04955_);
  and (_04958_, _04957_, _04954_);
  and (_04959_, _04958_, _04952_);
  and (_04960_, _04879_, \oc8051_golden_model_1.SP [7]);
  and (_04961_, _04882_, \oc8051_golden_model_1.DPL [7]);
  nor (_04962_, _04961_, _04960_);
  and (_04963_, _04597_, \oc8051_golden_model_1.TCON [7]);
  and (_04964_, _04612_, \oc8051_golden_model_1.TH0 [7]);
  nor (_04965_, _04964_, _04963_);
  and (_04966_, _04590_, \oc8051_golden_model_1.TL1 [7]);
  and (_04967_, _04637_, \oc8051_golden_model_1.P1 [7]);
  nor (_04968_, _04967_, _04966_);
  and (_04969_, _04968_, _04965_);
  and (_04970_, _04594_, \oc8051_golden_model_1.TH1 [7]);
  and (_04971_, _04615_, \oc8051_golden_model_1.SCON [7]);
  nor (_04972_, _04971_, _04970_);
  and (_04973_, _04605_, \oc8051_golden_model_1.TMOD [7]);
  and (_04974_, _04608_, \oc8051_golden_model_1.TL0 [7]);
  nor (_04975_, _04974_, _04973_);
  and (_04976_, _04975_, _04972_);
  and (_04977_, _04976_, _04969_);
  and (_04978_, _04977_, _04962_);
  and (_04979_, _04978_, _04959_);
  and (_04980_, _04979_, _04949_);
  and (_04981_, _04980_, _04946_);
  and (_04982_, _04981_, _04427_);
  and (_04983_, _04982_, _04937_);
  and (_04984_, _04983_, _04889_);
  and (_04985_, _04984_, _04789_);
  or (_04986_, _04985_, _03102_);
  nand (_04987_, _04984_, _04789_);
  or (_04988_, _04987_, _02596_);
  and (_04989_, _04988_, _02661_);
  and (_04990_, _04989_, _04986_);
  nor (_04991_, _02672_, _02572_);
  nor (_04992_, _04991_, _01994_);
  or (_04993_, _04992_, _04990_);
  or (_04994_, _04993_, _04547_);
  and (_04995_, _03163_, _01995_);
  nor (_04996_, _04992_, _04545_);
  or (_04997_, _04996_, _01914_);
  and (_04998_, _04997_, _04995_);
  and (_04999_, _04998_, _04994_);
  nor (_05000_, _01989_, _01925_);
  nor (_05001_, _04995_, _02556_);
  or (_05002_, _05001_, _05000_);
  or (_05003_, _05002_, _04999_);
  not (_05004_, _05000_);
  or (_05005_, _05004_, _01914_);
  and (_05006_, _05005_, _03179_);
  and (_05007_, _05006_, _05003_);
  or (_05008_, _05007_, _04501_);
  nor (_05009_, _04991_, _01989_);
  not (_05010_, _05009_);
  and (_05011_, _05010_, _05008_);
  and (_05012_, _05009_, _01914_);
  and (_05013_, _03428_, _01990_);
  not (_05014_, _05013_);
  or (_05015_, _05014_, _05012_);
  or (_05016_, _05015_, _05011_);
  or (_05017_, _05013_, _02555_);
  and (_05018_, _05017_, _05016_);
  or (_05019_, _05018_, _04498_);
  and (_05020_, _05019_, _04500_);
  or (_05021_, _05020_, _02675_);
  and (_05022_, _05021_, _04280_);
  or (_05023_, _05022_, _02664_);
  not (_05024_, _02673_);
  and (_05025_, _04640_, \oc8051_golden_model_1.P2INREG [1]);
  not (_05026_, _05025_);
  and (_05027_, _04637_, \oc8051_golden_model_1.P1INREG [1]);
  and (_05028_, _04642_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_05029_, _05028_, _05027_);
  and (_05030_, _05029_, _05026_);
  and (_05031_, _04634_, \oc8051_golden_model_1.P0INREG [1]);
  nor (_05032_, _05031_, _04829_);
  and (_05033_, _05032_, _05030_);
  and (_05034_, _05033_, _04822_);
  and (_05035_, _05034_, _04808_);
  and (_05036_, _05035_, _04790_);
  nor (_05037_, _05036_, \oc8051_golden_model_1.ACC [1]);
  and (_05038_, _05036_, \oc8051_golden_model_1.ACC [1]);
  nor (_05039_, _05038_, _05037_);
  not (_05040_, _04963_);
  not (_05041_, _04948_);
  and (_05042_, _04962_, _05041_);
  and (_05043_, _05042_, _05040_);
  nor (_05044_, _04964_, _04966_);
  and (_05045_, _05044_, _04975_);
  and (_05046_, _04640_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05047_, _04642_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05048_, _05047_, _05046_);
  and (_05049_, _04637_, \oc8051_golden_model_1.P1INREG [7]);
  and (_05050_, _04871_, \oc8051_golden_model_1.P0INREG [7]);
  nor (_05051_, _05050_, _05049_);
  and (_05052_, _05051_, _05048_);
  and (_05053_, _05052_, _05045_);
  and (_05054_, _05053_, _05043_);
  not (_05055_, _04956_);
  and (_05056_, _05055_, _04972_);
  and (_05057_, _05056_, _04952_);
  and (_05058_, _05057_, _04946_);
  and (_05059_, _05058_, _05054_);
  and (_05060_, _05059_, _04427_);
  nor (_05061_, _05060_, \oc8051_golden_model_1.ACC [7]);
  and (_05062_, _05060_, \oc8051_golden_model_1.ACC [7]);
  nor (_05063_, _05062_, _05061_);
  and (_05064_, _05063_, _05039_);
  and (_05065_, _04640_, \oc8051_golden_model_1.P2INREG [2]);
  and (_05066_, _04642_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_05067_, _05066_, _05065_);
  and (_05068_, _04637_, \oc8051_golden_model_1.P1INREG [2]);
  and (_05069_, _04871_, \oc8051_golden_model_1.P0INREG [2]);
  nor (_05070_, _05069_, _05068_);
  and (_05071_, _05070_, _05067_);
  and (_05072_, _05071_, _04685_);
  and (_05073_, _05072_, _04671_);
  and (_05074_, _05073_, _04650_);
  nor (_05075_, _05074_, \oc8051_golden_model_1.ACC [2]);
  and (_05076_, _05074_, \oc8051_golden_model_1.ACC [2]);
  nor (_05077_, _05076_, _05075_);
  and (_05078_, _04640_, \oc8051_golden_model_1.P2INREG [6]);
  and (_05079_, _04642_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_05080_, _05079_, _05078_);
  and (_05081_, _04637_, \oc8051_golden_model_1.P1INREG [6]);
  and (_05082_, _04871_, \oc8051_golden_model_1.P0INREG [6]);
  nor (_05083_, _05082_, _05081_);
  and (_05084_, _05083_, _05080_);
  and (_05085_, _05084_, _04925_);
  and (_05086_, _05085_, _04911_);
  and (_05087_, _05086_, _04890_);
  nor (_05088_, _05087_, \oc8051_golden_model_1.ACC [6]);
  and (_05089_, _05087_, \oc8051_golden_model_1.ACC [6]);
  nor (_05090_, _05089_, _05088_);
  and (_05091_, _05090_, _05077_);
  and (_05092_, _05091_, _05064_);
  not (_05093_, _04855_);
  and (_05094_, _04885_, _05093_);
  and (_05095_, _04640_, \oc8051_golden_model_1.P2INREG [0]);
  and (_05096_, _04642_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_05097_, _05096_, _05095_);
  and (_05098_, _04637_, \oc8051_golden_model_1.P1INREG [0]);
  and (_05099_, _04871_, \oc8051_golden_model_1.P0INREG [0]);
  nor (_05100_, _05099_, _05098_);
  and (_05101_, _05100_, _05097_);
  nor (_05102_, _04857_, _04854_);
  and (_05103_, _05102_, _04863_);
  and (_05104_, _05103_, _05101_);
  and (_05105_, _05104_, _05094_);
  and (_05106_, _04866_, _04842_);
  and (_05107_, _05106_, _04853_);
  and (_05108_, _05107_, _05105_);
  and (_05109_, _05108_, _04836_);
  nor (_05110_, _05109_, \oc8051_golden_model_1.ACC [0]);
  and (_05111_, _05109_, \oc8051_golden_model_1.ACC [0]);
  nor (_05112_, _05111_, _05110_);
  and (_05113_, _04642_, \oc8051_golden_model_1.P3INREG [4]);
  not (_05114_, _05113_);
  and (_05115_, _04637_, \oc8051_golden_model_1.P1INREG [4]);
  and (_05116_, _04640_, \oc8051_golden_model_1.P2INREG [4]);
  nor (_05117_, _05116_, _05115_);
  and (_05118_, _05117_, _05114_);
  and (_05119_, _04634_, \oc8051_golden_model_1.P0INREG [4]);
  nor (_05120_, _05119_, _04735_);
  and (_05121_, _05120_, _05118_);
  and (_05122_, _05121_, _04729_);
  and (_05123_, _05122_, _04715_);
  and (_05124_, _05123_, _04697_);
  nor (_05125_, _05124_, \oc8051_golden_model_1.ACC [4]);
  and (_05126_, _05124_, \oc8051_golden_model_1.ACC [4]);
  nor (_05127_, _05126_, _05125_);
  and (_05128_, _05127_, _05112_);
  and (_05129_, _04640_, \oc8051_golden_model_1.P2INREG [3]);
  and (_05130_, _04642_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_05131_, _05130_, _05129_);
  and (_05132_, _04637_, \oc8051_golden_model_1.P1INREG [3]);
  and (_05133_, _04871_, \oc8051_golden_model_1.P0INREG [3]);
  nor (_05134_, _05133_, _05132_);
  and (_05135_, _05134_, _05131_);
  and (_05136_, _05135_, _04632_);
  and (_05137_, _05136_, _04621_);
  and (_05138_, _05137_, _04548_);
  nor (_05139_, _05138_, \oc8051_golden_model_1.ACC [3]);
  and (_05140_, _05138_, \oc8051_golden_model_1.ACC [3]);
  nor (_05141_, _05140_, _05139_);
  and (_05142_, _04640_, \oc8051_golden_model_1.P2INREG [5]);
  and (_05143_, _04642_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_05144_, _05143_, _05142_);
  and (_05145_, _04637_, \oc8051_golden_model_1.P1INREG [5]);
  and (_05146_, _04871_, \oc8051_golden_model_1.P0INREG [5]);
  nor (_05147_, _05146_, _05145_);
  and (_05148_, _05147_, _05144_);
  and (_05149_, _05148_, _04777_);
  and (_05150_, _05149_, _04763_);
  and (_05151_, _05150_, _04742_);
  nor (_05152_, _05151_, \oc8051_golden_model_1.ACC [5]);
  and (_05153_, _05151_, \oc8051_golden_model_1.ACC [5]);
  nor (_05154_, _05153_, _05152_);
  and (_05155_, _05154_, _05141_);
  and (_05156_, _05155_, _05128_);
  and (_05157_, _05156_, _05092_);
  not (_05158_, _05157_);
  and (_05159_, _05158_, _03102_);
  and (_05160_, _05157_, _02596_);
  or (_05161_, _05160_, _03387_);
  or (_05162_, _05161_, _05159_);
  and (_05163_, _05162_, _05024_);
  and (_05164_, _05163_, _05023_);
  or (_05165_, _05164_, _03106_);
  and (_05166_, _05165_, _02599_);
  nand (_05167_, _02598_, _01914_);
  not (_05168_, _03144_);
  nor (_05169_, _01920_, _02636_);
  nor (_05170_, _05169_, _01992_);
  not (_05171_, _05170_);
  and (_05172_, _03118_, _01917_);
  and (_05173_, _05172_, _01981_);
  not (_05174_, _05173_);
  nor (_05175_, _03143_, _03119_);
  and (_05176_, _05175_, _05174_);
  and (_05177_, _05176_, _05171_);
  and (_05178_, _05177_, _02000_);
  and (_05179_, _05178_, _05168_);
  nand (_05180_, _05179_, _05167_);
  or (_05181_, _05180_, _05166_);
  or (_05182_, _05179_, _02555_);
  not (_05183_, _02023_);
  and (_05184_, _04991_, _05183_);
  nor (_05185_, _05184_, _01992_);
  not (_05186_, _05185_);
  and (_05187_, _05186_, _05182_);
  and (_05188_, _05187_, _05181_);
  and (_05189_, _05185_, _01914_);
  and (_05190_, _03207_, _01993_);
  not (_05191_, _05190_);
  or (_05192_, _05191_, _05189_);
  or (_05193_, _05192_, _05188_);
  nor (_05194_, _01984_, _01925_);
  not (_05195_, _05194_);
  or (_05196_, _05190_, _02555_);
  and (_05197_, _05196_, _05195_);
  and (_05198_, _05197_, _05193_);
  and (_05199_, _04513_, _01983_);
  and (_05200_, _05194_, _01914_);
  or (_05201_, _05200_, _05199_);
  or (_05202_, _05201_, _05198_);
  not (_05203_, _05199_);
  or (_05204_, _05203_, _02555_);
  and (_05205_, _05204_, _01985_);
  and (_05206_, _05205_, _05202_);
  and (_05207_, _02047_, _01914_);
  nor (_05208_, _03140_, _02025_);
  not (_05209_, _05208_);
  or (_05210_, _05209_, _05207_);
  or (_05211_, _05210_, _05206_);
  not (_05212_, _02670_);
  or (_05213_, _05208_, _02555_);
  and (_05214_, _05213_, _05212_);
  and (_05215_, _05214_, _05211_);
  and (_05216_, _02670_, _02596_);
  nor (_05217_, _02029_, _01925_);
  or (_05218_, _05217_, _05216_);
  or (_05219_, _05218_, _05215_);
  not (_05220_, _05217_);
  or (_05221_, _05220_, _02555_);
  and (_05222_, _05221_, _03139_);
  and (_05223_, _05222_, _05219_);
  or (_05224_, _05223_, _02597_);
  nor (_05225_, _04991_, _02029_);
  not (_05226_, _05225_);
  and (_05227_, _05226_, _05224_);
  nor (_05228_, _03135_, _01960_);
  not (_05229_, _05228_);
  and (_05230_, _05225_, _01914_);
  or (_05231_, _05230_, _05229_);
  or (_05232_, _05231_, _05227_);
  and (_05233_, _02566_, _01959_);
  not (_05234_, _05233_);
  or (_05235_, _05228_, _02555_);
  and (_05236_, _05235_, _05234_);
  and (_05237_, _05236_, _05232_);
  and (_05238_, _05233_, _02562_);
  or (_05239_, _05238_, _02577_);
  or (_05240_, _05239_, _05237_);
  and (_05241_, _05240_, _02578_);
  or (_05242_, _05241_, _02575_);
  and (_05243_, _02672_, _01966_);
  not (_05244_, _05243_);
  not (_05245_, _02575_);
  or (_05246_, _02596_, _05245_);
  and (_05247_, _05246_, _05244_);
  and (_05248_, _05247_, _05242_);
  and (_05249_, _05243_, _02555_);
  or (_05250_, _05249_, _05248_);
  and (_05251_, _05250_, _02574_);
  nor (_05252_, _03134_, _01967_);
  not (_05253_, _05252_);
  not (_05254_, \oc8051_golden_model_1.DPH [0]);
  and (_05255_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_05256_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and (_05257_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_05258_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_05259_, _05258_, _05257_);
  not (_05260_, _05259_);
  and (_05261_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_05262_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_05263_, _05262_, _05261_);
  not (_05264_, _05263_);
  and (_05265_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_05266_, _02116_, _02112_);
  nor (_05267_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_05268_, _05267_, _05265_);
  not (_05269_, _05268_);
  nor (_05270_, _05269_, _05266_);
  nor (_05271_, _05270_, _05265_);
  nor (_05272_, _05271_, _05264_);
  nor (_05273_, _05272_, _05261_);
  nor (_05274_, _05273_, _05260_);
  nor (_05275_, _05274_, _05257_);
  nor (_05276_, _05275_, _05256_);
  nor (_05277_, _05276_, _05255_);
  nor (_05278_, _05277_, _05254_);
  and (_05279_, _05278_, \oc8051_golden_model_1.DPH [1]);
  and (_05280_, _05279_, \oc8051_golden_model_1.DPH [2]);
  and (_05281_, _05280_, \oc8051_golden_model_1.DPH [3]);
  and (_05282_, _05281_, \oc8051_golden_model_1.DPH [4]);
  and (_05283_, _05282_, \oc8051_golden_model_1.DPH [5]);
  and (_05284_, _05283_, \oc8051_golden_model_1.DPH [6]);
  nand (_05285_, _05284_, \oc8051_golden_model_1.DPH [7]);
  or (_05286_, _05284_, \oc8051_golden_model_1.DPH [7]);
  and (_05287_, _05286_, _02573_);
  and (_05288_, _05287_, _05285_);
  or (_05289_, _05288_, _05253_);
  or (_05290_, _05289_, _05251_);
  not (_05291_, _02567_);
  or (_05292_, _05252_, _02555_);
  and (_05293_, _05292_, _05291_);
  and (_05294_, _05293_, _05290_);
  or (_05295_, _05294_, _02571_);
  not (_05296_, _01973_);
  nor (_05297_, _05296_, _01925_);
  not (_05298_, _05297_);
  and (_05299_, _05298_, _05295_);
  and (_05300_, _05297_, _01914_);
  and (_05302_, _04513_, _01973_);
  or (_05303_, _05302_, _05300_);
  or (_05304_, _05303_, _05299_);
  not (_05305_, _02656_);
  not (_05306_, _05302_);
  or (_05307_, _05306_, _02555_);
  and (_05308_, _05307_, _05305_);
  and (_05309_, _05308_, _05304_);
  and (_05310_, _02656_, _02596_);
  nor (_05311_, _03251_, _01974_);
  not (_05312_, _05311_);
  or (_05313_, _05312_, _05310_);
  or (_05314_, _05313_, _05309_);
  and (_05315_, _02566_, _01973_);
  not (_05316_, _05315_);
  or (_05317_, _05311_, _02555_);
  and (_05318_, _05317_, _05316_);
  and (_05319_, _05318_, _05314_);
  or (_05320_, _02562_, _02568_);
  or (_05321_, _02555_, _01953_);
  and (_05322_, _05321_, _05315_);
  and (_05323_, _05322_, _05320_);
  or (_05324_, _05323_, _05319_);
  nor (_05325_, _03359_, _01925_);
  not (_05326_, _05325_);
  and (_05327_, _05326_, _05324_);
  and (_05328_, _05325_, _01914_);
  and (_05329_, _04513_, _01964_);
  or (_05330_, _05329_, _05328_);
  or (_05331_, _05330_, _05327_);
  not (_05332_, _02669_);
  not (_05333_, _05329_);
  or (_05334_, _05333_, _02555_);
  and (_05335_, _05334_, _05332_);
  and (_05336_, _05335_, _05331_);
  and (_05337_, _02669_, _02596_);
  nor (_05338_, _03243_, _01965_);
  not (_05339_, _05338_);
  or (_05340_, _05339_, _05337_);
  or (_05341_, _05340_, _05336_);
  and (_05342_, _02566_, _01964_);
  not (_05343_, _05342_);
  or (_05344_, _05338_, _02555_);
  and (_05345_, _05344_, _05343_);
  and (_05346_, _05345_, _05341_);
  or (_05347_, _02562_, \oc8051_golden_model_1.PSW [7]);
  not (_05348_, \oc8051_golden_model_1.PSW [7]);
  or (_05349_, _02555_, _05348_);
  and (_05350_, _05349_, _05342_);
  and (_05351_, _05350_, _05347_);
  or (_05352_, _05351_, _01944_);
  or (_05353_, _05352_, _05346_);
  and (_05354_, _05353_, _01946_);
  and (_05355_, _04513_, _01942_);
  or (_05356_, _05355_, _05354_);
  not (_05357_, _02654_);
  not (_05358_, _05355_);
  or (_05359_, _05358_, _02555_);
  and (_05360_, _05359_, _05357_);
  and (_05361_, _05360_, _05356_);
  and (_05362_, _02654_, _02596_);
  nor (_05363_, _03239_, _01957_);
  not (_05364_, _05363_);
  or (_05365_, _05364_, _05362_);
  or (_05366_, _05365_, _05361_);
  and (_05367_, _02566_, _01942_);
  not (_05368_, _05367_);
  or (_05369_, _05363_, _02555_);
  and (_05370_, _05369_, _05368_);
  and (_05371_, _05370_, _05366_);
  or (_05372_, _02562_, _05348_);
  or (_05373_, _02555_, \oc8051_golden_model_1.PSW [7]);
  and (_05374_, _05373_, _05367_);
  and (_05375_, _05374_, _05372_);
  or (_05376_, _05375_, _05371_);
  and (_05377_, _02674_, _03399_);
  or (_05378_, _05377_, _02633_);
  not (_05379_, _05378_);
  and (_05380_, _03354_, _01918_);
  not (_05381_, _02640_);
  and (_05382_, _05381_, _05380_);
  and (_05383_, _05382_, _05379_);
  nor (_05384_, _05383_, _03482_);
  not (_05385_, _05384_);
  and (_05386_, _03395_, _01935_);
  and (_05387_, _01935_, _03339_);
  nor (_05388_, _05387_, _05386_);
  and (_05389_, _05388_, _05385_);
  and (_05390_, _05389_, _05376_);
  not (_05391_, _05389_);
  and (_05392_, _05391_, _01914_);
  and (_05393_, _04513_, _01935_);
  or (_05394_, _05393_, _05392_);
  or (_05395_, _05394_, _05390_);
  and (_05396_, _02572_, _01935_);
  not (_05397_, _05396_);
  not (_05398_, _05393_);
  or (_05399_, _05398_, _02555_);
  and (_05400_, _05399_, _05397_);
  and (_05401_, _05400_, _05395_);
  and (_05402_, _05396_, _01914_);
  or (_05403_, _05402_, _03109_);
  or (_05404_, _05403_, _05401_);
  nand (_05405_, _04426_, _03109_);
  and (_05406_, _05405_, _05404_);
  or (_05407_, _05406_, _01936_);
  not (_05408_, _01936_);
  or (_05409_, _02555_, _05408_);
  and (_05410_, _05409_, _03267_);
  and (_05411_, _05410_, _05407_);
  not (_05412_, _01930_);
  not (_05413_, _04554_);
  nor (_05414_, _03521_, _03391_);
  nor (_05415_, _03303_, _03133_);
  and (_05416_, _05415_, _05414_);
  and (_05417_, _04573_, _05416_);
  and (_05418_, _05417_, \oc8051_golden_model_1.PSW [2]);
  and (_05419_, _04599_, _05416_);
  and (_05420_, _05419_, \oc8051_golden_model_1.B [2]);
  nor (_05421_, _05420_, _05418_);
  not (_05422_, _03303_);
  and (_05423_, _05414_, _03133_);
  and (_05424_, _05423_, _05422_);
  and (_05425_, _05424_, _04580_);
  and (_05426_, _05425_, \oc8051_golden_model_1.IP [2]);
  and (_05427_, _04584_, _05416_);
  and (_05428_, _05427_, \oc8051_golden_model_1.ACC [2]);
  nor (_05429_, _05428_, _05426_);
  and (_05430_, _05429_, _05421_);
  and (_05431_, _05424_, _04614_);
  and (_05432_, _05431_, \oc8051_golden_model_1.SCON [2]);
  and (_05433_, _05424_, _04628_);
  and (_05434_, _05433_, \oc8051_golden_model_1.IE [2]);
  nor (_05435_, _05434_, _05432_);
  and (_05436_, _04628_, _05416_);
  and (_05437_, _05436_, \oc8051_golden_model_1.P2INREG [2]);
  not (_05438_, _05437_);
  and (_05439_, _04552_, \oc8051_golden_model_1.P0INREG [2]);
  and (_05440_, _05423_, _04551_);
  and (_05441_, _05440_, \oc8051_golden_model_1.TCON [2]);
  nor (_05442_, _05441_, _05439_);
  and (_05443_, _05442_, _05438_);
  and (_05444_, _04614_, _05416_);
  and (_05445_, _05444_, \oc8051_golden_model_1.P1INREG [2]);
  and (_05446_, _04580_, _05416_);
  and (_05447_, _05446_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_05448_, _05447_, _05445_);
  and (_05449_, _05448_, _05443_);
  and (_05450_, _05449_, _05435_);
  and (_05451_, _05450_, _05430_);
  and (_05452_, _05451_, _04650_);
  nor (_05453_, _05452_, _05413_);
  not (_05454_, _04563_);
  and (_05455_, _05425_, \oc8051_golden_model_1.IP [1]);
  and (_05456_, _05419_, \oc8051_golden_model_1.B [1]);
  nor (_05457_, _05456_, _05455_);
  and (_05458_, _05417_, \oc8051_golden_model_1.PSW [1]);
  and (_05459_, _05427_, \oc8051_golden_model_1.ACC [1]);
  nor (_05460_, _05459_, _05458_);
  and (_05461_, _05460_, _05457_);
  and (_05462_, _05431_, \oc8051_golden_model_1.SCON [1]);
  and (_05463_, _05433_, \oc8051_golden_model_1.IE [1]);
  nor (_05464_, _05463_, _05462_);
  and (_05465_, _05436_, \oc8051_golden_model_1.P2INREG [1]);
  and (_05466_, _05446_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_05467_, _05466_, _05465_);
  and (_05468_, _05444_, \oc8051_golden_model_1.P1INREG [1]);
  not (_05469_, _05468_);
  and (_05470_, _04552_, \oc8051_golden_model_1.P0INREG [1]);
  and (_05471_, _05440_, \oc8051_golden_model_1.TCON [1]);
  nor (_05472_, _05471_, _05470_);
  and (_05473_, _05472_, _05469_);
  and (_05474_, _05473_, _05467_);
  and (_05475_, _05474_, _05464_);
  and (_05476_, _05475_, _05461_);
  and (_05477_, _05476_, _04790_);
  nor (_05478_, _05477_, _05454_);
  nor (_05479_, _05478_, _05453_);
  and (_05480_, _05425_, \oc8051_golden_model_1.IP [4]);
  and (_05481_, _05427_, \oc8051_golden_model_1.ACC [4]);
  nor (_05482_, _05481_, _05480_);
  and (_05483_, _05433_, \oc8051_golden_model_1.IE [4]);
  and (_05484_, _05417_, \oc8051_golden_model_1.PSW [4]);
  nor (_05485_, _05484_, _05483_);
  and (_05486_, _05431_, \oc8051_golden_model_1.SCON [4]);
  and (_05487_, _05419_, \oc8051_golden_model_1.B [4]);
  nor (_05488_, _05487_, _05486_);
  and (_05489_, _05488_, _05485_);
  and (_05490_, _05489_, _05482_);
  and (_05491_, _05436_, \oc8051_golden_model_1.P2INREG [4]);
  and (_05492_, _05446_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_05493_, _05492_, _05491_);
  and (_05494_, _05444_, \oc8051_golden_model_1.P1INREG [4]);
  not (_05495_, _05494_);
  and (_05496_, _04552_, \oc8051_golden_model_1.P0INREG [4]);
  and (_05497_, _05440_, \oc8051_golden_model_1.TCON [4]);
  nor (_05498_, _05497_, _05496_);
  and (_05499_, _05498_, _05495_);
  and (_05500_, _05499_, _05493_);
  and (_05501_, _05500_, _05490_);
  and (_05502_, _05501_, _04697_);
  and (_05503_, _04568_, _04123_);
  not (_05504_, _05503_);
  nor (_05505_, _05504_, _05502_);
  not (_05506_, _04622_);
  and (_05507_, _05417_, \oc8051_golden_model_1.PSW [7]);
  and (_05508_, _05419_, \oc8051_golden_model_1.B [7]);
  nor (_05509_, _05508_, _05507_);
  and (_05510_, _05425_, \oc8051_golden_model_1.IP [7]);
  and (_05511_, _05427_, \oc8051_golden_model_1.ACC [7]);
  nor (_05512_, _05511_, _05510_);
  and (_05513_, _05512_, _05509_);
  and (_05514_, _05431_, \oc8051_golden_model_1.SCON [7]);
  and (_05515_, _05433_, \oc8051_golden_model_1.IE [7]);
  nor (_05516_, _05515_, _05514_);
  and (_05517_, _05436_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05518_, _05446_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05519_, _05518_, _05517_);
  and (_05520_, _05444_, \oc8051_golden_model_1.P1INREG [7]);
  not (_05521_, _05520_);
  and (_05522_, _04552_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05523_, _05440_, \oc8051_golden_model_1.TCON [7]);
  nor (_05524_, _05523_, _05522_);
  and (_05525_, _05524_, _05521_);
  and (_05526_, _05525_, _05519_);
  and (_05527_, _05526_, _05516_);
  and (_05528_, _05527_, _05513_);
  and (_05529_, _05528_, _04427_);
  nor (_05530_, _05529_, _05506_);
  nor (_05531_, _05530_, _05505_);
  and (_05532_, _05531_, _05479_);
  not (_05533_, _04633_);
  and (_05534_, _05425_, \oc8051_golden_model_1.IP [0]);
  and (_05535_, _05419_, \oc8051_golden_model_1.B [0]);
  nor (_05536_, _05535_, _05534_);
  and (_05537_, _05417_, \oc8051_golden_model_1.PSW [0]);
  and (_05538_, _05427_, \oc8051_golden_model_1.ACC [0]);
  nor (_05539_, _05538_, _05537_);
  and (_05540_, _05539_, _05536_);
  and (_05541_, _05431_, \oc8051_golden_model_1.SCON [0]);
  and (_05542_, _05433_, \oc8051_golden_model_1.IE [0]);
  nor (_05543_, _05542_, _05541_);
  and (_05544_, _05436_, \oc8051_golden_model_1.P2INREG [0]);
  and (_05545_, _05446_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_05546_, _05545_, _05544_);
  and (_05547_, _05444_, \oc8051_golden_model_1.P1INREG [0]);
  not (_05548_, _05547_);
  and (_05549_, _04552_, \oc8051_golden_model_1.P0INREG [0]);
  and (_05550_, _05440_, \oc8051_golden_model_1.TCON [0]);
  nor (_05551_, _05550_, _05549_);
  and (_05552_, _05551_, _05548_);
  and (_05553_, _05552_, _05546_);
  and (_05554_, _05553_, _05543_);
  and (_05555_, _05554_, _05540_);
  and (_05556_, _05555_, _04836_);
  nor (_05557_, _05556_, _05533_);
  and (_05558_, _05425_, \oc8051_golden_model_1.IP [6]);
  and (_05559_, _05419_, \oc8051_golden_model_1.B [6]);
  nor (_05560_, _05559_, _05558_);
  and (_05561_, _05433_, \oc8051_golden_model_1.IE [6]);
  and (_05562_, _05417_, \oc8051_golden_model_1.PSW [6]);
  nor (_05563_, _05562_, _05561_);
  and (_05564_, _05431_, \oc8051_golden_model_1.SCON [6]);
  and (_05566_, _05427_, \oc8051_golden_model_1.ACC [6]);
  nor (_05568_, _05566_, _05564_);
  and (_05570_, _05568_, _05563_);
  and (_05572_, _05570_, _05560_);
  and (_05574_, _05436_, \oc8051_golden_model_1.P2INREG [6]);
  and (_05576_, _05446_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_05578_, _05576_, _05574_);
  and (_05580_, _05444_, \oc8051_golden_model_1.P1INREG [6]);
  not (_05582_, _05580_);
  and (_05584_, _04552_, \oc8051_golden_model_1.P0INREG [6]);
  and (_05586_, _05440_, \oc8051_golden_model_1.TCON [6]);
  nor (_05588_, _05586_, _05584_);
  and (_05590_, _05588_, _05582_);
  and (_05592_, _05590_, _05578_);
  and (_05594_, _05592_, _05572_);
  and (_05596_, _05594_, _04890_);
  and (_05598_, _04553_, _04123_);
  not (_05600_, _05598_);
  nor (_05602_, _05600_, _05596_);
  nor (_05604_, _05602_, _05557_);
  not (_05606_, _04559_);
  and (_05608_, _05425_, \oc8051_golden_model_1.IP [3]);
  and (_05610_, _05427_, \oc8051_golden_model_1.ACC [3]);
  nor (_05612_, _05610_, _05608_);
  and (_05614_, _05417_, \oc8051_golden_model_1.PSW [3]);
  and (_05616_, _05419_, \oc8051_golden_model_1.B [3]);
  nor (_05618_, _05616_, _05614_);
  and (_05620_, _05618_, _05612_);
  and (_05622_, _05431_, \oc8051_golden_model_1.SCON [3]);
  and (_05624_, _05433_, \oc8051_golden_model_1.IE [3]);
  nor (_05626_, _05624_, _05622_);
  and (_05627_, _05436_, \oc8051_golden_model_1.P2INREG [3]);
  not (_05629_, _05627_);
  and (_05630_, _04552_, \oc8051_golden_model_1.P0INREG [3]);
  and (_05632_, _05440_, \oc8051_golden_model_1.TCON [3]);
  nor (_05633_, _05632_, _05630_);
  and (_05635_, _05633_, _05629_);
  and (_05637_, _05444_, \oc8051_golden_model_1.P1INREG [3]);
  and (_05638_, _05446_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_05640_, _05638_, _05637_);
  and (_05641_, _05640_, _05635_);
  and (_05643_, _05641_, _05626_);
  and (_05644_, _05643_, _05620_);
  and (_05646_, _05644_, _04548_);
  nor (_05647_, _05646_, _05606_);
  and (_05649_, _05425_, \oc8051_golden_model_1.IP [5]);
  and (_05650_, _05419_, \oc8051_golden_model_1.B [5]);
  nor (_05652_, _05650_, _05649_);
  and (_05653_, _05417_, \oc8051_golden_model_1.PSW [5]);
  and (_05655_, _05427_, \oc8051_golden_model_1.ACC [5]);
  nor (_05656_, _05655_, _05653_);
  and (_05658_, _05656_, _05652_);
  and (_05660_, _05431_, \oc8051_golden_model_1.SCON [5]);
  and (_05662_, _05433_, \oc8051_golden_model_1.IE [5]);
  nor (_05664_, _05662_, _05660_);
  and (_05666_, _05436_, \oc8051_golden_model_1.P2INREG [5]);
  and (_05668_, _05446_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_05670_, _05668_, _05666_);
  and (_05672_, _05444_, \oc8051_golden_model_1.P1INREG [5]);
  not (_05674_, _05672_);
  and (_05676_, _04552_, \oc8051_golden_model_1.P0INREG [5]);
  and (_05678_, _05440_, \oc8051_golden_model_1.TCON [5]);
  nor (_05680_, _05678_, _05676_);
  and (_05682_, _05680_, _05674_);
  and (_05684_, _05682_, _05670_);
  and (_05686_, _05684_, _05664_);
  and (_05688_, _05686_, _05658_);
  and (_05690_, _05688_, _04742_);
  and (_05692_, _04562_, _04123_);
  not (_05694_, _05692_);
  nor (_05696_, _05694_, _05690_);
  nor (_05698_, _05696_, _05647_);
  and (_05700_, _05698_, _05604_);
  and (_05702_, _05700_, _05532_);
  not (_05704_, _05702_);
  or (_05706_, _05704_, _03102_);
  or (_05708_, _05702_, _02596_);
  and (_05710_, _05708_, _02653_);
  and (_05712_, _05710_, _05706_);
  or (_05714_, _05712_, _05412_);
  or (_05716_, _05714_, _05411_);
  and (_05718_, _05716_, _01931_);
  and (_05720_, _04513_, _01898_);
  or (_05722_, _05720_, _05718_);
  and (_05724_, _02572_, _01898_);
  not (_05726_, _05724_);
  not (_05728_, _05720_);
  or (_05730_, _05728_, _02555_);
  and (_05732_, _05730_, _05726_);
  and (_05734_, _05732_, _05722_);
  and (_05736_, _05724_, _01914_);
  or (_05738_, _05736_, _03108_);
  or (_05740_, _05738_, _05734_);
  nand (_05742_, _04426_, _03108_);
  and (_05744_, _05742_, _05740_);
  or (_05746_, _05744_, _01899_);
  not (_05748_, _01899_);
  or (_05750_, _02555_, _05748_);
  and (_05752_, _05750_, _03125_);
  and (_05754_, _05752_, _05746_);
  nand (_05756_, _05702_, _03096_);
  or (_05758_, _05702_, _03102_);
  and (_05760_, _05758_, _05756_);
  and (_05762_, _05760_, _02647_);
  nor (_05764_, _03502_, _01925_);
  or (_05766_, _05764_, _05762_);
  or (_05768_, _05766_, _05754_);
  not (_05770_, _05764_);
  or (_05772_, _05770_, _01914_);
  and (_05774_, _05772_, _03124_);
  and (_05776_, _05774_, _05768_);
  and (_05778_, _03123_, _02555_);
  nor (_05780_, _04991_, _03502_);
  or (_05782_, _05780_, _05778_);
  or (_05784_, _05782_, _05776_);
  not (_05786_, _02646_);
  not (_05788_, _05780_);
  or (_05790_, _05788_, _01914_);
  and (_05792_, _05790_, _05786_);
  and (_05794_, _05792_, _05784_);
  nor (_05796_, _05786_, _02204_);
  or (_05798_, _05796_, _01971_);
  or (_05800_, _05798_, _05794_);
  not (_05802_, _01971_);
  or (_05804_, _02555_, _05802_);
  and (_05806_, _05804_, _03122_);
  and (_05808_, _05806_, _05800_);
  and (_05810_, _05760_, _02650_);
  and (_05812_, _01954_, _02674_);
  not (_05814_, _05812_);
  and (_05816_, _01954_, _02640_);
  nor (_05818_, _02633_, _01927_);
  nor (_05820_, _05818_, _03510_);
  nor (_05822_, _05820_, _05816_);
  and (_05824_, _05822_, _05814_);
  not (_05826_, _05824_);
  or (_05828_, _05826_, _05810_);
  or (_05830_, _05828_, _05808_);
  or (_05832_, _05824_, _01914_);
  and (_05834_, _05832_, _03513_);
  and (_05836_, _05834_, _05830_);
  and (_05838_, _03121_, _02555_);
  nor (_05840_, _04991_, _03510_);
  or (_05842_, _05840_, _05838_);
  or (_05844_, _05842_, _05836_);
  not (_05846_, _02649_);
  not (_05848_, _05840_);
  or (_05850_, _05848_, _01914_);
  and (_05852_, _05850_, _05846_);
  and (_05854_, _05852_, _05844_);
  nor (_05856_, _05846_, _02204_);
  or (_05858_, _05856_, _01955_);
  or (_05860_, _05858_, _05854_);
  and (_05862_, _02566_, _01954_);
  not (_05864_, _05862_);
  or (_05866_, _02555_, _01956_);
  and (_05868_, _05866_, _05864_);
  and (_05870_, _05868_, _05860_);
  and (_05872_, _05862_, _01914_);
  or (_05874_, _05872_, _05870_);
  or (_05876_, _05874_, _27789_);
  or (_05878_, _27788_, \oc8051_golden_model_1.PC [15]);
  and (_05880_, _05878_, _27053_);
  and (_26394_, _05880_, _05876_);
  not (_05883_, _03239_);
  not (_05885_, \oc8051_golden_model_1.TMOD [7]);
  nor (_05887_, _04605_, _05885_);
  not (_05889_, _02752_);
  and (_05891_, _04605_, _05889_);
  nor (_05893_, _05891_, _05887_);
  and (_05895_, _05893_, _02575_);
  and (_05897_, _04605_, \oc8051_golden_model_1.ACC [7]);
  nor (_05899_, _05897_, _05887_);
  nor (_05901_, _05899_, _03179_);
  not (_05903_, _04505_);
  nor (_05905_, _05899_, _05903_);
  nor (_05907_, _04505_, _05885_);
  or (_05909_, _05907_, _05905_);
  and (_05911_, _05909_, _02662_);
  not (_05913_, _04605_);
  not (_05915_, _04888_);
  and (_05917_, _05915_, _04835_);
  and (_05919_, _05917_, _04789_);
  and (_05921_, _05919_, _04937_);
  nor (_05923_, _05921_, _04982_);
  and (_05925_, _05921_, _04982_);
  nor (_05927_, _05925_, _05923_);
  nor (_05929_, _05927_, _05913_);
  nor (_05931_, _05929_, _05887_);
  nor (_05933_, _05931_, _02662_);
  or (_05935_, _05933_, _05911_);
  and (_05937_, _05935_, _03365_);
  nor (_05939_, _05913_, _04426_);
  nor (_05941_, _05939_, _05887_);
  nor (_05943_, _05941_, _03365_);
  nor (_05945_, _05943_, _05937_);
  nor (_05947_, _05945_, _03168_);
  and (_05949_, _01959_, _01704_);
  or (_05951_, _05949_, _05947_);
  nor (_05953_, _05951_, _05901_);
  and (_05955_, _05949_, _05941_);
  nor (_05957_, _05955_, _05953_);
  and (_05959_, _01959_, _02674_);
  nor (_05961_, _05959_, _05957_);
  and (_05962_, _04605_, _04067_);
  not (_05963_, _05959_);
  nor (_05964_, _05963_, _05887_);
  not (_05965_, _05964_);
  nor (_05966_, _05965_, _05962_);
  or (_05967_, _05966_, _02024_);
  nor (_05968_, _05967_, _05961_);
  nor (_05969_, _04426_, _05889_);
  and (_05970_, _02981_, _02945_);
  and (_05971_, _03048_, _03016_);
  and (_05972_, _05971_, _05970_);
  and (_05973_, _02834_, _05889_);
  not (_05974_, _02910_);
  and (_05975_, _05974_, _02873_);
  and (_05976_, _05975_, _05973_);
  and (_05977_, _05976_, _05972_);
  and (_05978_, _05977_, \oc8051_golden_model_1.P1INREG [7]);
  not (_05979_, _05978_);
  and (_05980_, _02910_, _02873_);
  and (_05981_, _05980_, _05973_);
  and (_05982_, _05981_, _05972_);
  and (_05983_, _05982_, \oc8051_golden_model_1.P0INREG [7]);
  not (_05984_, _03016_);
  and (_05985_, _03048_, _05984_);
  not (_05986_, _02945_);
  and (_05987_, _02981_, _05986_);
  and (_05988_, _05987_, _05985_);
  and (_05989_, _05988_, _05981_);
  and (_05990_, _05989_, \oc8051_golden_model_1.TL0 [7]);
  nor (_05991_, _05990_, _05983_);
  and (_05992_, _05991_, _05979_);
  and (_05993_, _05987_, _05971_);
  and (_05994_, _05993_, _05981_);
  and (_05995_, _05994_, \oc8051_golden_model_1.TCON [7]);
  not (_05996_, _03048_);
  and (_05997_, _05996_, _03016_);
  and (_05998_, _05997_, _05987_);
  and (_05999_, _05998_, _05981_);
  and (_06000_, _05999_, \oc8051_golden_model_1.TMOD [7]);
  nor (_06001_, _06000_, _05995_);
  and (_06002_, _05993_, _05976_);
  and (_06003_, _06002_, \oc8051_golden_model_1.SCON [7]);
  and (_06004_, _05998_, _05976_);
  and (_06005_, _06004_, \oc8051_golden_model_1.SBUF [7]);
  nor (_06006_, _06005_, _06003_);
  and (_06007_, _06006_, _06001_);
  and (_06008_, _06007_, _05992_);
  not (_06009_, _02981_);
  nor (_06010_, _03048_, _03016_);
  and (_06011_, _06010_, _05981_);
  and (_06012_, _06011_, _02945_);
  and (_06013_, _06012_, _06009_);
  and (_06014_, _06013_, \oc8051_golden_model_1.PCON [7]);
  and (_06015_, _06012_, _02981_);
  and (_06016_, _06015_, \oc8051_golden_model_1.DPH [7]);
  nor (_06017_, _06016_, _06014_);
  and (_06018_, _06017_, _06008_);
  and (_06019_, _05981_, _05970_);
  and (_06020_, _06019_, _05997_);
  and (_06021_, _06020_, \oc8051_golden_model_1.SP [7]);
  not (_06022_, _06021_);
  nor (_06023_, _02981_, _02945_);
  and (_06024_, _06023_, _05981_);
  and (_06025_, _06024_, _05997_);
  and (_06026_, _06025_, \oc8051_golden_model_1.TH1 [7]);
  and (_06027_, _06011_, _05987_);
  and (_06028_, _06027_, \oc8051_golden_model_1.TL1 [7]);
  nor (_06029_, _06028_, _06026_);
  and (_06030_, _06029_, _06022_);
  nor (_06031_, _02910_, _02873_);
  and (_06032_, _06031_, _05973_);
  and (_06033_, _06032_, _05972_);
  and (_06034_, _06033_, \oc8051_golden_model_1.P3INREG [7]);
  not (_06035_, _06034_);
  not (_06036_, _02873_);
  and (_06037_, _02910_, _06036_);
  and (_06038_, _06037_, _05973_);
  and (_06039_, _06038_, _05972_);
  and (_06040_, _06039_, \oc8051_golden_model_1.P2INREG [7]);
  and (_06041_, _06032_, _05993_);
  and (_06042_, _06041_, \oc8051_golden_model_1.IP [7]);
  nor (_06043_, _06042_, _06040_);
  and (_06044_, _06043_, _06035_);
  and (_06045_, _06037_, _05972_);
  nor (_06046_, _02834_, _02752_);
  and (_06047_, _06046_, _06045_);
  and (_06048_, _06047_, \oc8051_golden_model_1.ACC [7]);
  and (_06049_, _06046_, _06031_);
  and (_06050_, _06049_, _05972_);
  and (_06051_, _06050_, \oc8051_golden_model_1.B [7]);
  nor (_06052_, _06051_, _06048_);
  and (_06053_, _06038_, _05993_);
  and (_06054_, _06053_, \oc8051_golden_model_1.IE [7]);
  and (_06055_, _06046_, _05975_);
  and (_06056_, _06055_, _05972_);
  and (_06057_, _06056_, \oc8051_golden_model_1.PSW [7]);
  nor (_06058_, _06057_, _06054_);
  and (_06059_, _06058_, _06052_);
  and (_06060_, _06059_, _06044_);
  and (_06061_, _06019_, _05985_);
  and (_06062_, _06061_, \oc8051_golden_model_1.DPL [7]);
  and (_06063_, _06024_, _05971_);
  and (_06064_, _06063_, \oc8051_golden_model_1.TH0 [7]);
  nor (_06065_, _06064_, _06062_);
  and (_06066_, _06065_, _06060_);
  and (_06067_, _06066_, _06030_);
  and (_06068_, _06067_, _06018_);
  not (_06069_, _06068_);
  nor (_06070_, _06069_, _05969_);
  nor (_06071_, _06070_, _05913_);
  nor (_06072_, _06071_, _05887_);
  nor (_06073_, _06072_, _03139_);
  or (_06074_, _06073_, _02575_);
  nor (_06075_, _06074_, _05968_);
  nor (_06076_, _06075_, _05895_);
  or (_06077_, _06076_, _02656_);
  and (_06078_, _04982_, _02752_);
  nor (_06079_, _04982_, _02752_);
  nor (_06080_, _06079_, _06078_);
  and (_06081_, _06080_, _04605_);
  or (_06082_, _06081_, _05887_);
  or (_06083_, _06082_, _05305_);
  and (_06084_, _06083_, _03252_);
  and (_06085_, _06084_, _06077_);
  not (_06086_, \oc8051_golden_model_1.ACC [7]);
  and (_06087_, _04982_, _06086_);
  nor (_06088_, _04982_, _06086_);
  nor (_06089_, _06088_, _06087_);
  and (_06090_, _06089_, _04605_);
  nor (_06091_, _06090_, _05887_);
  nor (_06092_, _06091_, _03252_);
  nor (_06093_, _06092_, _06085_);
  nor (_06094_, _06093_, _02669_);
  not (_06095_, _05887_);
  and (_06096_, _06095_, _04982_);
  not (_06097_, _06096_);
  nor (_06098_, _05893_, _05332_);
  and (_06099_, _06098_, _06097_);
  nor (_06100_, _06099_, _06094_);
  nor (_06101_, _06100_, _03243_);
  or (_06102_, _06096_, _03244_);
  nor (_06103_, _06102_, _05899_);
  or (_06104_, _06103_, _02654_);
  nor (_06105_, _06104_, _06101_);
  nor (_06106_, _06078_, _05913_);
  nor (_06107_, _06106_, _05887_);
  and (_06108_, _06107_, _02654_);
  nor (_06109_, _06108_, _06105_);
  and (_06110_, _06109_, _05883_);
  nor (_06111_, _06087_, _05913_);
  nor (_06112_, _06111_, _05887_);
  nor (_06113_, _06112_, _05883_);
  or (_06114_, _06113_, _06110_);
  and (_06115_, _06114_, _03124_);
  nor (_06116_, _05931_, _03124_);
  or (_06117_, _06116_, _06115_);
  and (_06118_, _06117_, _03513_);
  not (_06119_, _04937_);
  not (_06120_, _04649_);
  not (_06121_, _04695_);
  not (_06122_, _04835_);
  and (_06123_, _04888_, _06122_);
  and (_06124_, _06123_, _06121_);
  and (_06125_, _06124_, _06120_);
  nor (_06126_, _04787_, _04741_);
  and (_06127_, _06126_, _06125_);
  and (_06128_, _06127_, _06119_);
  and (_06129_, _06128_, _04982_);
  nor (_06130_, _06128_, _04982_);
  or (_06131_, _06130_, _06129_);
  and (_06132_, _06131_, _04605_);
  nor (_06133_, _06132_, _05887_);
  nor (_06134_, _06133_, _03513_);
  or (_06135_, _06134_, _06118_);
  or (_06136_, _06135_, _27789_);
  or (_06137_, _27788_, \oc8051_golden_model_1.TMOD [7]);
  and (_06138_, _06137_, _27053_);
  and (_26395_, _06138_, _06136_);
  not (_06139_, \oc8051_golden_model_1.TL1 [7]);
  nor (_06140_, _04590_, _06139_);
  and (_06141_, _04590_, _05889_);
  nor (_06142_, _06141_, _06140_);
  and (_06143_, _06142_, _02575_);
  and (_06144_, _04590_, \oc8051_golden_model_1.ACC [7]);
  nor (_06145_, _06144_, _06140_);
  nor (_06146_, _06145_, _03179_);
  nor (_06147_, _06145_, _05903_);
  nor (_06148_, _04505_, _06139_);
  or (_06149_, _06148_, _06147_);
  and (_06150_, _06149_, _02662_);
  not (_06151_, _04590_);
  nor (_06152_, _05927_, _06151_);
  nor (_06153_, _06152_, _06140_);
  nor (_06154_, _06153_, _02662_);
  or (_06155_, _06154_, _06150_);
  and (_06156_, _06155_, _03365_);
  nor (_06157_, _06151_, _04426_);
  nor (_06158_, _06157_, _06140_);
  nor (_06159_, _06158_, _03365_);
  nor (_06160_, _06159_, _06156_);
  nor (_06161_, _06160_, _03168_);
  or (_06162_, _06161_, _05949_);
  nor (_06163_, _06162_, _06146_);
  and (_06164_, _06158_, _05949_);
  nor (_06165_, _06164_, _06163_);
  nor (_06166_, _06165_, _05959_);
  and (_06167_, _04590_, _04067_);
  nor (_06168_, _06140_, _05963_);
  not (_06169_, _06168_);
  nor (_06170_, _06169_, _06167_);
  or (_06171_, _06170_, _02024_);
  nor (_06172_, _06171_, _06166_);
  nor (_06173_, _06070_, _06151_);
  nor (_06174_, _06173_, _06140_);
  nor (_06175_, _06174_, _03139_);
  or (_06176_, _06175_, _02575_);
  nor (_06177_, _06176_, _06172_);
  nor (_06178_, _06177_, _06143_);
  or (_06179_, _06178_, _02656_);
  and (_06180_, _06080_, _04590_);
  or (_06181_, _06180_, _06140_);
  or (_06182_, _06181_, _05305_);
  and (_06183_, _06182_, _03252_);
  and (_06184_, _06183_, _06179_);
  and (_06185_, _06089_, _04590_);
  nor (_06186_, _06185_, _06140_);
  nor (_06187_, _06186_, _03252_);
  nor (_06188_, _06187_, _06184_);
  nor (_06189_, _06188_, _02669_);
  not (_06190_, _06140_);
  and (_06191_, _06190_, _04982_);
  not (_06192_, _06191_);
  nor (_06193_, _06142_, _05332_);
  and (_06194_, _06193_, _06192_);
  nor (_06195_, _06194_, _06189_);
  nor (_06196_, _06195_, _03243_);
  or (_06197_, _06191_, _03244_);
  nor (_06198_, _06197_, _06145_);
  or (_06199_, _06198_, _02654_);
  nor (_06200_, _06199_, _06196_);
  nor (_06201_, _06078_, _06151_);
  nor (_06202_, _06201_, _06140_);
  and (_06203_, _06202_, _02654_);
  nor (_06204_, _06203_, _06200_);
  and (_06205_, _06204_, _05883_);
  nor (_06206_, _06087_, _06151_);
  nor (_06207_, _06206_, _06140_);
  nor (_06208_, _06207_, _05883_);
  or (_06209_, _06208_, _06205_);
  and (_06210_, _06209_, _03124_);
  nor (_06211_, _06153_, _03124_);
  or (_06212_, _06211_, _06210_);
  and (_06213_, _06212_, _03513_);
  and (_06214_, _06131_, _04590_);
  nor (_06215_, _06214_, _06140_);
  nor (_06216_, _06215_, _03513_);
  or (_06217_, _06216_, _06213_);
  or (_06218_, _06217_, _27789_);
  or (_06219_, _27788_, \oc8051_golden_model_1.TL1 [7]);
  and (_06220_, _06219_, _27053_);
  and (_26397_, _06220_, _06218_);
  not (_06221_, \oc8051_golden_model_1.TL0 [7]);
  nor (_06222_, _04608_, _06221_);
  and (_06223_, _04608_, _05889_);
  nor (_06224_, _06223_, _06222_);
  and (_06225_, _06224_, _02575_);
  not (_06226_, _04608_);
  nor (_06227_, _06226_, _04426_);
  nor (_06228_, _06227_, _06222_);
  and (_06229_, _06228_, _05949_);
  and (_06230_, _04608_, \oc8051_golden_model_1.ACC [7]);
  nor (_06231_, _06230_, _06222_);
  nor (_06232_, _06231_, _05903_);
  nor (_06233_, _04505_, _06221_);
  or (_06234_, _06233_, _06232_);
  and (_06235_, _06234_, _02662_);
  nor (_06236_, _05927_, _06226_);
  nor (_06237_, _06236_, _06222_);
  nor (_06238_, _06237_, _02662_);
  or (_06239_, _06238_, _06235_);
  and (_06240_, _06239_, _03365_);
  nor (_06241_, _06228_, _03365_);
  nor (_06242_, _06241_, _06240_);
  nor (_06243_, _06242_, _03168_);
  nor (_06244_, _06231_, _03179_);
  nor (_06245_, _06244_, _05949_);
  not (_06246_, _06245_);
  nor (_06247_, _06246_, _06243_);
  nor (_06248_, _06247_, _06229_);
  nor (_06249_, _06248_, _05959_);
  and (_06250_, _04608_, _04067_);
  nor (_06251_, _06222_, _05963_);
  not (_06252_, _06251_);
  nor (_06253_, _06252_, _06250_);
  or (_06254_, _06253_, _02024_);
  nor (_06255_, _06254_, _06249_);
  nor (_06256_, _06070_, _06226_);
  nor (_06257_, _06256_, _06222_);
  nor (_06258_, _06257_, _03139_);
  or (_06259_, _06258_, _02575_);
  nor (_06260_, _06259_, _06255_);
  nor (_06261_, _06260_, _06225_);
  or (_06262_, _06261_, _02656_);
  and (_06263_, _06080_, _04608_);
  or (_06264_, _06263_, _06222_);
  or (_06265_, _06264_, _05305_);
  and (_06266_, _06265_, _03252_);
  and (_06267_, _06266_, _06262_);
  and (_06268_, _06089_, _04608_);
  nor (_06269_, _06268_, _06222_);
  nor (_06270_, _06269_, _03252_);
  nor (_06271_, _06270_, _06267_);
  nor (_06272_, _06271_, _02669_);
  not (_06273_, _06222_);
  and (_06274_, _06273_, _04982_);
  not (_06275_, _06274_);
  nor (_06276_, _06224_, _05332_);
  and (_06277_, _06276_, _06275_);
  nor (_06278_, _06277_, _06272_);
  nor (_06279_, _06278_, _03243_);
  or (_06280_, _06274_, _03244_);
  nor (_06281_, _06280_, _06231_);
  or (_06282_, _06281_, _02654_);
  nor (_06283_, _06282_, _06279_);
  nor (_06284_, _06078_, _06226_);
  nor (_06285_, _06284_, _06222_);
  and (_06286_, _06285_, _02654_);
  nor (_06287_, _06286_, _06283_);
  and (_06288_, _06287_, _05883_);
  nor (_06289_, _06087_, _06226_);
  nor (_06290_, _06289_, _06222_);
  nor (_06291_, _06290_, _05883_);
  or (_06292_, _06291_, _06288_);
  and (_06293_, _06292_, _03124_);
  nor (_06294_, _06237_, _03124_);
  or (_06295_, _06294_, _06293_);
  and (_06296_, _06295_, _03513_);
  and (_06297_, _06131_, _04608_);
  nor (_06298_, _06297_, _06222_);
  nor (_06299_, _06298_, _03513_);
  or (_06300_, _06299_, _06296_);
  or (_06301_, _06300_, _27789_);
  or (_06302_, _27788_, \oc8051_golden_model_1.TL0 [7]);
  and (_06303_, _06302_, _27053_);
  and (_26398_, _06303_, _06301_);
  not (_06304_, \oc8051_golden_model_1.TH1 [7]);
  nor (_06305_, _04594_, _06304_);
  and (_06306_, _04594_, _05889_);
  nor (_06307_, _06306_, _06305_);
  and (_06308_, _06307_, _02575_);
  and (_06309_, _04594_, \oc8051_golden_model_1.ACC [7]);
  nor (_06310_, _06309_, _06305_);
  nor (_06311_, _06310_, _03179_);
  nor (_06312_, _06310_, _05903_);
  nor (_06313_, _04505_, _06304_);
  or (_06314_, _06313_, _06312_);
  and (_06315_, _06314_, _02662_);
  not (_06316_, _04594_);
  nor (_06317_, _05927_, _06316_);
  nor (_06318_, _06317_, _06305_);
  nor (_06319_, _06318_, _02662_);
  or (_06320_, _06319_, _06315_);
  and (_06321_, _06320_, _03365_);
  nor (_06322_, _06316_, _04426_);
  nor (_06323_, _06322_, _06305_);
  nor (_06324_, _06323_, _03365_);
  nor (_06325_, _06324_, _06321_);
  nor (_06326_, _06325_, _03168_);
  or (_06327_, _06326_, _05949_);
  nor (_06328_, _06327_, _06311_);
  and (_06329_, _06323_, _05949_);
  nor (_06330_, _06329_, _06328_);
  nor (_06331_, _06330_, _05959_);
  and (_06332_, _04594_, _04067_);
  nor (_06333_, _06305_, _05963_);
  not (_06334_, _06333_);
  nor (_06335_, _06334_, _06332_);
  or (_06336_, _06335_, _02024_);
  nor (_06337_, _06336_, _06331_);
  nor (_06338_, _06070_, _06316_);
  nor (_06339_, _06338_, _06305_);
  nor (_06340_, _06339_, _03139_);
  or (_06341_, _06340_, _02575_);
  nor (_06342_, _06341_, _06337_);
  nor (_06343_, _06342_, _06308_);
  or (_06344_, _06343_, _02656_);
  and (_06345_, _06080_, _04594_);
  or (_06346_, _06345_, _06305_);
  or (_06347_, _06346_, _05305_);
  and (_06348_, _06347_, _03252_);
  and (_06349_, _06348_, _06344_);
  and (_06350_, _06089_, _04594_);
  nor (_06351_, _06350_, _06305_);
  nor (_06352_, _06351_, _03252_);
  nor (_06353_, _06352_, _06349_);
  nor (_06354_, _06353_, _02669_);
  not (_06355_, _06305_);
  and (_06356_, _06355_, _04982_);
  not (_06357_, _06356_);
  nor (_06358_, _06307_, _05332_);
  and (_06359_, _06358_, _06357_);
  nor (_06360_, _06359_, _06354_);
  nor (_06361_, _06360_, _03243_);
  or (_06363_, _06356_, _03244_);
  nor (_06364_, _06363_, _06310_);
  or (_06365_, _06364_, _02654_);
  nor (_06366_, _06365_, _06361_);
  nor (_06367_, _06078_, _06316_);
  nor (_06368_, _06367_, _06305_);
  and (_06369_, _06368_, _02654_);
  nor (_06370_, _06369_, _06366_);
  and (_06371_, _06370_, _05883_);
  nor (_06372_, _06087_, _06316_);
  nor (_06374_, _06372_, _06305_);
  nor (_06375_, _06374_, _05883_);
  or (_06376_, _06375_, _06371_);
  and (_06377_, _06376_, _03124_);
  nor (_06378_, _06318_, _03124_);
  or (_06379_, _06378_, _06377_);
  and (_06380_, _06379_, _03513_);
  and (_06381_, _06131_, _04594_);
  nor (_06382_, _06381_, _06305_);
  nor (_06383_, _06382_, _03513_);
  or (_06385_, _06383_, _06380_);
  or (_06386_, _06385_, _27789_);
  or (_06387_, _27788_, \oc8051_golden_model_1.TH1 [7]);
  and (_06388_, _06387_, _27053_);
  and (_26399_, _06388_, _06386_);
  not (_06389_, \oc8051_golden_model_1.TH0 [7]);
  nor (_06390_, _04612_, _06389_);
  and (_06391_, _04612_, _05889_);
  nor (_06392_, _06391_, _06390_);
  and (_06393_, _06392_, _02575_);
  and (_06395_, _04612_, \oc8051_golden_model_1.ACC [7]);
  nor (_06396_, _06395_, _06390_);
  nor (_06397_, _06396_, _03179_);
  nor (_06398_, _06396_, _05903_);
  nor (_06399_, _04505_, _06389_);
  or (_06400_, _06399_, _06398_);
  and (_06401_, _06400_, _02662_);
  not (_06402_, _04612_);
  nor (_06403_, _05927_, _06402_);
  nor (_06404_, _06403_, _06390_);
  nor (_06406_, _06404_, _02662_);
  or (_06407_, _06406_, _06401_);
  and (_06408_, _06407_, _03365_);
  nor (_06409_, _06402_, _04426_);
  nor (_06410_, _06409_, _06390_);
  nor (_06411_, _06410_, _03365_);
  nor (_06412_, _06411_, _06408_);
  nor (_06413_, _06412_, _03168_);
  or (_06414_, _06413_, _05949_);
  nor (_06415_, _06414_, _06397_);
  and (_06417_, _06410_, _05949_);
  nor (_06418_, _06417_, _06415_);
  nor (_06419_, _06418_, _05959_);
  and (_06420_, _04612_, _04067_);
  nor (_06421_, _06390_, _05963_);
  not (_06422_, _06421_);
  nor (_06423_, _06422_, _06420_);
  or (_06424_, _06423_, _02024_);
  nor (_06425_, _06424_, _06419_);
  nor (_06426_, _06070_, _06402_);
  nor (_06427_, _06426_, _06390_);
  nor (_06428_, _06427_, _03139_);
  or (_06429_, _06428_, _02575_);
  nor (_06430_, _06429_, _06425_);
  nor (_06431_, _06430_, _06393_);
  or (_06432_, _06431_, _02656_);
  and (_06433_, _06080_, _04612_);
  or (_06434_, _06433_, _06390_);
  or (_06435_, _06434_, _05305_);
  and (_06436_, _06435_, _03252_);
  and (_06437_, _06436_, _06432_);
  and (_06438_, _06089_, _04612_);
  nor (_06439_, _06438_, _06390_);
  nor (_06440_, _06439_, _03252_);
  nor (_06441_, _06440_, _06437_);
  nor (_06442_, _06441_, _02669_);
  not (_06443_, _06390_);
  and (_06444_, _06443_, _04982_);
  not (_06445_, _06444_);
  nor (_06446_, _06392_, _05332_);
  and (_06447_, _06446_, _06445_);
  nor (_06448_, _06447_, _06442_);
  nor (_06449_, _06448_, _03243_);
  or (_06450_, _06444_, _03244_);
  nor (_06451_, _06450_, _06396_);
  or (_06452_, _06451_, _02654_);
  nor (_06453_, _06452_, _06449_);
  nor (_06454_, _06078_, _06402_);
  nor (_06455_, _06454_, _06390_);
  and (_06456_, _06455_, _02654_);
  nor (_06457_, _06456_, _06453_);
  and (_06458_, _06457_, _05883_);
  nor (_06459_, _06087_, _06402_);
  nor (_06460_, _06459_, _06390_);
  nor (_06461_, _06460_, _05883_);
  or (_06462_, _06461_, _06458_);
  and (_06463_, _06462_, _03124_);
  nor (_06464_, _06404_, _03124_);
  or (_06465_, _06464_, _06463_);
  and (_06466_, _06465_, _03513_);
  and (_06467_, _06131_, _04612_);
  nor (_06468_, _06467_, _06390_);
  nor (_06469_, _06468_, _03513_);
  or (_06470_, _06469_, _06466_);
  or (_06471_, _06470_, _27789_);
  or (_06472_, _27788_, \oc8051_golden_model_1.TH0 [7]);
  and (_06473_, _06472_, _27053_);
  and (_26400_, _06473_, _06471_);
  not (_06474_, \oc8051_golden_model_1.TCON [7]);
  nor (_06475_, _04597_, _06474_);
  not (_06476_, _04597_);
  nor (_06477_, _06476_, _04426_);
  nor (_06478_, _06477_, _06475_);
  and (_06479_, _06478_, _05949_);
  nor (_06480_, _05440_, _06474_);
  not (_06481_, _06480_);
  and (_06482_, _05446_, \oc8051_golden_model_1.P3 [7]);
  not (_06483_, _06482_);
  and (_06484_, _04552_, \oc8051_golden_model_1.P0 [7]);
  nor (_06485_, _06484_, _05523_);
  and (_06486_, _06485_, _06483_);
  and (_06487_, _05444_, \oc8051_golden_model_1.P1 [7]);
  and (_06488_, _05436_, \oc8051_golden_model_1.P2 [7]);
  nor (_06489_, _06488_, _06487_);
  and (_06490_, _06489_, _06486_);
  and (_06491_, _06490_, _05516_);
  and (_06492_, _06491_, _05513_);
  and (_06493_, _06492_, _04427_);
  nor (_06494_, _06493_, _05506_);
  and (_06495_, _06494_, _06481_);
  nand (_06496_, _06493_, _05506_);
  and (_06497_, _06496_, _05440_);
  nor (_06498_, _06497_, _06480_);
  or (_06499_, _06498_, _05168_);
  nor (_06500_, _06499_, _06495_);
  nor (_06501_, _05927_, _06476_);
  nor (_06502_, _06501_, _06475_);
  and (_06503_, _06502_, _02661_);
  not (_06504_, _03163_);
  and (_06505_, _04597_, \oc8051_golden_model_1.ACC [7]);
  nor (_06506_, _06505_, _06475_);
  nor (_06507_, _06506_, _05903_);
  nor (_06508_, _04505_, _06474_);
  or (_06509_, _06508_, _02661_);
  nor (_06510_, _06509_, _06507_);
  or (_06511_, _06510_, _06504_);
  nor (_06512_, _06511_, _06503_);
  nor (_06513_, _06478_, _03365_);
  nor (_06514_, _06498_, _03390_);
  nor (_06515_, _06514_, _06513_);
  nand (_06516_, _06515_, _03179_);
  or (_06517_, _06516_, _06512_);
  nand (_06518_, _06506_, _03168_);
  and (_06519_, _06518_, _06517_);
  and (_06520_, _06519_, _03177_);
  nor (_06521_, _06493_, _04622_);
  and (_06522_, _06521_, _05440_);
  nor (_06523_, _06522_, _06480_);
  nor (_06524_, _06523_, _03177_);
  or (_06525_, _06524_, _06520_);
  and (_06526_, _06525_, _05168_);
  nor (_06527_, _06526_, _06500_);
  nor (_06528_, _06527_, _03140_);
  not (_06529_, _05440_);
  nor (_06530_, _05529_, _04622_);
  and (_06531_, _04558_, \oc8051_golden_model_1.PSW [7]);
  and (_06532_, _06531_, _04123_);
  nor (_06533_, _06532_, _06530_);
  nor (_06534_, _06533_, _06529_);
  nor (_06535_, _06534_, _06480_);
  nor (_06536_, _06535_, _03141_);
  nor (_06537_, _06536_, _05949_);
  not (_06538_, _06537_);
  nor (_06539_, _06538_, _06528_);
  nor (_06540_, _06539_, _06479_);
  nor (_06541_, _06540_, _05959_);
  and (_06542_, _04597_, _04067_);
  nor (_06543_, _06475_, _05963_);
  not (_06544_, _06543_);
  nor (_06545_, _06544_, _06542_);
  nor (_06546_, _06545_, _02024_);
  not (_06547_, _06546_);
  nor (_06548_, _06547_, _06541_);
  not (_06549_, _02657_);
  nor (_06550_, _06070_, _06476_);
  nor (_06551_, _06550_, _06475_);
  nor (_06552_, _06551_, _03139_);
  or (_06553_, _06552_, _06549_);
  or (_06554_, _06553_, _06548_);
  and (_06555_, _06080_, _04597_);
  or (_06556_, _06475_, _05305_);
  or (_06557_, _06556_, _06555_);
  and (_06558_, _04597_, _05889_);
  nor (_06559_, _06558_, _06475_);
  and (_06560_, _06559_, _02575_);
  nor (_06561_, _06560_, _03251_);
  and (_06562_, _06561_, _06557_);
  and (_06563_, _06562_, _06554_);
  and (_06564_, _06089_, _04597_);
  nor (_06565_, _06564_, _06475_);
  nor (_06566_, _06565_, _03252_);
  nor (_06567_, _06566_, _06563_);
  nor (_06568_, _06567_, _02669_);
  not (_06569_, _06475_);
  and (_06570_, _06569_, _04982_);
  not (_06571_, _06570_);
  nor (_06572_, _06559_, _05332_);
  and (_06573_, _06572_, _06571_);
  nor (_06574_, _06573_, _06568_);
  nor (_06575_, _06574_, _03243_);
  or (_06576_, _06570_, _03244_);
  nor (_06577_, _06576_, _06506_);
  or (_06578_, _06577_, _02654_);
  nor (_06579_, _06578_, _06575_);
  nor (_06580_, _06078_, _06476_);
  nor (_06581_, _06580_, _06475_);
  and (_06582_, _06581_, _02654_);
  nor (_06583_, _06582_, _06579_);
  and (_06584_, _06583_, _05883_);
  nor (_06585_, _06087_, _06476_);
  nor (_06586_, _06585_, _06475_);
  nor (_06587_, _06586_, _05883_);
  or (_06588_, _06587_, _06584_);
  and (_06589_, _06588_, _03124_);
  nor (_06590_, _06502_, _03124_);
  or (_06591_, _06590_, _02650_);
  or (_06592_, _06591_, _06589_);
  nand (_06593_, _06523_, _02650_);
  and (_06594_, _06593_, _06592_);
  nor (_06595_, _06594_, _03121_);
  and (_06596_, _06131_, _04597_);
  nor (_06597_, _06596_, _06475_);
  and (_06598_, _06597_, _03121_);
  nor (_06599_, _06598_, _06595_);
  or (_06600_, _06599_, _27789_);
  or (_06601_, _27788_, \oc8051_golden_model_1.TCON [7]);
  and (_06602_, _06601_, _27053_);
  and (_26402_, _06602_, _06600_);
  not (_06603_, \oc8051_golden_model_1.SP [7]);
  nor (_06604_, _04879_, _06603_);
  and (_06605_, _06131_, _04564_);
  nor (_06606_, _06605_, _06604_);
  nor (_06607_, _06606_, _03513_);
  not (_06608_, _04564_);
  nor (_06609_, _05927_, _06608_);
  nor (_06610_, _06609_, _06604_);
  nor (_06611_, _06610_, _03124_);
  not (_06612_, _03109_);
  and (_06613_, _06089_, _04564_);
  nor (_06614_, _06613_, _06604_);
  nor (_06615_, _06614_, _03252_);
  nor (_06616_, _04505_, _06603_);
  and (_06617_, _04879_, \oc8051_golden_model_1.ACC [7]);
  nor (_06618_, _06617_, _06604_);
  nor (_06619_, _06618_, _05903_);
  or (_06620_, _06619_, _06616_);
  and (_06621_, _06620_, _01988_);
  and (_06622_, \oc8051_golden_model_1.SP [3], \oc8051_golden_model_1.SP [2]);
  and (_06623_, _06622_, \oc8051_golden_model_1.SP [1]);
  and (_06624_, _06623_, \oc8051_golden_model_1.SP [4]);
  and (_06625_, _06624_, \oc8051_golden_model_1.SP [5]);
  and (_06626_, _06625_, \oc8051_golden_model_1.SP [6]);
  nor (_06627_, _06626_, \oc8051_golden_model_1.SP [7]);
  and (_06628_, _06626_, \oc8051_golden_model_1.SP [7]);
  nor (_06629_, _06628_, _06627_);
  not (_06630_, _06629_);
  nor (_06631_, _06630_, _01988_);
  nor (_06632_, _06631_, _06621_);
  nor (_06633_, _06632_, _02661_);
  nor (_06634_, _06610_, _02662_);
  or (_06635_, _06634_, _06633_);
  and (_06636_, _06635_, _01995_);
  nor (_06637_, _06630_, _01995_);
  or (_06638_, _06637_, _06636_);
  and (_06639_, _06638_, _03365_);
  not (_06640_, \oc8051_golden_model_1.SP [6]);
  not (_06641_, \oc8051_golden_model_1.SP [5]);
  not (_06642_, \oc8051_golden_model_1.SP [4]);
  and (_06643_, _03803_, _06642_);
  and (_06644_, _06643_, _06641_);
  and (_06645_, _06644_, _06640_);
  and (_06646_, _06645_, _03417_);
  nor (_06647_, _06646_, _06603_);
  and (_06648_, _06646_, _06603_);
  nor (_06649_, _06648_, _06647_);
  nor (_06650_, _06649_, _03365_);
  or (_06651_, _06650_, _06639_);
  and (_06652_, _06651_, _03179_);
  nor (_06653_, _06618_, _03179_);
  or (_06654_, _06653_, _06652_);
  and (_06655_, _06654_, _03430_);
  nand (_06656_, _06622_, _03782_);
  nor (_06657_, _06656_, _06642_);
  and (_06658_, _06657_, \oc8051_golden_model_1.SP [5]);
  and (_06659_, _06658_, \oc8051_golden_model_1.SP [6]);
  nor (_06660_, _06659_, \oc8051_golden_model_1.SP [7]);
  and (_06661_, _06659_, \oc8051_golden_model_1.SP [7]);
  nor (_06662_, _06661_, _06660_);
  and (_06663_, _06662_, _03187_);
  not (_06664_, _02000_);
  nor (_06665_, _02025_, _06664_);
  not (_06666_, _06665_);
  nor (_06667_, _06666_, _06663_);
  not (_06668_, _06667_);
  nor (_06669_, _06668_, _06655_);
  nor (_06670_, _06665_, _06629_);
  or (_06671_, _06670_, _05949_);
  nor (_06672_, _06671_, _06669_);
  not (_06673_, _05949_);
  nor (_06674_, _06608_, _04426_);
  nor (_06675_, _06674_, _06604_);
  nor (_06676_, _06675_, _06673_);
  nor (_06677_, _06676_, _05959_);
  not (_06678_, _06677_);
  nor (_06679_, _06678_, _06672_);
  nor (_06680_, _06604_, _05963_);
  or (_06681_, _06608_, _04069_);
  and (_06682_, _06681_, _06680_);
  nor (_06683_, _06682_, _02024_);
  not (_06684_, _06683_);
  nor (_06685_, _06684_, _06679_);
  nor (_06686_, _06070_, _06608_);
  nor (_06687_, _06686_, _06604_);
  nor (_06688_, _06687_, _03139_);
  or (_06689_, _06688_, _02575_);
  or (_06690_, _06689_, _06685_);
  and (_06691_, _04879_, _05889_);
  nor (_06692_, _06691_, _06604_);
  nand (_06693_, _06692_, _02575_);
  and (_06694_, _06693_, _06690_);
  nor (_06695_, _06694_, _01967_);
  and (_06696_, _06630_, _01967_);
  nor (_06697_, _06696_, _06695_);
  and (_06698_, _06697_, _05305_);
  and (_06699_, _06080_, _04879_);
  nor (_06700_, _06699_, _06604_);
  nor (_06701_, _06700_, _05305_);
  or (_06702_, _06701_, _06698_);
  and (_06703_, _06702_, _03252_);
  nor (_06704_, _06703_, _06615_);
  nor (_06705_, _06704_, _02669_);
  not (_06706_, _06604_);
  and (_06707_, _06706_, _04982_);
  or (_06708_, _06707_, _05332_);
  nor (_06709_, _06708_, _06692_);
  nor (_06710_, _06709_, _06705_);
  nor (_06711_, _06710_, _05339_);
  and (_06712_, _06629_, _01965_);
  nor (_06713_, _06712_, _02654_);
  or (_06714_, _06618_, _03244_);
  or (_06715_, _06714_, _06707_);
  nand (_06716_, _06715_, _06713_);
  nor (_06717_, _06716_, _06711_);
  not (_06718_, _04879_);
  nor (_06719_, _06078_, _06718_);
  nor (_06720_, _06719_, _06604_);
  and (_06721_, _06720_, _02654_);
  nor (_06722_, _06721_, _06717_);
  and (_06723_, _06722_, _05883_);
  nor (_06724_, _06087_, _06718_);
  nor (_06725_, _06724_, _06604_);
  nor (_06726_, _06725_, _05883_);
  or (_06727_, _06726_, _06723_);
  and (_06728_, _06727_, _06612_);
  nor (_06729_, _06645_, \oc8051_golden_model_1.SP [7]);
  and (_06730_, _06645_, \oc8051_golden_model_1.SP [7]);
  nor (_06731_, _06730_, _06729_);
  and (_06732_, _06731_, _03109_);
  or (_06733_, _06732_, _01936_);
  or (_06734_, _06733_, _06728_);
  nand (_06735_, _06630_, _01936_);
  and (_06736_, _06735_, _06734_);
  and (_06737_, _06736_, _03126_);
  and (_06738_, _06731_, _03108_);
  or (_06739_, _06738_, _06737_);
  and (_06740_, _06739_, _03124_);
  nor (_06741_, _02646_, _01971_);
  not (_06742_, _06741_);
  or (_06743_, _06742_, _06740_);
  nor (_06744_, _06743_, _06611_);
  nor (_06745_, _06741_, _06629_);
  nor (_06746_, _06745_, _03121_);
  not (_06747_, _06746_);
  nor (_06748_, _06747_, _06744_);
  nor (_06749_, _06748_, _06607_);
  nand (_06750_, _06749_, _27788_);
  or (_06751_, _27788_, \oc8051_golden_model_1.SP [7]);
  and (_06752_, _06751_, _27053_);
  and (_26403_, _06752_, _06750_);
  not (_06753_, \oc8051_golden_model_1.SCON [7]);
  nor (_06754_, _04615_, _06753_);
  not (_06755_, _04615_);
  nor (_06756_, _06755_, _04426_);
  nor (_06757_, _06756_, _06754_);
  and (_06758_, _06757_, _05949_);
  nor (_06759_, _05431_, _06753_);
  not (_06760_, _06759_);
  and (_06761_, _06760_, _06494_);
  and (_06762_, _06496_, _05431_);
  nor (_06763_, _06762_, _06759_);
  or (_06764_, _06763_, _05168_);
  nor (_06765_, _06764_, _06761_);
  nor (_06766_, _05927_, _06755_);
  nor (_06767_, _06766_, _06754_);
  and (_06768_, _06767_, _02661_);
  and (_06769_, _04615_, \oc8051_golden_model_1.ACC [7]);
  nor (_06770_, _06769_, _06754_);
  nor (_06771_, _06770_, _05903_);
  nor (_06772_, _04505_, _06753_);
  or (_06773_, _06772_, _02661_);
  nor (_06774_, _06773_, _06771_);
  or (_06775_, _06774_, _06504_);
  nor (_06776_, _06775_, _06768_);
  nor (_06777_, _06757_, _03365_);
  nor (_06778_, _06763_, _03390_);
  nor (_06779_, _06778_, _06777_);
  nand (_06780_, _06779_, _03179_);
  or (_06781_, _06780_, _06776_);
  nand (_06782_, _06770_, _03168_);
  and (_06783_, _06782_, _06781_);
  and (_06784_, _06783_, _03177_);
  and (_06785_, _06521_, _05431_);
  nor (_06786_, _06785_, _06759_);
  nor (_06787_, _06786_, _03177_);
  or (_06788_, _06787_, _06784_);
  and (_06789_, _06788_, _05168_);
  nor (_06790_, _06789_, _06765_);
  nor (_06791_, _06790_, _03140_);
  not (_06792_, _05431_);
  nor (_06793_, _06533_, _06792_);
  nor (_06794_, _06793_, _06759_);
  nor (_06795_, _06794_, _03141_);
  nor (_06796_, _06795_, _05949_);
  not (_06797_, _06796_);
  nor (_06798_, _06797_, _06791_);
  nor (_06799_, _06798_, _06758_);
  nor (_06800_, _06799_, _05959_);
  and (_06801_, _04615_, _04067_);
  nor (_06802_, _06754_, _05963_);
  not (_06803_, _06802_);
  nor (_06804_, _06803_, _06801_);
  nor (_06805_, _06804_, _02024_);
  not (_06806_, _06805_);
  nor (_06807_, _06806_, _06800_);
  nor (_06808_, _06070_, _06755_);
  nor (_06809_, _06808_, _06754_);
  nor (_06810_, _06809_, _03139_);
  or (_06811_, _06810_, _06549_);
  or (_06812_, _06811_, _06807_);
  and (_06813_, _06080_, _04615_);
  or (_06814_, _06754_, _05305_);
  or (_06815_, _06814_, _06813_);
  and (_06816_, _04615_, _05889_);
  nor (_06817_, _06816_, _06754_);
  and (_06818_, _06817_, _02575_);
  nor (_06819_, _06818_, _03251_);
  and (_06820_, _06819_, _06815_);
  and (_06821_, _06820_, _06812_);
  and (_06822_, _06089_, _04615_);
  nor (_06823_, _06822_, _06754_);
  nor (_06824_, _06823_, _03252_);
  nor (_06825_, _06824_, _06821_);
  nor (_06826_, _06825_, _02669_);
  not (_06827_, _06754_);
  and (_06828_, _06827_, _04982_);
  not (_06829_, _06828_);
  nor (_06830_, _06817_, _05332_);
  and (_06831_, _06830_, _06829_);
  nor (_06832_, _06831_, _06826_);
  nor (_06833_, _06832_, _03243_);
  or (_06834_, _06828_, _03244_);
  nor (_06835_, _06834_, _06770_);
  or (_06836_, _06835_, _02654_);
  nor (_06837_, _06836_, _06833_);
  nor (_06838_, _06078_, _06755_);
  nor (_06839_, _06838_, _06754_);
  and (_06840_, _06839_, _02654_);
  nor (_06841_, _06840_, _06837_);
  and (_06842_, _06841_, _05883_);
  nor (_06843_, _06087_, _06755_);
  nor (_06844_, _06843_, _06754_);
  nor (_06845_, _06844_, _05883_);
  or (_06846_, _06845_, _06842_);
  and (_06847_, _06846_, _03124_);
  nor (_06848_, _06767_, _03124_);
  or (_06849_, _06848_, _02650_);
  or (_06850_, _06849_, _06847_);
  nand (_06851_, _06786_, _02650_);
  and (_06852_, _06851_, _06850_);
  nor (_06853_, _06852_, _03121_);
  and (_06854_, _06131_, _04615_);
  nor (_06855_, _06854_, _06754_);
  and (_06856_, _06855_, _03121_);
  nor (_06857_, _06856_, _06853_);
  or (_06858_, _06857_, _27789_);
  or (_06859_, _27788_, \oc8051_golden_model_1.SCON [7]);
  and (_06860_, _06859_, _27053_);
  and (_26404_, _06860_, _06858_);
  not (_06861_, \oc8051_golden_model_1.SBUF [7]);
  nor (_06862_, _04626_, _06861_);
  and (_06863_, _04626_, _05889_);
  nor (_06864_, _06863_, _06862_);
  and (_06865_, _06864_, _02575_);
  not (_06866_, _04626_);
  nor (_06867_, _06866_, _04426_);
  nor (_06868_, _06867_, _06862_);
  and (_06869_, _06868_, _05949_);
  and (_06870_, _04626_, \oc8051_golden_model_1.ACC [7]);
  nor (_06871_, _06870_, _06862_);
  nor (_06872_, _06871_, _05903_);
  nor (_06873_, _04505_, _06861_);
  or (_06874_, _06873_, _06872_);
  and (_06875_, _06874_, _02662_);
  nor (_06876_, _05927_, _06866_);
  nor (_06877_, _06876_, _06862_);
  nor (_06878_, _06877_, _02662_);
  or (_06879_, _06878_, _06875_);
  and (_06880_, _06879_, _03365_);
  nor (_06881_, _06868_, _03365_);
  nor (_06882_, _06881_, _06880_);
  nor (_06883_, _06882_, _03168_);
  nor (_06884_, _06871_, _03179_);
  nor (_06885_, _06884_, _05949_);
  not (_06886_, _06885_);
  nor (_06887_, _06886_, _06883_);
  nor (_06888_, _06887_, _06869_);
  nor (_06889_, _06888_, _05959_);
  and (_06890_, _04626_, _04067_);
  nor (_06891_, _06862_, _05963_);
  not (_06892_, _06891_);
  nor (_06893_, _06892_, _06890_);
  or (_06894_, _06893_, _02024_);
  nor (_06895_, _06894_, _06889_);
  nor (_06896_, _06070_, _06866_);
  nor (_06897_, _06896_, _06862_);
  nor (_06898_, _06897_, _03139_);
  or (_06899_, _06898_, _02575_);
  nor (_06900_, _06899_, _06895_);
  nor (_06901_, _06900_, _06865_);
  or (_06902_, _06901_, _02656_);
  and (_06903_, _06080_, _04626_);
  or (_06904_, _06903_, _06862_);
  or (_06905_, _06904_, _05305_);
  and (_06906_, _06905_, _03252_);
  and (_06907_, _06906_, _06902_);
  and (_06908_, _06089_, _04626_);
  nor (_06909_, _06908_, _06862_);
  nor (_06910_, _06909_, _03252_);
  nor (_06911_, _06910_, _06907_);
  nor (_06912_, _06911_, _02669_);
  not (_06913_, _06862_);
  and (_06914_, _06913_, _04982_);
  not (_06915_, _06914_);
  nor (_06916_, _06864_, _05332_);
  and (_06917_, _06916_, _06915_);
  nor (_06918_, _06917_, _06912_);
  nor (_06919_, _06918_, _03243_);
  or (_06920_, _06914_, _03244_);
  nor (_06921_, _06920_, _06871_);
  or (_06922_, _06921_, _02654_);
  nor (_06923_, _06922_, _06919_);
  nor (_06924_, _06078_, _06866_);
  nor (_06925_, _06924_, _06862_);
  and (_06926_, _06925_, _02654_);
  nor (_06927_, _06926_, _06923_);
  and (_06928_, _06927_, _05883_);
  nor (_06929_, _06087_, _06866_);
  nor (_06930_, _06929_, _06862_);
  nor (_06931_, _06930_, _05883_);
  or (_06932_, _06931_, _06928_);
  and (_06933_, _06932_, _03124_);
  nor (_06934_, _06877_, _03124_);
  or (_06935_, _06934_, _06933_);
  and (_06936_, _06935_, _03513_);
  and (_06937_, _06131_, _04626_);
  nor (_06938_, _06937_, _06862_);
  nor (_06939_, _06938_, _03513_);
  or (_06940_, _06939_, _06936_);
  or (_06941_, _06940_, _27789_);
  or (_06942_, _27788_, \oc8051_golden_model_1.SBUF [7]);
  and (_06943_, _06942_, _27053_);
  and (_26406_, _06943_, _06941_);
  not (_06944_, \oc8051_golden_model_1.PCON [7]);
  nor (_06945_, _04623_, _06944_);
  and (_06946_, _04623_, _05889_);
  nor (_06947_, _06946_, _06945_);
  and (_06948_, _06947_, _02575_);
  and (_06949_, _04623_, \oc8051_golden_model_1.ACC [7]);
  nor (_06950_, _06949_, _06945_);
  nor (_06951_, _06950_, _03179_);
  nor (_06952_, _06950_, _05903_);
  nor (_06953_, _04505_, _06944_);
  or (_06954_, _06953_, _06952_);
  and (_06955_, _06954_, _02662_);
  not (_06956_, _04623_);
  nor (_06957_, _05927_, _06956_);
  nor (_06958_, _06957_, _06945_);
  nor (_06959_, _06958_, _02662_);
  or (_06960_, _06959_, _06955_);
  and (_06961_, _06960_, _03365_);
  nor (_06962_, _06956_, _04426_);
  nor (_06963_, _06962_, _06945_);
  nor (_06964_, _06963_, _03365_);
  nor (_06965_, _06964_, _06961_);
  nor (_06966_, _06965_, _03168_);
  or (_06967_, _06966_, _05949_);
  nor (_06968_, _06967_, _06951_);
  and (_06969_, _06963_, _05949_);
  nor (_06970_, _06969_, _06968_);
  nor (_06971_, _06970_, _05959_);
  and (_06972_, _04623_, _04067_);
  nor (_06973_, _06945_, _05963_);
  not (_06974_, _06973_);
  nor (_06975_, _06974_, _06972_);
  or (_06976_, _06975_, _02024_);
  nor (_06977_, _06976_, _06971_);
  nor (_06978_, _06070_, _06956_);
  nor (_06979_, _06978_, _06945_);
  nor (_06980_, _06979_, _03139_);
  or (_06981_, _06980_, _02575_);
  nor (_06982_, _06981_, _06977_);
  nor (_06983_, _06982_, _06948_);
  or (_06984_, _06983_, _02656_);
  and (_06985_, _06080_, _04623_);
  or (_06986_, _06985_, _06945_);
  or (_06987_, _06986_, _05305_);
  and (_06988_, _06987_, _03252_);
  and (_06989_, _06988_, _06984_);
  and (_06990_, _06089_, _04623_);
  nor (_06991_, _06990_, _06945_);
  nor (_06992_, _06991_, _03252_);
  nor (_06993_, _06992_, _06989_);
  nor (_06994_, _06993_, _02669_);
  not (_06995_, _06945_);
  and (_06996_, _06995_, _04982_);
  not (_06997_, _06996_);
  nor (_06998_, _06947_, _05332_);
  and (_06999_, _06998_, _06997_);
  nor (_07000_, _06999_, _06994_);
  nor (_07001_, _07000_, _03243_);
  or (_07002_, _06996_, _03244_);
  nor (_07003_, _07002_, _06950_);
  or (_07004_, _07003_, _02654_);
  nor (_07005_, _07004_, _07001_);
  nor (_07006_, _06078_, _06956_);
  nor (_07007_, _07006_, _06945_);
  and (_07008_, _07007_, _02654_);
  nor (_07009_, _07008_, _07005_);
  and (_07010_, _07009_, _05883_);
  nor (_07011_, _06087_, _06956_);
  nor (_07012_, _07011_, _06945_);
  nor (_07013_, _07012_, _05883_);
  or (_07014_, _07013_, _07010_);
  and (_07015_, _07014_, _03124_);
  nor (_07016_, _06958_, _03124_);
  or (_07017_, _07016_, _07015_);
  and (_07018_, _07017_, _03513_);
  and (_07019_, _06131_, _04623_);
  nor (_07020_, _07019_, _06945_);
  nor (_07021_, _07020_, _03513_);
  or (_07022_, _07021_, _07018_);
  or (_07023_, _07022_, _27789_);
  or (_07024_, _27788_, \oc8051_golden_model_1.PCON [7]);
  and (_07025_, _07024_, _27053_);
  and (_26407_, _07025_, _07023_);
  or (_07026_, _05348_, rst);
  nor (_26409_, _07026_, _27788_);
  not (_07027_, \oc8051_golden_model_1.P3 [7]);
  nor (_07028_, _27788_, _07027_);
  or (_26410_, _07028_, rst);
  and (_00001_, _27788_, _27053_);
  nor (_07029_, \oc8051_golden_model_1.P2 [7], rst);
  nor (_26411_, _07029_, _00001_);
  nor (_07030_, \oc8051_golden_model_1.P1 [7], rst);
  nor (_26412_, _07030_, _00001_);
  nor (_07031_, \oc8051_golden_model_1.P0 [7], rst);
  nor (_26414_, _07031_, _00001_);
  not (_07032_, \oc8051_golden_model_1.IP [7]);
  nor (_07033_, _04581_, _07032_);
  not (_07034_, _04581_);
  nor (_07035_, _07034_, _04426_);
  nor (_07036_, _07035_, _07033_);
  and (_07037_, _07036_, _05949_);
  nor (_07038_, _05425_, _07032_);
  not (_07039_, _07038_);
  and (_07040_, _07039_, _06494_);
  and (_07041_, _06496_, _05425_);
  nor (_07042_, _07041_, _07038_);
  or (_07043_, _07042_, _05168_);
  nor (_07044_, _07043_, _07040_);
  nor (_07045_, _05927_, _07034_);
  nor (_07046_, _07045_, _07033_);
  and (_07047_, _07046_, _02661_);
  and (_07048_, _04581_, \oc8051_golden_model_1.ACC [7]);
  nor (_07049_, _07048_, _07033_);
  nor (_07050_, _07049_, _05903_);
  nor (_07051_, _04505_, _07032_);
  or (_07052_, _07051_, _02661_);
  nor (_07053_, _07052_, _07050_);
  or (_07054_, _07053_, _06504_);
  nor (_07055_, _07054_, _07047_);
  nor (_07056_, _07036_, _03365_);
  nor (_07057_, _07042_, _03390_);
  nor (_07058_, _07057_, _07056_);
  nand (_07059_, _07058_, _03179_);
  or (_07060_, _07059_, _07055_);
  nand (_07061_, _07049_, _03168_);
  and (_07062_, _07061_, _07060_);
  and (_07063_, _07062_, _03177_);
  and (_07064_, _06521_, _05425_);
  nor (_07065_, _07064_, _07038_);
  nor (_07066_, _07065_, _03177_);
  or (_07067_, _07066_, _07063_);
  and (_07068_, _07067_, _05168_);
  nor (_07069_, _07068_, _07044_);
  nor (_07070_, _07069_, _03140_);
  not (_07071_, _05425_);
  nor (_07072_, _06533_, _07071_);
  nor (_07073_, _07072_, _07038_);
  nor (_07074_, _07073_, _03141_);
  nor (_07075_, _07074_, _05949_);
  not (_07076_, _07075_);
  nor (_07077_, _07076_, _07070_);
  nor (_07078_, _07077_, _07037_);
  nor (_07079_, _07078_, _05959_);
  and (_07080_, _04581_, _04067_);
  nor (_07081_, _07033_, _05963_);
  not (_07082_, _07081_);
  nor (_07083_, _07082_, _07080_);
  nor (_07084_, _07083_, _02024_);
  not (_07085_, _07084_);
  nor (_07086_, _07085_, _07079_);
  nor (_07087_, _06070_, _07034_);
  nor (_07088_, _07087_, _07033_);
  nor (_07089_, _07088_, _03139_);
  or (_07090_, _07089_, _06549_);
  or (_07091_, _07090_, _07086_);
  and (_07092_, _06080_, _04581_);
  or (_07093_, _07033_, _05305_);
  or (_07094_, _07093_, _07092_);
  and (_07095_, _04581_, _05889_);
  nor (_07096_, _07095_, _07033_);
  and (_07097_, _07096_, _02575_);
  nor (_07098_, _07097_, _03251_);
  and (_07099_, _07098_, _07094_);
  and (_07100_, _07099_, _07091_);
  and (_07101_, _06089_, _04581_);
  nor (_07102_, _07101_, _07033_);
  nor (_07103_, _07102_, _03252_);
  nor (_07104_, _07103_, _07100_);
  nor (_07105_, _07104_, _02669_);
  not (_07106_, _07033_);
  and (_07107_, _07106_, _04982_);
  not (_07108_, _07107_);
  nor (_07109_, _07096_, _05332_);
  and (_07110_, _07109_, _07108_);
  nor (_07111_, _07110_, _07105_);
  nor (_07112_, _07111_, _03243_);
  or (_07113_, _07107_, _03244_);
  nor (_07114_, _07113_, _07049_);
  or (_07115_, _07114_, _02654_);
  nor (_07116_, _07115_, _07112_);
  nor (_07117_, _06078_, _07034_);
  nor (_07118_, _07117_, _07033_);
  and (_07119_, _07118_, _02654_);
  nor (_07120_, _07119_, _07116_);
  and (_07121_, _07120_, _05883_);
  nor (_07122_, _06087_, _07034_);
  nor (_07123_, _07122_, _07033_);
  nor (_07124_, _07123_, _05883_);
  or (_07126_, _07124_, _07121_);
  and (_07127_, _07126_, _03124_);
  nor (_07128_, _07046_, _03124_);
  or (_07129_, _07128_, _02650_);
  or (_07130_, _07129_, _07127_);
  nand (_07131_, _07065_, _02650_);
  and (_07132_, _07131_, _07130_);
  nor (_07133_, _07132_, _03121_);
  and (_07134_, _06131_, _04581_);
  nor (_07135_, _07134_, _07033_);
  and (_07136_, _07135_, _03121_);
  nor (_07137_, _07136_, _07133_);
  or (_07138_, _07137_, _27789_);
  or (_07139_, _27788_, \oc8051_golden_model_1.IP [7]);
  and (_07140_, _07139_, _27053_);
  and (_26415_, _07140_, _07138_);
  not (_07141_, \oc8051_golden_model_1.IE [7]);
  nor (_07142_, _04629_, _07141_);
  not (_07143_, _04629_);
  nor (_07144_, _07143_, _04426_);
  nor (_07145_, _07144_, _07142_);
  and (_07146_, _07145_, _05949_);
  nor (_07147_, _05433_, _07141_);
  not (_07148_, _07147_);
  and (_07149_, _07148_, _06494_);
  and (_07150_, _06496_, _05433_);
  nor (_07151_, _07150_, _07147_);
  or (_07152_, _07151_, _05168_);
  nor (_07153_, _07152_, _07149_);
  nor (_07154_, _05927_, _07143_);
  nor (_07155_, _07154_, _07142_);
  and (_07156_, _07155_, _02661_);
  and (_07157_, _04629_, \oc8051_golden_model_1.ACC [7]);
  nor (_07158_, _07157_, _07142_);
  nor (_07159_, _07158_, _05903_);
  nor (_07160_, _04505_, _07141_);
  or (_07161_, _07160_, _02661_);
  nor (_07162_, _07161_, _07159_);
  or (_07163_, _07162_, _06504_);
  nor (_07164_, _07163_, _07156_);
  nor (_07165_, _07145_, _03365_);
  nor (_07166_, _07151_, _03390_);
  nor (_07167_, _07166_, _07165_);
  nand (_07168_, _07167_, _03179_);
  or (_07169_, _07168_, _07164_);
  nand (_07170_, _07158_, _03168_);
  and (_07171_, _07170_, _07169_);
  and (_07172_, _07171_, _03177_);
  and (_07173_, _06521_, _05433_);
  nor (_07174_, _07173_, _07147_);
  nor (_07175_, _07174_, _03177_);
  or (_07176_, _07175_, _07172_);
  and (_07177_, _07176_, _05168_);
  nor (_07178_, _07177_, _07153_);
  nor (_07179_, _07178_, _03140_);
  not (_07180_, _05433_);
  nor (_07181_, _06533_, _07180_);
  nor (_07182_, _07181_, _07147_);
  nor (_07183_, _07182_, _03141_);
  nor (_07184_, _07183_, _05949_);
  not (_07185_, _07184_);
  nor (_07186_, _07185_, _07179_);
  nor (_07187_, _07186_, _07146_);
  nor (_07188_, _07187_, _05959_);
  and (_07189_, _04629_, _04067_);
  nor (_07190_, _07142_, _05963_);
  not (_07191_, _07190_);
  nor (_07192_, _07191_, _07189_);
  nor (_07193_, _07192_, _02024_);
  not (_07194_, _07193_);
  nor (_07195_, _07194_, _07188_);
  nor (_07196_, _06070_, _07143_);
  nor (_07197_, _07196_, _07142_);
  nor (_07198_, _07197_, _03139_);
  or (_07199_, _07198_, _06549_);
  or (_07200_, _07199_, _07195_);
  and (_07201_, _06080_, _04629_);
  or (_07202_, _07142_, _05305_);
  or (_07203_, _07202_, _07201_);
  and (_07204_, _04629_, _05889_);
  nor (_07205_, _07204_, _07142_);
  and (_07206_, _07205_, _02575_);
  nor (_07207_, _07206_, _03251_);
  and (_07208_, _07207_, _07203_);
  and (_07209_, _07208_, _07200_);
  and (_07210_, _06089_, _04629_);
  nor (_07211_, _07210_, _07142_);
  nor (_07212_, _07211_, _03252_);
  nor (_07213_, _07212_, _07209_);
  nor (_07214_, _07213_, _02669_);
  not (_07215_, _07142_);
  and (_07216_, _07215_, _04982_);
  not (_07217_, _07216_);
  nor (_07218_, _07205_, _05332_);
  and (_07219_, _07218_, _07217_);
  nor (_07220_, _07219_, _07214_);
  nor (_07221_, _07220_, _03243_);
  or (_07222_, _07216_, _03244_);
  nor (_07223_, _07222_, _07158_);
  or (_07224_, _07223_, _02654_);
  nor (_07225_, _07224_, _07221_);
  nor (_07226_, _06078_, _07143_);
  nor (_07227_, _07226_, _07142_);
  and (_07228_, _07227_, _02654_);
  nor (_07229_, _07228_, _07225_);
  and (_07230_, _07229_, _05883_);
  nor (_07231_, _06087_, _07143_);
  nor (_07232_, _07231_, _07142_);
  nor (_07233_, _07232_, _05883_);
  or (_07234_, _07233_, _07230_);
  and (_07235_, _07234_, _03124_);
  nor (_07236_, _07155_, _03124_);
  or (_07237_, _07236_, _02650_);
  or (_07238_, _07237_, _07235_);
  nand (_07239_, _07174_, _02650_);
  and (_07240_, _07239_, _07238_);
  nor (_07241_, _07240_, _03121_);
  and (_07242_, _06131_, _04629_);
  nor (_07243_, _07242_, _07142_);
  and (_07244_, _07243_, _03121_);
  nor (_07245_, _07244_, _07241_);
  or (_07246_, _07245_, _27789_);
  or (_07247_, _27788_, \oc8051_golden_model_1.IE [7]);
  and (_07248_, _07247_, _27053_);
  and (_26417_, _07248_, _07246_);
  nand (_07249_, \oc8051_golden_model_1.DPH [7], _27053_);
  nor (_26418_, _07249_, _27788_);
  nand (_07250_, \oc8051_golden_model_1.DPL [7], _27053_);
  nor (_26419_, _07250_, _27788_);
  or (_07251_, _06086_, rst);
  nor (_26420_, _07251_, _27788_);
  nand (_07252_, \oc8051_golden_model_1.B [7], _27053_);
  nor (_26422_, _07252_, _27788_);
  not (_07253_, _03287_);
  and (_07254_, _02204_, _01959_);
  and (_07255_, _07254_, _01704_);
  and (_07256_, _05959_, _02204_);
  nor (_07257_, _07256_, _07255_);
  and (_07258_, _02204_, _02024_);
  not (_07259_, _07258_);
  and (_07260_, _07259_, _07257_);
  nor (_07261_, _07260_, _03452_);
  and (_07262_, _01966_, _03421_);
  and (_07263_, _03187_, _03417_);
  not (_07264_, _07263_);
  and (_07265_, _03176_, _02204_);
  and (_07266_, _03391_, _03150_);
  nor (_07267_, _01988_, _03417_);
  nor (_07268_, _07267_, _03407_);
  not (_07269_, _07268_);
  and (_07270_, _04505_, _02204_);
  and (_07271_, _03394_, _03421_);
  nor (_07272_, _07271_, _07270_);
  not (_07273_, _07272_);
  and (_07274_, _07270_, _03452_);
  nor (_07275_, _07274_, _04504_);
  and (_07276_, _07275_, _07273_);
  nor (_07277_, _07276_, _07269_);
  not (_07278_, _07277_);
  and (_07279_, _03394_, _02674_);
  nor (_07280_, _04545_, _07279_);
  nor (_07281_, _07280_, _03716_);
  nor (_07282_, _07281_, _07278_);
  and (_07283_, _02661_, _02204_);
  and (_07284_, _07283_, _02503_);
  nor (_07285_, _07284_, _03288_);
  and (_07286_, _07285_, _07282_);
  nor (_07287_, _07286_, _07266_);
  nor (_07288_, _01995_, _03417_);
  nor (_07289_, _07288_, _07287_);
  and (_07290_, _03162_, _02204_);
  and (_07291_, _07290_, _02503_);
  nor (_07292_, _07291_, _03422_);
  and (_07293_, _07292_, _07289_);
  and (_07294_, _03168_, _02204_);
  and (_07295_, _03167_, _02674_);
  and (_07296_, _07295_, _04485_);
  nor (_07297_, _07296_, _07294_);
  and (_07298_, _07297_, _07293_);
  and (_07299_, _07294_, _03452_);
  nor (_07300_, _07299_, _07298_);
  nor (_07301_, _07300_, _07265_);
  not (_07302_, _07301_);
  and (_07303_, _07302_, _03432_);
  or (_07304_, _07303_, _03187_);
  and (_07305_, _07304_, _07264_);
  and (_07306_, _03144_, _02204_);
  and (_07307_, _07306_, _03127_);
  nor (_07308_, _07307_, _07305_);
  nor (_07309_, _02000_, _03417_);
  and (_07310_, _03118_, _03421_);
  nor (_07311_, _07310_, _07309_);
  and (_07312_, _07311_, _07308_);
  and (_07313_, _04485_, _03119_);
  nor (_07314_, _07313_, _03300_);
  and (_07315_, _07314_, _07312_);
  nor (_07316_, _07315_, _03456_);
  nor (_07317_, _07316_, _02025_);
  and (_07318_, _02025_, _03417_);
  nor (_07319_, _07318_, _07317_);
  or (_07320_, _07319_, _07262_);
  nor (_07321_, _07320_, _07261_);
  and (_07322_, _01966_, _02674_);
  and (_07323_, _04485_, _07322_);
  not (_07324_, _07323_);
  and (_07325_, _07324_, _07321_);
  and (_07326_, _02575_, _02204_);
  and (_07327_, _07326_, _02503_);
  nor (_07328_, _07327_, _01967_);
  and (_07329_, _07328_, _07325_);
  and (_07330_, _01967_, _03417_);
  nor (_07331_, _07330_, _07329_);
  and (_07332_, _03251_, _02204_);
  and (_07333_, _02656_, _02204_);
  nor (_07334_, _07333_, _07332_);
  and (_07335_, _03243_, _02204_);
  and (_07336_, _02669_, _02204_);
  nor (_07337_, _07336_, _07335_);
  and (_07338_, _07337_, _07334_);
  nor (_07339_, _07338_, _03452_);
  nor (_07340_, _07339_, _01965_);
  not (_07341_, _07340_);
  nor (_07342_, _07341_, _07331_);
  and (_07343_, _01965_, _03417_);
  nor (_07344_, _07343_, _07342_);
  nand (_07345_, _03241_, _02204_);
  nor (_07346_, _07345_, _03452_);
  nor (_07347_, _07346_, _07344_);
  and (_07348_, _01970_, _03421_);
  and (_07349_, _01936_, \oc8051_golden_model_1.SP [0]);
  nor (_07350_, _07349_, _07348_);
  and (_07351_, _07350_, _07347_);
  and (_07352_, _03123_, _02204_);
  and (_07353_, _01970_, _02674_);
  and (_07354_, _04485_, _07353_);
  nor (_07355_, _07354_, _07352_);
  and (_07356_, _07355_, _07351_);
  and (_07357_, _07352_, _03452_);
  nor (_07358_, _07357_, _07356_);
  nor (_07359_, _06741_, _03417_);
  nor (_07360_, _07359_, _07358_);
  and (_07361_, _07360_, _07253_);
  nor (_07362_, _07361_, _03508_);
  and (_07363_, _01954_, _03421_);
  nor (_07364_, _07363_, _07362_);
  and (_07365_, _03121_, _02204_);
  and (_07366_, _05812_, _04485_);
  nor (_07367_, _07366_, _07365_);
  and (_07368_, _07367_, _07364_);
  and (_07369_, _07365_, _03452_);
  nor (_07370_, _07369_, _07368_);
  not (_07371_, _07370_);
  and (_07372_, _03521_, _02650_);
  and (_07373_, _03783_, _01936_);
  and (_07374_, _07326_, _04220_);
  and (_07375_, _03521_, _03150_);
  and (_07376_, _07283_, _04220_);
  not (_07377_, _03777_);
  or (_07378_, _07280_, _07377_);
  not (_07379_, _07283_);
  or (_07380_, _01767_, _02021_);
  nor (_07381_, _07380_, _01987_);
  nor (_07382_, _07381_, _07270_);
  and (_07383_, _07270_, _04220_);
  or (_07384_, _07383_, _04504_);
  or (_07385_, _07384_, _07382_);
  nor (_07386_, _07380_, _01994_);
  nor (_07387_, _03783_, _01988_);
  nor (_07388_, _07387_, _07386_);
  and (_07389_, _07388_, _07385_);
  and (_07390_, _07389_, _07379_);
  and (_07391_, _07390_, _07378_);
  nor (_07392_, _07391_, _07376_);
  nor (_07393_, _07392_, _03288_);
  nor (_07394_, _07393_, _07375_);
  nor (_07395_, _03783_, _01995_);
  nor (_07396_, _07395_, _07394_);
  and (_07397_, _07290_, _02471_);
  nor (_07398_, _07380_, _01989_);
  nor (_07399_, _07398_, _07397_);
  and (_07400_, _07399_, _07396_);
  and (_07401_, _07295_, _03777_);
  nor (_07402_, _07401_, _07294_);
  and (_07403_, _07402_, _07400_);
  and (_07404_, _07294_, _04220_);
  nor (_07405_, _07404_, _07403_);
  and (_07406_, _07265_, _02370_);
  or (_07407_, _07406_, _03187_);
  nor (_07408_, _07407_, _07405_);
  and (_07409_, _03783_, _03187_);
  nor (_07410_, _07409_, _07408_);
  and (_07411_, _07306_, _02370_);
  nor (_07412_, _07411_, _07410_);
  nor (_07413_, _03783_, _02000_);
  nor (_07414_, _07380_, _01992_);
  nor (_07415_, _07414_, _07413_);
  and (_07416_, _07415_, _07412_);
  and (_07417_, _03777_, _03119_);
  nor (_07418_, _07417_, _03300_);
  and (_07419_, _07418_, _07416_);
  nor (_07420_, _07419_, _03519_);
  nor (_07421_, _07420_, _02025_);
  and (_07422_, _03783_, _02025_);
  nor (_07423_, _07422_, _07421_);
  nor (_07424_, _07260_, _04220_);
  not (_07425_, _07380_);
  and (_07426_, _07425_, _01966_);
  or (_07427_, _07426_, _07424_);
  nor (_07428_, _07427_, _07423_);
  and (_07429_, _03777_, _07322_);
  nor (_07430_, _07429_, _07326_);
  and (_07431_, _07430_, _07428_);
  nor (_07432_, _07431_, _07374_);
  nor (_07433_, _07432_, _01967_);
  and (_07434_, _03783_, _01967_);
  nor (_07435_, _07434_, _07433_);
  nor (_07436_, _07338_, _04220_);
  nor (_07437_, _07436_, _01965_);
  not (_07438_, _07437_);
  nor (_07439_, _07438_, _07435_);
  and (_07440_, _03783_, _01965_);
  nor (_07441_, _07440_, _07439_);
  nor (_07442_, _07345_, _04220_);
  nor (_07443_, _07442_, _01936_);
  not (_07444_, _07443_);
  nor (_07445_, _07444_, _07441_);
  nor (_07446_, _07445_, _07373_);
  and (_07447_, _07425_, _01970_);
  nor (_07448_, _07447_, _07446_);
  and (_07449_, _03777_, _07353_);
  nor (_07450_, _07449_, _07352_);
  and (_07451_, _07450_, _07448_);
  and (_07452_, _07352_, _04220_);
  nor (_07453_, _07452_, _07451_);
  nor (_07454_, _06741_, _03783_);
  nor (_07455_, _07454_, _03287_);
  not (_07456_, _07455_);
  nor (_07457_, _07456_, _07453_);
  nor (_07458_, _07457_, _07372_);
  and (_07459_, _07425_, _01954_);
  nor (_07460_, _07459_, _07458_);
  and (_07461_, _05812_, _03777_);
  nor (_07462_, _07461_, _07365_);
  and (_07463_, _07462_, _07460_);
  and (_07464_, _07365_, _04220_);
  nor (_07465_, _07464_, _07463_);
  not (_07466_, _00001_);
  and (_07467_, _07255_, _01673_);
  not (_07468_, _07467_);
  nor (_07469_, _07256_, _03300_);
  nor (_07470_, _07365_, _07352_);
  and (_07471_, _07470_, _07469_);
  and (_07472_, _07471_, _07338_);
  and (_07473_, _07472_, _07468_);
  and (_07474_, _07345_, _03289_);
  and (_07475_, _07254_, _02023_);
  and (_07476_, _07254_, _01917_);
  nor (_07477_, _07476_, _07475_);
  and (_07478_, _07477_, _07474_);
  nor (_07479_, _07283_, _07270_);
  nor (_07480_, _07294_, _07290_);
  and (_07481_, _07480_, _07479_);
  nor (_07482_, _07306_, _07265_);
  not (_07483_, _07326_);
  nand (_07484_, _01917_, _01980_);
  nor (_07485_, _02576_, _07484_);
  not (_07486_, _01917_);
  or (_07487_, _02565_, _07486_);
  nor (_07488_, _07487_, _01989_);
  nor (_07489_, _07488_, _07485_);
  nand (_07490_, _01970_, _01928_);
  not (_07491_, _07490_);
  and (_07492_, _01992_, _01989_);
  nor (_07493_, _07492_, _01926_);
  nor (_07494_, _07493_, _07491_);
  and (_07495_, _07494_, _07489_);
  nor (_07496_, _06742_, _03548_);
  nor (_07497_, _04504_, _01936_);
  and (_07498_, _07497_, _06665_);
  and (_07499_, _07498_, _07496_);
  and (_07500_, _07499_, _07495_);
  nor (_07501_, _02634_, _03510_);
  nor (_07502_, _07501_, _05816_);
  and (_07503_, _01954_, _02636_);
  nor (_07504_, _02674_, _01920_);
  or (_07505_, _07504_, _01987_);
  not (_07506_, _07505_);
  nor (_07507_, _07506_, _07503_);
  nor (_07508_, _01992_, _01918_);
  and (_07509_, _03167_, _02640_);
  nor (_07510_, _07509_, _07508_);
  and (_07511_, _07510_, _07507_);
  and (_07512_, _07511_, _07502_);
  and (_07513_, _07512_, _07500_);
  and (_07514_, _02660_, _01917_);
  not (_07515_, _07514_);
  nor (_07516_, _01992_, _07484_);
  nor (_07517_, _07516_, _03119_);
  and (_07518_, _07517_, _07515_);
  nor (_07519_, _05812_, _04545_);
  nor (_07520_, _07295_, _07322_);
  and (_07521_, _07520_, _07519_);
  not (_07522_, _03546_);
  nor (_07523_, _03342_, _03187_);
  and (_07524_, _07523_, _07522_);
  and (_07525_, _07524_, _07521_);
  and (_07526_, _01995_, _01968_);
  and (_07527_, _01895_, _01833_);
  and (_07528_, _07527_, _01920_);
  nor (_07529_, _02576_, _01918_);
  nor (_07530_, _07529_, _07528_);
  and (_07531_, _01966_, _01920_);
  and (_07532_, _03394_, _01917_);
  nor (_07533_, _07532_, _07531_);
  and (_07534_, _07533_, _07530_);
  and (_07535_, _07534_, _07526_);
  and (_07536_, _07535_, _07525_);
  and (_07537_, _07536_, _07518_);
  and (_07538_, _07537_, _07513_);
  and (_07539_, _07538_, _07483_);
  and (_07540_, _07539_, _07482_);
  and (_07541_, _07540_, _07481_);
  and (_07542_, _07541_, _07478_);
  and (_07543_, _07542_, _07473_);
  nor (_07544_, _07543_, _07466_);
  not (_07545_, _07544_);
  nor (_07546_, _07545_, _07465_);
  and (_07547_, _07546_, _07371_);
  and (_07548_, _05812_, _03859_);
  and (_07549_, _03859_, _07353_);
  and (_07550_, _03859_, _07322_);
  and (_07551_, _03859_, _03119_);
  and (_07552_, _03782_, \oc8051_golden_model_1.SP [2]);
  or (_07553_, _07552_, \oc8051_golden_model_1.SP [3]);
  and (_07554_, _07553_, _06656_);
  not (_07555_, _07554_);
  nor (_07556_, _07555_, _02000_);
  and (_07557_, _07295_, _03859_);
  not (_07558_, _01995_);
  and (_07559_, _03288_, _02295_);
  and (_07560_, _04545_, _03859_);
  nor (_07561_, _07555_, _01988_);
  nor (_07562_, _07279_, \oc8051_golden_model_1.PSW [3]);
  and (_07563_, _07279_, _03859_);
  nor (_07564_, _07563_, _07562_);
  nor (_07565_, _07564_, _07270_);
  and (_07566_, _07270_, _03127_);
  nor (_07567_, _07566_, _04504_);
  not (_07568_, _07567_);
  nor (_07569_, _07568_, _07565_);
  or (_07570_, _07569_, _04545_);
  nor (_07571_, _07570_, _07561_);
  or (_07572_, _07571_, _07283_);
  nor (_07573_, _07572_, _07560_);
  and (_07574_, _07283_, _02405_);
  or (_07575_, _07574_, _03288_);
  nor (_07576_, _07575_, _07573_);
  nor (_07577_, _07576_, _07559_);
  nor (_07578_, _07577_, _07558_);
  nor (_07579_, _07554_, _01995_);
  nor (_07580_, _07579_, _07290_);
  not (_07581_, _07580_);
  nor (_07582_, _07581_, _07578_);
  and (_07583_, _07290_, _02405_);
  or (_07584_, _07583_, _07295_);
  nor (_07585_, _07584_, _07582_);
  or (_07586_, _07585_, _07294_);
  nor (_07587_, _07586_, _07557_);
  and (_07588_, _07294_, _02405_);
  or (_07589_, _07588_, _07265_);
  nor (_07590_, _07589_, _07587_);
  and (_07591_, _07265_, _02295_);
  nor (_07592_, _07591_, _07590_);
  and (_07593_, _07592_, _03430_);
  and (_07594_, _07554_, _03187_);
  nor (_07595_, _07594_, _07593_);
  nor (_07596_, _07595_, _07306_);
  and (_07597_, _07306_, _03133_);
  or (_07598_, _07597_, _07596_);
  and (_07599_, _07598_, _02000_);
  or (_07600_, _07599_, _03119_);
  nor (_07601_, _07600_, _07556_);
  or (_07602_, _07601_, _03300_);
  nor (_07603_, _07602_, _07551_);
  and (_07604_, _03300_, _03909_);
  nor (_07605_, _07604_, _07603_);
  nor (_07606_, _07605_, _02025_);
  and (_07607_, _07554_, _02025_);
  not (_07608_, _07607_);
  and (_07609_, _07608_, _07260_);
  not (_07610_, _07609_);
  nor (_07611_, _07610_, _07606_);
  nor (_07612_, _07260_, _02405_);
  nor (_07613_, _07612_, _07611_);
  nor (_07614_, _07613_, _07322_);
  or (_07615_, _07614_, _07326_);
  nor (_07616_, _07615_, _07550_);
  and (_07617_, _03391_, _02575_);
  nor (_07618_, _07617_, _07616_);
  nor (_07619_, _07618_, _01967_);
  and (_07620_, _07554_, _01967_);
  not (_07621_, _07620_);
  and (_07622_, _07621_, _07338_);
  not (_07623_, _07622_);
  nor (_07624_, _07623_, _07619_);
  nor (_07625_, _07338_, _02405_);
  nor (_07626_, _07625_, _01965_);
  not (_07627_, _07626_);
  nor (_07628_, _07627_, _07624_);
  and (_07629_, _07554_, _01965_);
  not (_07630_, _07629_);
  and (_07631_, _07630_, _07345_);
  not (_07632_, _07631_);
  nor (_07633_, _07632_, _07628_);
  nor (_07634_, _07345_, _02405_);
  nor (_07635_, _07634_, _01936_);
  not (_07636_, _07635_);
  nor (_07637_, _07636_, _07633_);
  and (_07638_, _07554_, _01936_);
  nor (_07639_, _07638_, _07353_);
  not (_07640_, _07639_);
  nor (_07641_, _07640_, _07637_);
  or (_07642_, _07641_, _07352_);
  nor (_07643_, _07642_, _07549_);
  and (_07644_, _07352_, _02405_);
  nor (_07645_, _07644_, _06742_);
  not (_07646_, _07645_);
  nor (_07647_, _07646_, _07643_);
  nor (_07648_, _07554_, _06741_);
  nor (_07649_, _07648_, _03287_);
  not (_07650_, _07649_);
  nor (_07651_, _07650_, _07647_);
  and (_07652_, _03287_, _03909_);
  or (_07653_, _07652_, _05812_);
  nor (_07654_, _07653_, _07651_);
  or (_07655_, _07654_, _07365_);
  nor (_07656_, _07655_, _07548_);
  and (_07657_, _07365_, _02405_);
  nor (_07658_, _07657_, _07656_);
  and (_07659_, _07365_, _04123_);
  and (_07660_, _01954_, _01917_);
  and (_07661_, _03303_, _02650_);
  nor (_07662_, _03782_, \oc8051_golden_model_1.SP [2]);
  nor (_07663_, _07662_, _07552_);
  and (_07664_, _07663_, _01936_);
  and (_07665_, _07326_, _04123_);
  nor (_07666_, _07663_, _02000_);
  nor (_07667_, _07666_, _05172_);
  and (_07668_, _03303_, _03150_);
  and (_07669_, _07283_, _04123_);
  not (_07670_, _03644_);
  or (_07671_, _07280_, _07670_);
  and (_07672_, _07270_, _04123_);
  or (_07673_, _07672_, _04504_);
  nor (_07674_, _07270_, _07532_);
  or (_07675_, _07674_, _07673_);
  nor (_07676_, _07663_, _01988_);
  nor (_07677_, _07676_, _07514_);
  and (_07678_, _07677_, _07675_);
  and (_07679_, _07678_, _07379_);
  and (_07680_, _07679_, _07671_);
  nor (_07681_, _07680_, _07669_);
  nor (_07682_, _07681_, _03288_);
  nor (_07683_, _07682_, _07668_);
  nor (_07684_, _07663_, _01995_);
  nor (_07685_, _07684_, _07683_);
  and (_07686_, _03167_, _01917_);
  and (_07687_, _07290_, _02439_);
  nor (_07688_, _07687_, _07686_);
  and (_07689_, _07688_, _07685_);
  and (_07690_, _07295_, _03644_);
  nor (_07691_, _07690_, _07294_);
  and (_07692_, _07691_, _07689_);
  and (_07693_, _07294_, _04123_);
  nor (_07694_, _07693_, _07692_);
  and (_07695_, _07265_, _02333_);
  nor (_07696_, _07695_, _07694_);
  and (_07697_, _07696_, _03430_);
  and (_07698_, _07663_, _03187_);
  nor (_07699_, _07698_, _07697_);
  and (_07700_, _07306_, _02333_);
  nor (_07701_, _07700_, _07699_);
  and (_07702_, _07701_, _07667_);
  and (_07703_, _03644_, _03119_);
  nor (_07704_, _07703_, _03300_);
  and (_07705_, _07704_, _07702_);
  nor (_07706_, _07705_, _03301_);
  nor (_07707_, _07706_, _02025_);
  and (_07708_, _07663_, _02025_);
  nor (_07709_, _07708_, _07707_);
  and (_07710_, _01966_, _01917_);
  nor (_07711_, _07260_, _04123_);
  nor (_07712_, _07711_, _07710_);
  not (_07713_, _07712_);
  nor (_07714_, _07713_, _07709_);
  and (_07715_, _03644_, _07322_);
  nor (_07716_, _07715_, _07326_);
  and (_07717_, _07716_, _07714_);
  nor (_07718_, _07717_, _07665_);
  nor (_07719_, _07718_, _01967_);
  and (_07720_, _07663_, _01967_);
  nor (_07721_, _07720_, _07719_);
  nor (_07722_, _07338_, _04123_);
  nor (_07723_, _07722_, _01965_);
  not (_07724_, _07723_);
  nor (_07725_, _07724_, _07721_);
  and (_07726_, _07663_, _01965_);
  nor (_07727_, _07726_, _07725_);
  nor (_07728_, _07345_, _04123_);
  nor (_07729_, _07728_, _01936_);
  not (_07730_, _07729_);
  nor (_07731_, _07730_, _07727_);
  nor (_07732_, _07731_, _07664_);
  nor (_07733_, _07732_, _03547_);
  and (_07734_, _03644_, _07353_);
  nor (_07735_, _07734_, _07352_);
  and (_07736_, _07735_, _07733_);
  and (_07737_, _07352_, _04123_);
  nor (_07738_, _07737_, _07736_);
  nor (_07739_, _07663_, _06741_);
  nor (_07740_, _07739_, _07738_);
  and (_07741_, _07740_, _07253_);
  nor (_07742_, _07741_, _07661_);
  nor (_07743_, _07742_, _07660_);
  and (_07744_, _05812_, _03644_);
  nor (_07745_, _07744_, _07365_);
  and (_07746_, _07745_, _07743_);
  nor (_07747_, _07746_, _07659_);
  nor (_07748_, _07747_, _07545_);
  not (_07749_, _07748_);
  nor (_07750_, _07749_, _07658_);
  and (_07751_, _07750_, _07547_);
  or (_07752_, _07751_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_07753_, _06741_, _06665_);
  and (_07754_, _07753_, _07497_);
  and (_07755_, _07754_, _07526_);
  nor (_07756_, _07755_, _07466_);
  and (_07757_, _07756_, \oc8051_golden_model_1.SP [0]);
  and (_07758_, _07757_, _03565_);
  and (_07759_, \oc8051_golden_model_1.SP [1], _03417_);
  and (_07760_, _07759_, \oc8051_golden_model_1.SP [2]);
  nor (_07761_, _07759_, _07663_);
  nor (_07762_, _07761_, _07760_);
  and (_07763_, _06623_, _03417_);
  nor (_07764_, _07760_, _07554_);
  nor (_07765_, _07764_, _07763_);
  and (_07766_, _07765_, _07756_);
  and (_07767_, _07766_, _07762_);
  and (_07768_, _07767_, _07758_);
  not (_07769_, _07768_);
  and (_07770_, _07769_, _07752_);
  not (_07771_, _07465_);
  nor (_07772_, _07545_, _07370_);
  and (_07773_, _07772_, _07771_);
  not (_07774_, _07747_);
  nor (_07775_, _07658_, _07545_);
  and (_07776_, _07775_, _07774_);
  nand (_07777_, _07776_, _07773_);
  and (_07778_, _07365_, _06131_);
  and (_07779_, _04218_, _04268_);
  and (_07780_, _07779_, _04170_);
  and (_07781_, _07780_, _04120_);
  and (_07782_, _07781_, _04012_);
  and (_07783_, _07782_, _03904_);
  and (_07784_, _07783_, _03960_);
  nor (_07785_, _07784_, _04069_);
  and (_07786_, _07784_, _04069_);
  nor (_07787_, _07786_, _07785_);
  and (_07788_, _07787_, _05812_);
  not (_07789_, _07335_);
  and (_07790_, _07336_, _06079_);
  not (_07791_, _02025_);
  not (_07792_, _03300_);
  nor (_07793_, _06533_, _07792_);
  not (_07794_, _07265_);
  or (_07795_, _06521_, _07794_);
  not (_07796_, _03288_);
  or (_07797_, _06496_, _07796_);
  not (_07798_, _04545_);
  or (_07799_, _07798_, _04067_);
  not (_07800_, _04426_);
  and (_07801_, _03777_, _04485_);
  and (_07802_, _07801_, _04535_);
  and (_07803_, _07802_, _04531_);
  and (_07804_, _07803_, _04373_);
  or (_07805_, _07804_, _07800_);
  nand (_07806_, _07804_, _07800_);
  and (_07807_, _07806_, _07805_);
  and (_07808_, _07807_, _03406_);
  and (_07809_, _01988_, \oc8051_golden_model_1.ACC [7]);
  nor (_07810_, _02260_, _01988_);
  or (_07811_, _07810_, _07809_);
  and (_07812_, _07811_, _04539_);
  or (_07813_, _07812_, _04545_);
  or (_07814_, _07813_, _07808_);
  and (_07815_, _07814_, _07799_);
  or (_07816_, _07815_, _07283_);
  nand (_07817_, _07283_, _05927_);
  and (_07818_, _07817_, _07816_);
  or (_07819_, _07818_, _03288_);
  and (_07820_, _07819_, _07797_);
  or (_07821_, _07820_, _07558_);
  nor (_07822_, _02259_, _01995_);
  nor (_07823_, _07822_, _07290_);
  and (_07824_, _07823_, _07821_);
  and (_07825_, _07290_, _07800_);
  or (_07826_, _07825_, _07265_);
  or (_07827_, _07826_, _07824_);
  and (_07828_, _07827_, _07795_);
  or (_07829_, _07828_, _03187_);
  not (_07830_, _07306_);
  nand (_07831_, _05060_, _03187_);
  and (_07832_, _07831_, _07830_);
  and (_07833_, _07832_, _07829_);
  nand (_07834_, _07306_, _06496_);
  nor (_07835_, _07834_, _06494_);
  or (_07836_, _07835_, _07833_);
  and (_07837_, _07836_, _02000_);
  nor (_07838_, _02260_, _02000_);
  or (_07839_, _07838_, _03200_);
  or (_07840_, _07839_, _07837_);
  nand (_07841_, _05060_, _03200_);
  and (_07842_, _07841_, _07840_);
  or (_07843_, _07842_, _03119_);
  and (_07844_, _05059_, _03119_);
  nand (_07845_, _07844_, _04070_);
  and (_07846_, _07845_, _07792_);
  and (_07847_, _07846_, _07843_);
  or (_07848_, _07847_, _07793_);
  and (_07849_, _07848_, _07791_);
  and (_07850_, _02259_, _02025_);
  or (_07851_, _07850_, _07255_);
  or (_07852_, _07851_, _07849_);
  nand (_07853_, _07255_, _04426_);
  and (_07854_, _07853_, _07852_);
  or (_07855_, _07854_, _07256_);
  not (_07856_, _07256_);
  or (_07857_, _07856_, _04067_);
  and (_07858_, _07857_, _07259_);
  and (_07859_, _07858_, _07855_);
  nor (_07860_, _07259_, _06070_);
  or (_07861_, _07860_, _02577_);
  or (_07862_, _07861_, _07859_);
  and (_07863_, _02577_, _02204_);
  nor (_07864_, _07863_, _07326_);
  and (_07865_, _07864_, _07862_);
  and (_07866_, _07326_, _05889_);
  or (_07867_, _07866_, _01967_);
  or (_07868_, _07867_, _07865_);
  and (_07869_, _02260_, _01967_);
  nor (_07870_, _07869_, _07333_);
  and (_07871_, _07870_, _07868_);
  nor (_07872_, _07332_, _06080_);
  nor (_07873_, _07872_, _07334_);
  or (_07874_, _07873_, _07871_);
  not (_07875_, _07336_);
  not (_07876_, _07332_);
  or (_07877_, _07876_, _06089_);
  and (_07878_, _07877_, _07875_);
  and (_07879_, _07878_, _07874_);
  or (_07880_, _07879_, _07790_);
  and (_07881_, _07880_, _07789_);
  and (_07882_, _07335_, _06088_);
  or (_07883_, _07882_, _01965_);
  or (_07884_, _07883_, _07881_);
  and (_07885_, _02654_, _02204_);
  and (_07886_, _02260_, _01965_);
  nor (_07887_, _07886_, _07885_);
  and (_07888_, _07887_, _07884_);
  and (_07889_, _03239_, _02204_);
  not (_07890_, _07889_);
  and (_07891_, _07890_, _06078_);
  nor (_07892_, _07891_, _07345_);
  or (_07893_, _07892_, _07888_);
  nand (_07894_, _07889_, _06087_);
  and (_07895_, _07894_, _05408_);
  and (_07896_, _07895_, _07893_);
  and (_07897_, _02259_, _01936_);
  nand (_07898_, _01970_, _01704_);
  not (_07899_, _07898_);
  or (_07900_, _07899_, _07897_);
  or (_07901_, _07900_, _07896_);
  or (_07902_, _07898_, _07807_);
  and (_07903_, _07902_, _07901_);
  or (_07904_, _07903_, _07353_);
  not (_07905_, _07352_);
  not (_07906_, _07353_);
  and (_07907_, _04221_, _04270_);
  and (_07908_, _07907_, _04168_);
  and (_07909_, _07908_, _04118_);
  and (_07910_, _07909_, _04014_);
  and (_07911_, _07910_, _03906_);
  and (_07912_, _07911_, _03958_);
  nor (_07913_, _07912_, _04069_);
  and (_07914_, _07912_, _04069_);
  or (_07915_, _07914_, _07913_);
  or (_07916_, _07915_, _07906_);
  and (_07917_, _07916_, _07905_);
  and (_07918_, _07917_, _07904_);
  nor (_07919_, _07905_, _05927_);
  or (_07920_, _07919_, _02646_);
  or (_07921_, _07920_, _07918_);
  nand (_07922_, _02801_, _02646_);
  and (_07923_, _07922_, _07921_);
  or (_07924_, _07923_, _01971_);
  and (_07925_, _02260_, _01971_);
  nor (_07926_, _07925_, _03287_);
  and (_07927_, _07926_, _07924_);
  not (_07928_, _05822_);
  and (_07929_, _06530_, _03287_);
  nor (_07930_, _07929_, _07928_);
  not (_07931_, _07930_);
  nor (_07932_, _07931_, _07927_);
  not (_07933_, _04373_);
  not (_07934_, _04480_);
  not (_07935_, _04325_);
  not (_07936_, _03859_);
  nor (_07937_, _03777_, _04485_);
  and (_07938_, _07937_, _07670_);
  and (_07939_, _07938_, _07936_);
  and (_07940_, _07939_, _07935_);
  and (_07941_, _07940_, _07934_);
  and (_07942_, _07941_, _07933_);
  nor (_07943_, _07942_, _04426_);
  and (_07944_, _07942_, _04426_);
  or (_07945_, _07944_, _07943_);
  nor (_07946_, _07945_, _05822_);
  nor (_07947_, _07946_, _07932_);
  nor (_07948_, _07947_, _05812_);
  or (_07949_, _07948_, _07365_);
  nor (_07950_, _07949_, _07788_);
  nor (_07951_, _07950_, _07778_);
  nor (_07952_, _07951_, _07545_);
  or (_07953_, _07952_, _07777_);
  and (_07954_, _07953_, _07770_);
  and (_07955_, _05786_, _02555_);
  and (_07956_, _02646_, _02596_);
  or (_07957_, _07956_, _07955_);
  and (_07958_, _07957_, _07756_);
  and (_07959_, _07958_, _07768_);
  or (_30758_[7], _07959_, _07954_);
  nor (_07960_, _07772_, _07546_);
  nor (_07961_, _07775_, _07748_);
  and (_07962_, _07961_, _07960_);
  and (_07963_, _07962_, _07544_);
  not (_07964_, _07963_);
  nand (_07965_, _01971_, _01647_);
  and (_07966_, _04888_, _05996_);
  nor (_07967_, _04888_, _05996_);
  nor (_07968_, _07967_, _07966_);
  and (_07969_, _07968_, _07333_);
  not (_07970_, _07255_);
  or (_07971_, _07970_, _03716_);
  and (_07972_, _04268_, _02204_);
  nand (_07973_, _05108_, _03119_);
  or (_07974_, _07973_, _07972_);
  and (_07975_, _07290_, _03716_);
  nor (_07976_, _07379_, _04888_);
  or (_07977_, _04485_, _04539_);
  nor (_07978_, _01988_, _01647_);
  and (_07979_, _01988_, \oc8051_golden_model_1.ACC [0]);
  or (_07980_, _07979_, _07978_);
  nor (_07981_, _07980_, _03406_);
  nor (_07982_, _07981_, _07283_);
  and (_07983_, _07982_, _07977_);
  or (_07984_, _07983_, _07976_);
  and (_07985_, _07984_, _07796_);
  and (_07986_, _05446_, \oc8051_golden_model_1.P3 [0]);
  nor (_07987_, _07986_, _05550_);
  and (_07988_, _07987_, _05543_);
  and (_07989_, _05444_, \oc8051_golden_model_1.P1 [0]);
  and (_07990_, _05436_, \oc8051_golden_model_1.P2 [0]);
  and (_07991_, _04552_, \oc8051_golden_model_1.P0 [0]);
  or (_07992_, _07991_, _07990_);
  nor (_07993_, _07992_, _07989_);
  and (_07994_, _07993_, _05540_);
  and (_07995_, _07994_, _07988_);
  and (_07996_, _07995_, _04836_);
  nand (_07997_, _07996_, _05533_);
  and (_07998_, _07997_, _03288_);
  or (_07999_, _07998_, _07558_);
  or (_08000_, _07999_, _07985_);
  nor (_08001_, _01995_, \oc8051_golden_model_1.PC [0]);
  nor (_08002_, _08001_, _07290_);
  and (_08003_, _08002_, _08000_);
  or (_08004_, _08003_, _07975_);
  and (_08005_, _08004_, _07794_);
  or (_08006_, _04633_, _07794_);
  nor (_08007_, _08006_, _07996_);
  or (_08008_, _08007_, _03187_);
  or (_08009_, _08008_, _08005_);
  nand (_08010_, _05109_, _03187_);
  and (_08011_, _08010_, _07830_);
  and (_08012_, _08011_, _08009_);
  or (_08013_, _07996_, _05533_);
  and (_08014_, _07997_, _07306_);
  and (_08015_, _08014_, _08013_);
  or (_08016_, _08015_, _08012_);
  and (_08017_, _08016_, _02000_);
  nor (_08018_, _02000_, _01647_);
  nor (_08019_, _05818_, _01992_);
  or (_08020_, _08019_, _08018_);
  or (_08021_, _08020_, _08017_);
  and (_08022_, _03118_, _02640_);
  not (_08023_, _08022_);
  nand (_08024_, _08019_, _05109_);
  and (_08025_, _08024_, _08023_);
  and (_08026_, _08025_, _08021_);
  nor (_08027_, _05109_, _08023_);
  or (_08028_, _08027_, _03119_);
  or (_08029_, _08028_, _08026_);
  and (_08030_, _08029_, _07974_);
  or (_08031_, _08030_, _03300_);
  nor (_08032_, _05556_, _04633_);
  and (_08033_, _04568_, \oc8051_golden_model_1.PSW [7]);
  and (_08034_, _08033_, _02439_);
  nor (_08035_, _08034_, _08032_);
  nand (_08036_, _08035_, _03300_);
  and (_08037_, _08036_, _07791_);
  and (_08038_, _08037_, _08031_);
  and (_08039_, _02025_, \oc8051_golden_model_1.PC [0]);
  or (_08040_, _07255_, _08039_);
  or (_08041_, _08040_, _08038_);
  and (_08042_, _08041_, _07971_);
  or (_08043_, _08042_, _07256_);
  or (_08044_, _07856_, _04268_);
  and (_08045_, _08044_, _07259_);
  and (_08046_, _08045_, _08043_);
  and (_08047_, _03716_, _02752_);
  and (_08048_, _06002_, \oc8051_golden_model_1.SCON [0]);
  not (_08049_, _08048_);
  and (_08050_, _05994_, \oc8051_golden_model_1.TCON [0]);
  and (_08051_, _06004_, \oc8051_golden_model_1.SBUF [0]);
  nor (_08052_, _08051_, _08050_);
  and (_08053_, _08052_, _08049_);
  and (_08054_, _05999_, \oc8051_golden_model_1.TMOD [0]);
  and (_08055_, _05977_, \oc8051_golden_model_1.P1INREG [0]);
  nor (_08056_, _08055_, _08054_);
  and (_08057_, _05982_, \oc8051_golden_model_1.P0INREG [0]);
  and (_08058_, _05989_, \oc8051_golden_model_1.TL0 [0]);
  nor (_08059_, _08058_, _08057_);
  and (_08060_, _08059_, _08056_);
  and (_08061_, _08060_, _08053_);
  and (_08062_, _06013_, \oc8051_golden_model_1.PCON [0]);
  and (_08063_, _06015_, \oc8051_golden_model_1.DPH [0]);
  nor (_08064_, _08063_, _08062_);
  and (_08065_, _08064_, _08061_);
  and (_08066_, _06027_, \oc8051_golden_model_1.TL1 [0]);
  not (_08067_, _08066_);
  and (_08068_, _06061_, \oc8051_golden_model_1.DPL [0]);
  and (_08069_, _06020_, \oc8051_golden_model_1.SP [0]);
  nor (_08070_, _08069_, _08068_);
  and (_08071_, _08070_, _08067_);
  and (_08072_, _06039_, \oc8051_golden_model_1.P2INREG [0]);
  not (_08073_, _08072_);
  and (_08074_, _06033_, \oc8051_golden_model_1.P3INREG [0]);
  and (_08075_, _06050_, \oc8051_golden_model_1.B [0]);
  nor (_08076_, _08075_, _08074_);
  and (_08077_, _08076_, _08073_);
  and (_08078_, _06053_, \oc8051_golden_model_1.IE [0]);
  and (_08079_, _06056_, \oc8051_golden_model_1.PSW [0]);
  nor (_08080_, _08079_, _08078_);
  and (_08081_, _06041_, \oc8051_golden_model_1.IP [0]);
  and (_08082_, _06047_, \oc8051_golden_model_1.ACC [0]);
  nor (_08083_, _08082_, _08081_);
  and (_08084_, _08083_, _08080_);
  and (_08085_, _08084_, _08077_);
  and (_08086_, _06025_, \oc8051_golden_model_1.TH1 [0]);
  and (_08087_, _06063_, \oc8051_golden_model_1.TH0 [0]);
  nor (_08088_, _08087_, _08086_);
  and (_08089_, _08088_, _08085_);
  and (_08090_, _08089_, _08071_);
  and (_08091_, _08090_, _08065_);
  not (_08092_, _08091_);
  nor (_08093_, _08092_, _08047_);
  nor (_08094_, _08093_, _07259_);
  or (_08095_, _08094_, _02577_);
  or (_08096_, _08095_, _08046_);
  and (_08097_, _02577_, _02503_);
  nor (_08098_, _08097_, _07326_);
  and (_08099_, _08098_, _08096_);
  and (_08100_, _07326_, _05996_);
  or (_08101_, _08100_, _01967_);
  or (_08102_, _08101_, _08099_);
  and (_08103_, _01967_, _01647_);
  nor (_08104_, _08103_, _07333_);
  and (_08105_, _08104_, _08102_);
  or (_08106_, _08105_, _07969_);
  and (_08107_, _08106_, _07876_);
  and (_08108_, _04888_, \oc8051_golden_model_1.ACC [0]);
  nor (_08109_, _04888_, \oc8051_golden_model_1.ACC [0]);
  nor (_08110_, _08109_, _08108_);
  and (_08111_, _08110_, _07332_);
  or (_08112_, _08111_, _08107_);
  and (_08113_, _08112_, _07875_);
  and (_08114_, _07966_, _07336_);
  or (_08115_, _08114_, _07335_);
  or (_08116_, _08115_, _08113_);
  or (_08117_, _08108_, _07789_);
  and (_08118_, _08117_, _08116_);
  or (_08119_, _08118_, _01965_);
  and (_08120_, _01965_, _01647_);
  nor (_08121_, _08120_, _07885_);
  and (_08122_, _08121_, _08119_);
  and (_08123_, _07967_, _07890_);
  nor (_08124_, _08123_, _07345_);
  or (_08125_, _08124_, _08122_);
  nand (_08126_, _08109_, _07889_);
  and (_08127_, _08126_, _08125_);
  or (_08128_, _08127_, _01936_);
  nand (_08129_, _01936_, _01647_);
  and (_08130_, _08129_, _07898_);
  and (_08131_, _08130_, _08128_);
  and (_08132_, _07899_, _04485_);
  or (_08133_, _08132_, _07353_);
  or (_08134_, _08133_, _08131_);
  or (_08135_, _04270_, _07906_);
  and (_08136_, _08135_, _08134_);
  or (_08137_, _08136_, _07352_);
  nand (_08138_, _07352_, _04888_);
  and (_08139_, _08138_, _05786_);
  and (_08140_, _08139_, _08137_);
  and (_08141_, _02646_, _01647_);
  or (_08142_, _08141_, _01971_);
  or (_08143_, _08142_, _08140_);
  and (_08144_, _08143_, _07965_);
  or (_08145_, _08144_, _03287_);
  or (_08146_, _08032_, _07253_);
  and (_08147_, _08146_, _05822_);
  and (_08148_, _08147_, _08145_);
  and (_08149_, _07928_, _04485_);
  or (_08150_, _08149_, _08148_);
  and (_08151_, _08150_, _05814_);
  and (_08152_, _05812_, _04270_);
  or (_08153_, _08152_, _07365_);
  or (_08154_, _08153_, _08151_);
  nand (_08155_, _07365_, _04888_);
  and (_08156_, _08155_, _07544_);
  and (_08157_, _08156_, _08154_);
  or (_08158_, _08157_, _07964_);
  and (_08159_, _07762_, _07756_);
  nor (_08160_, _07766_, _08159_);
  and (_08161_, _08160_, _07756_);
  and (_08162_, _08161_, _07759_);
  not (_08163_, _08162_);
  or (_08164_, _07963_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_08165_, _08164_, _08163_);
  and (_08166_, _08165_, _08158_);
  nor (_08167_, _02646_, _02529_);
  and (_08168_, _03073_, _02646_);
  or (_08169_, _08168_, _08167_);
  and (_08170_, _08169_, _08162_);
  or (_30702_, _08170_, _08166_);
  or (_08172_, _07963_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_08173_, _08172_, _08163_);
  nor (_08174_, _07937_, _07801_);
  and (_08175_, _08174_, _07928_);
  and (_08176_, _01970_, _02636_);
  nor (_08177_, _08176_, _03350_);
  and (_08178_, _01970_, _03339_);
  not (_08179_, _08178_);
  and (_08180_, _08179_, _08177_);
  not (_08181_, _08180_);
  nand (_08182_, _08181_, _08174_);
  and (_08183_, _04835_, _03016_);
  nor (_08184_, _04835_, _03016_);
  nor (_08185_, _08184_, _08183_);
  and (_08186_, _08185_, _07333_);
  nand (_08187_, _07255_, _03777_);
  nand (_08188_, _05036_, _03200_);
  and (_08189_, _05446_, \oc8051_golden_model_1.P3 [1]);
  nor (_08190_, _08189_, _05471_);
  and (_08191_, _08190_, _05464_);
  and (_08192_, _05444_, \oc8051_golden_model_1.P1 [1]);
  and (_08193_, _05436_, \oc8051_golden_model_1.P2 [1]);
  and (_08194_, _04552_, \oc8051_golden_model_1.P0 [1]);
  or (_08195_, _08194_, _08193_);
  nor (_08196_, _08195_, _08192_);
  and (_08197_, _08196_, _05461_);
  and (_08198_, _08197_, _08191_);
  and (_08199_, _08198_, _04790_);
  nor (_08200_, _08199_, _04563_);
  or (_08201_, _08200_, _07794_);
  nor (_08202_, _08174_, _04539_);
  nor (_08203_, _01988_, \oc8051_golden_model_1.PC [1]);
  and (_08204_, _01988_, \oc8051_golden_model_1.ACC [1]);
  or (_08205_, _08204_, _08203_);
  and (_08206_, _08205_, _04539_);
  or (_08207_, _08206_, _07283_);
  or (_08208_, _08207_, _08202_);
  nor (_08209_, _06123_, _05917_);
  nand (_08210_, _08209_, _07283_);
  and (_08211_, _08210_, _08208_);
  or (_08212_, _08211_, _03288_);
  nand (_08213_, _08199_, _05454_);
  or (_08214_, _08213_, _07796_);
  and (_08215_, _08214_, _08212_);
  or (_08216_, _08215_, _07558_);
  nor (_08217_, _01995_, _01620_);
  nor (_08218_, _08217_, _07290_);
  and (_08219_, _08218_, _08216_);
  and (_08220_, _07290_, _07377_);
  or (_08221_, _08220_, _07265_);
  or (_08222_, _08221_, _08219_);
  and (_08223_, _08222_, _08201_);
  or (_08224_, _08223_, _03187_);
  nand (_08225_, _05036_, _03187_);
  and (_08226_, _08225_, _07830_);
  and (_08227_, _08226_, _08224_);
  or (_08228_, _08199_, _05454_);
  and (_08229_, _08213_, _08228_);
  and (_08230_, _08229_, _07306_);
  or (_08231_, _08230_, _08227_);
  and (_08232_, _08231_, _02000_);
  nor (_08233_, _02000_, \oc8051_golden_model_1.PC [1]);
  or (_08234_, _03200_, _08233_);
  or (_08235_, _08234_, _08232_);
  and (_08236_, _08235_, _08188_);
  or (_08237_, _08236_, _03119_);
  and (_08238_, _04218_, _02204_);
  nand (_08239_, _05035_, _03119_);
  or (_08240_, _08239_, _08238_);
  and (_08241_, _08240_, _08237_);
  or (_08242_, _08241_, _03300_);
  nor (_08243_, _05477_, _04563_);
  and (_08244_, _04562_, \oc8051_golden_model_1.PSW [7]);
  and (_08245_, _08244_, _02439_);
  nor (_08246_, _08245_, _08243_);
  nand (_08247_, _08246_, _03300_);
  and (_08248_, _08247_, _07791_);
  and (_08249_, _08248_, _08242_);
  and (_08250_, _02025_, _01620_);
  or (_08251_, _07255_, _08250_);
  or (_08252_, _08251_, _08249_);
  and (_08253_, _08252_, _08187_);
  or (_08254_, _08253_, _07256_);
  or (_08255_, _07856_, _04218_);
  and (_08256_, _08255_, _07259_);
  and (_08257_, _08256_, _08254_);
  nor (_08258_, _03777_, _05889_);
  and (_08259_, _05982_, \oc8051_golden_model_1.P0INREG [1]);
  not (_08260_, _08259_);
  and (_08261_, _05994_, \oc8051_golden_model_1.TCON [1]);
  and (_08262_, _05999_, \oc8051_golden_model_1.TMOD [1]);
  nor (_08263_, _08262_, _08261_);
  and (_08264_, _08263_, _08260_);
  and (_08265_, _05989_, \oc8051_golden_model_1.TL0 [1]);
  and (_08266_, _06002_, \oc8051_golden_model_1.SCON [1]);
  nor (_08267_, _08266_, _08265_);
  and (_08269_, _05977_, \oc8051_golden_model_1.P1INREG [1]);
  and (_08270_, _06004_, \oc8051_golden_model_1.SBUF [1]);
  nor (_08272_, _08270_, _08269_);
  and (_08273_, _08272_, _08267_);
  and (_08275_, _08273_, _08264_);
  and (_08276_, _06013_, \oc8051_golden_model_1.PCON [1]);
  and (_08278_, _06015_, \oc8051_golden_model_1.DPH [1]);
  nor (_08279_, _08278_, _08276_);
  and (_08280_, _08279_, _08275_);
  and (_08281_, _06020_, \oc8051_golden_model_1.SP [1]);
  not (_08282_, _08281_);
  and (_08283_, _06061_, \oc8051_golden_model_1.DPL [1]);
  and (_08284_, _06063_, \oc8051_golden_model_1.TH0 [1]);
  nor (_08285_, _08284_, _08283_);
  and (_08286_, _08285_, _08282_);
  and (_08287_, _06047_, \oc8051_golden_model_1.ACC [1]);
  and (_08288_, _06039_, \oc8051_golden_model_1.P2INREG [1]);
  and (_08289_, _06033_, \oc8051_golden_model_1.P3INREG [1]);
  or (_08290_, _08289_, _08288_);
  or (_08291_, _08290_, _08287_);
  and (_08292_, _06041_, \oc8051_golden_model_1.IP [1]);
  and (_08293_, _06056_, \oc8051_golden_model_1.PSW [1]);
  nor (_08294_, _08293_, _08292_);
  and (_08295_, _06053_, \oc8051_golden_model_1.IE [1]);
  and (_08296_, _06050_, \oc8051_golden_model_1.B [1]);
  nor (_08297_, _08296_, _08295_);
  nand (_08298_, _08297_, _08294_);
  nor (_08299_, _08298_, _08291_);
  and (_08300_, _06025_, \oc8051_golden_model_1.TH1 [1]);
  and (_08301_, _06027_, \oc8051_golden_model_1.TL1 [1]);
  nor (_08302_, _08301_, _08300_);
  and (_08303_, _08302_, _08299_);
  and (_08304_, _08303_, _08286_);
  and (_08305_, _08304_, _08280_);
  not (_08306_, _08305_);
  nor (_08307_, _08306_, _08258_);
  nor (_08308_, _08307_, _07259_);
  or (_08309_, _08308_, _02577_);
  or (_08310_, _08309_, _08257_);
  and (_08311_, _02577_, _02471_);
  nor (_08312_, _08311_, _07326_);
  and (_08313_, _08312_, _08310_);
  and (_08314_, _07326_, _05984_);
  or (_08315_, _08314_, _01967_);
  or (_08316_, _08315_, _08313_);
  and (_08317_, _01967_, \oc8051_golden_model_1.PC [1]);
  nor (_08318_, _08317_, _07333_);
  and (_08319_, _08318_, _08316_);
  or (_08320_, _08319_, _08186_);
  and (_08321_, _08320_, _07876_);
  not (_08322_, \oc8051_golden_model_1.ACC [1]);
  nor (_08323_, _04835_, _08322_);
  and (_08324_, _04835_, _08322_);
  nor (_08325_, _08324_, _08323_);
  and (_08326_, _08325_, _07332_);
  or (_08327_, _08326_, _08321_);
  and (_08328_, _08327_, _07875_);
  and (_08329_, _08184_, _07336_);
  or (_08330_, _08329_, _07335_);
  or (_08331_, _08330_, _08328_);
  or (_08332_, _08323_, _07789_);
  and (_08333_, _08332_, _08331_);
  or (_08334_, _08333_, _01965_);
  and (_08335_, _01965_, \oc8051_golden_model_1.PC [1]);
  nor (_08336_, _08335_, _07885_);
  and (_08337_, _08336_, _08334_);
  and (_08338_, _08183_, _07890_);
  nor (_08339_, _08338_, _07345_);
  or (_08340_, _08339_, _08337_);
  nand (_08341_, _08324_, _07889_);
  and (_08342_, _08341_, _05408_);
  and (_08343_, _08342_, _08340_);
  nand (_08344_, _01936_, _01620_);
  nand (_08345_, _08180_, _08344_);
  or (_08346_, _08345_, _08343_);
  and (_08347_, _08346_, _08182_);
  and (_08348_, _03547_, _01981_);
  or (_08349_, _08348_, _08347_);
  nand (_08350_, _08348_, _08174_);
  and (_08351_, _08350_, _07906_);
  and (_08352_, _08351_, _08349_);
  nor (_08353_, _07779_, _07907_);
  nor (_08354_, _08353_, _07906_);
  or (_08355_, _08354_, _08352_);
  and (_08356_, _08355_, _07905_);
  nor (_08357_, _08209_, _07905_);
  or (_08358_, _08357_, _02646_);
  or (_08359_, _08358_, _08356_);
  nand (_08360_, _02646_, _02006_);
  and (_08361_, _08360_, _05802_);
  and (_08362_, _08361_, _08359_);
  and (_08363_, _01971_, _01620_);
  or (_08364_, _03287_, _08363_);
  or (_08365_, _08364_, _08362_);
  or (_08366_, _08243_, _07253_);
  and (_08367_, _08366_, _05822_);
  and (_08368_, _08367_, _08365_);
  or (_08369_, _08368_, _08175_);
  and (_08370_, _08369_, _05814_);
  and (_08371_, _08353_, _05812_);
  or (_08372_, _08371_, _07365_);
  or (_08373_, _08372_, _08370_);
  not (_08374_, _07365_);
  or (_08375_, _08209_, _08374_);
  and (_08376_, _08375_, _07544_);
  and (_08377_, _08376_, _08373_);
  or (_08378_, _08377_, _07964_);
  and (_08379_, _08378_, _08173_);
  nor (_08380_, _02646_, _02252_);
  and (_08381_, _02793_, _02646_);
  or (_08382_, _08381_, _08380_);
  and (_08383_, _08382_, _08162_);
  or (_30703_, _08383_, _08379_);
  not (_08384_, \oc8051_golden_model_1.ACC [2]);
  nor (_08385_, _04695_, _08384_);
  and (_08386_, _04695_, _08384_);
  nor (_08387_, _08386_, _08385_);
  and (_08388_, _08387_, _07332_);
  and (_08389_, _02086_, _02025_);
  and (_08390_, _04170_, _02204_);
  nand (_08391_, _05073_, _03119_);
  or (_08392_, _08391_, _08390_);
  and (_08393_, _05446_, \oc8051_golden_model_1.P3 [2]);
  nor (_08394_, _08393_, _05441_);
  and (_08395_, _08394_, _05435_);
  and (_08396_, _05444_, \oc8051_golden_model_1.P1 [2]);
  and (_08397_, _05436_, \oc8051_golden_model_1.P2 [2]);
  and (_08398_, _04552_, \oc8051_golden_model_1.P0 [2]);
  or (_08399_, _08398_, _08397_);
  nor (_08400_, _08399_, _08396_);
  and (_08401_, _08400_, _05430_);
  and (_08402_, _08401_, _08395_);
  and (_08403_, _08402_, _04650_);
  nor (_08404_, _08403_, _04554_);
  or (_08405_, _08404_, _07794_);
  nand (_08406_, _08403_, _05413_);
  or (_08407_, _08406_, _07796_);
  and (_08408_, _07801_, _03644_);
  nor (_08409_, _07801_, _03644_);
  or (_08410_, _08409_, _08408_);
  and (_08411_, _08410_, _03406_);
  nor (_08412_, _02408_, _01988_);
  and (_08413_, _01988_, \oc8051_golden_model_1.ACC [2]);
  or (_08414_, _08413_, _08412_);
  and (_08415_, _08414_, _04539_);
  or (_08416_, _08415_, _08411_);
  and (_08417_, _08416_, _07379_);
  and (_08418_, _05917_, _04695_);
  nor (_08419_, _05917_, _04695_);
  nor (_08420_, _08419_, _08418_);
  nor (_08421_, _08420_, _07379_);
  or (_08422_, _08421_, _08417_);
  or (_08423_, _08422_, _03288_);
  and (_08424_, _08423_, _08407_);
  or (_08425_, _08424_, _07558_);
  nor (_08426_, _02086_, _01995_);
  nor (_08427_, _08426_, _07290_);
  and (_08428_, _08427_, _08425_);
  and (_08430_, _07290_, _07670_);
  or (_08432_, _08430_, _07265_);
  or (_08434_, _08432_, _08428_);
  and (_08436_, _08434_, _08405_);
  or (_08438_, _08436_, _03187_);
  nand (_08440_, _05074_, _03187_);
  and (_08442_, _08440_, _07830_);
  and (_08444_, _08442_, _08438_);
  or (_08446_, _08403_, _05413_);
  and (_08447_, _08406_, _08446_);
  and (_08448_, _08447_, _07306_);
  or (_08449_, _08448_, _08444_);
  and (_08450_, _08449_, _02000_);
  nor (_08451_, _02408_, _02000_);
  or (_08452_, _08019_, _08451_);
  or (_08453_, _08452_, _08450_);
  nand (_08454_, _08019_, _05074_);
  and (_08455_, _08454_, _08023_);
  and (_08456_, _08455_, _08453_);
  nor (_08457_, _05074_, _08023_);
  or (_08458_, _08457_, _03119_);
  or (_08459_, _08458_, _08456_);
  and (_08460_, _08459_, _08392_);
  or (_08461_, _08460_, _03300_);
  nor (_08462_, _05452_, _04554_);
  and (_08463_, _04553_, \oc8051_golden_model_1.PSW [7]);
  and (_08464_, _08463_, _02439_);
  nor (_08465_, _08464_, _08462_);
  nand (_08466_, _08465_, _03300_);
  and (_08467_, _08466_, _07791_);
  and (_08468_, _08467_, _08461_);
  or (_08469_, _08468_, _08389_);
  and (_08470_, _08469_, _07970_);
  nor (_08471_, _07970_, _03644_);
  or (_08472_, _08471_, _07256_);
  or (_08473_, _08472_, _08470_);
  or (_08474_, _07856_, _04170_);
  and (_08475_, _08474_, _07259_);
  and (_08476_, _08475_, _08473_);
  nor (_08477_, _03644_, _05889_);
  and (_08478_, _05989_, \oc8051_golden_model_1.TL0 [2]);
  not (_08479_, _08478_);
  and (_08480_, _05994_, \oc8051_golden_model_1.TCON [2]);
  and (_08481_, _06002_, \oc8051_golden_model_1.SCON [2]);
  nor (_08482_, _08481_, _08480_);
  and (_08483_, _08482_, _08479_);
  and (_08484_, _05977_, \oc8051_golden_model_1.P1INREG [2]);
  and (_08485_, _06004_, \oc8051_golden_model_1.SBUF [2]);
  nor (_08486_, _08485_, _08484_);
  and (_08487_, _05982_, \oc8051_golden_model_1.P0INREG [2]);
  and (_08488_, _05999_, \oc8051_golden_model_1.TMOD [2]);
  nor (_08489_, _08488_, _08487_);
  and (_08490_, _08489_, _08486_);
  and (_08491_, _08490_, _08483_);
  and (_08492_, _06013_, \oc8051_golden_model_1.PCON [2]);
  and (_08493_, _06015_, \oc8051_golden_model_1.DPH [2]);
  nor (_08494_, _08493_, _08492_);
  and (_08495_, _08494_, _08491_);
  and (_08496_, _06063_, \oc8051_golden_model_1.TH0 [2]);
  not (_08497_, _08496_);
  and (_08498_, _06061_, \oc8051_golden_model_1.DPL [2]);
  and (_08499_, _06025_, \oc8051_golden_model_1.TH1 [2]);
  nor (_08500_, _08499_, _08498_);
  and (_08501_, _08500_, _08497_);
  and (_08502_, _06041_, \oc8051_golden_model_1.IP [2]);
  and (_08503_, _06056_, \oc8051_golden_model_1.PSW [2]);
  and (_08504_, _06047_, \oc8051_golden_model_1.ACC [2]);
  or (_08505_, _08504_, _08503_);
  or (_08506_, _08505_, _08502_);
  and (_08507_, _06033_, \oc8051_golden_model_1.P3INREG [2]);
  and (_08508_, _06050_, \oc8051_golden_model_1.B [2]);
  or (_08509_, _08508_, _08507_);
  and (_08510_, _06039_, \oc8051_golden_model_1.P2INREG [2]);
  and (_08511_, _06053_, \oc8051_golden_model_1.IE [2]);
  or (_08512_, _08511_, _08510_);
  or (_08513_, _08512_, _08509_);
  nor (_08514_, _08513_, _08506_);
  and (_08515_, _06027_, \oc8051_golden_model_1.TL1 [2]);
  and (_08516_, _06020_, \oc8051_golden_model_1.SP [2]);
  nor (_08517_, _08516_, _08515_);
  and (_08518_, _08517_, _08514_);
  and (_08519_, _08518_, _08501_);
  and (_08520_, _08519_, _08495_);
  not (_08521_, _08520_);
  nor (_08522_, _08521_, _08477_);
  nor (_08523_, _08522_, _07259_);
  or (_08524_, _08523_, _02577_);
  or (_08525_, _08524_, _08476_);
  and (_08526_, _02577_, _02439_);
  nor (_08527_, _08526_, _07326_);
  and (_08528_, _08527_, _08525_);
  and (_08529_, _07326_, _06009_);
  or (_08530_, _08529_, _01967_);
  or (_08531_, _08530_, _08528_);
  and (_08532_, _02408_, _01967_);
  nor (_08533_, _08532_, _07333_);
  and (_08534_, _08533_, _08531_);
  nor (_08535_, _04695_, _02981_);
  and (_08536_, _04695_, _02981_);
  nor (_08537_, _08536_, _08535_);
  and (_08538_, _08537_, _07333_);
  or (_08539_, _08538_, _08534_);
  and (_08540_, _08539_, _07876_);
  or (_08541_, _08540_, _08388_);
  and (_08542_, _08541_, _07875_);
  and (_08543_, _08535_, _07336_);
  or (_08544_, _08543_, _08542_);
  and (_08545_, _08544_, _07789_);
  and (_08546_, _08385_, _07335_);
  or (_08547_, _08546_, _01965_);
  or (_08548_, _08547_, _08545_);
  and (_08549_, _02408_, _01965_);
  nor (_08550_, _08549_, _07885_);
  and (_08551_, _08550_, _08548_);
  and (_08552_, _08536_, _07890_);
  nor (_08553_, _08552_, _07345_);
  or (_08554_, _08553_, _08551_);
  nand (_08555_, _08386_, _07889_);
  and (_08556_, _08555_, _05408_);
  and (_08557_, _08556_, _08554_);
  and (_08558_, _02086_, _01936_);
  or (_08559_, _07899_, _08558_);
  or (_08560_, _08559_, _08557_);
  or (_08561_, _08410_, _07898_);
  and (_08562_, _08561_, _07906_);
  and (_08563_, _08562_, _08560_);
  nor (_08564_, _07907_, _04168_);
  or (_08565_, _08564_, _07908_);
  and (_08566_, _08565_, _07353_);
  or (_08567_, _08566_, _08563_);
  and (_08568_, _08567_, _07905_);
  nor (_08569_, _08420_, _07905_);
  or (_08570_, _08569_, _02646_);
  or (_08571_, _08570_, _08568_);
  nand (_08572_, _02984_, _02646_);
  and (_08573_, _08572_, _05802_);
  and (_08574_, _08573_, _08571_);
  and (_08575_, _02086_, _01971_);
  or (_08576_, _03287_, _08575_);
  or (_08577_, _08576_, _08574_);
  not (_08578_, _05820_);
  or (_08579_, _08462_, _07253_);
  and (_08580_, _08579_, _08578_);
  and (_08581_, _08580_, _08577_);
  nor (_08582_, _07937_, _07670_);
  nor (_08583_, _08582_, _07938_);
  and (_08584_, _08583_, _07928_);
  or (_08585_, _08584_, _08581_);
  not (_08586_, _05816_);
  or (_08587_, _08583_, _08586_);
  and (_08588_, _08587_, _05814_);
  and (_08589_, _08588_, _08585_);
  or (_08590_, _07779_, _04170_);
  nor (_08591_, _07780_, _05814_);
  and (_08592_, _08591_, _08590_);
  or (_08593_, _08592_, _07365_);
  or (_08594_, _08593_, _08589_);
  nor (_08595_, _06123_, _06121_);
  nor (_08596_, _08595_, _06124_);
  or (_08597_, _08596_, _08374_);
  and (_08598_, _08597_, _07544_);
  and (_08599_, _08598_, _08594_);
  or (_08600_, _08599_, _07964_);
  or (_08601_, _07963_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_08602_, _08601_, _08163_);
  and (_08603_, _08602_, _08600_);
  and (_08604_, _02777_, _02646_);
  nor (_08605_, _02646_, _02239_);
  or (_08606_, _08605_, _08604_);
  and (_08607_, _08606_, _08162_);
  or (_30704_, _08607_, _08603_);
  or (_08608_, _07963_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_08609_, _08608_, _08163_);
  nor (_08610_, _07780_, _04120_);
  nor (_08611_, _08610_, _07781_);
  or (_08612_, _08611_, _05814_);
  nor (_08613_, _08408_, _03859_);
  or (_08614_, _08613_, _07802_);
  or (_08615_, _08614_, _07898_);
  nor (_08616_, _04649_, _02129_);
  and (_08617_, _04649_, _02129_);
  nor (_08618_, _08617_, _08616_);
  and (_08619_, _08618_, _07332_);
  nor (_08620_, _04649_, _02945_);
  and (_08621_, _04649_, _02945_);
  nor (_08622_, _08621_, _08620_);
  and (_08623_, _08622_, _07333_);
  nand (_08624_, _07255_, _03859_);
  nor (_08625_, _05646_, _04559_);
  and (_08626_, _06531_, _02439_);
  nor (_08627_, _08626_, _08625_);
  nor (_08628_, _08627_, _07792_);
  and (_08629_, _05446_, \oc8051_golden_model_1.P3 [3]);
  and (_08630_, _05444_, \oc8051_golden_model_1.P1 [3]);
  and (_08631_, _05436_, \oc8051_golden_model_1.P2 [3]);
  and (_08632_, _04552_, \oc8051_golden_model_1.P0 [3]);
  or (_08633_, _08632_, _08631_);
  or (_08634_, _08633_, _08630_);
  nor (_08635_, _08634_, _08629_);
  and (_08636_, _08635_, _05620_);
  nand (_08637_, _08636_, _05626_);
  nor (_08638_, _08637_, _05632_);
  and (_08639_, _08638_, _04548_);
  nor (_08640_, _08639_, _04559_);
  or (_08641_, _08640_, _07794_);
  nand (_08642_, _08639_, _05606_);
  or (_08643_, _08642_, _07796_);
  and (_08644_, _05917_, _04696_);
  nor (_08645_, _08418_, _04649_);
  nor (_08646_, _08645_, _08644_);
  nor (_08647_, _08646_, _07379_);
  or (_08648_, _08614_, _04539_);
  nor (_08649_, _02108_, _01988_);
  and (_08650_, _01988_, \oc8051_golden_model_1.ACC [3]);
  or (_08651_, _08650_, _08649_);
  nor (_08652_, _08651_, _03406_);
  nor (_08653_, _08652_, _07283_);
  and (_08654_, _08653_, _08648_);
  or (_08655_, _08654_, _03288_);
  or (_08656_, _08655_, _08647_);
  and (_08657_, _08656_, _08643_);
  or (_08658_, _08657_, _07558_);
  nor (_08659_, _02107_, _01995_);
  nor (_08660_, _08659_, _07290_);
  and (_08661_, _08660_, _08658_);
  and (_08662_, _07290_, _07936_);
  or (_08663_, _08662_, _07265_);
  or (_08664_, _08663_, _08661_);
  and (_08665_, _08664_, _08641_);
  or (_08666_, _08665_, _03187_);
  nand (_08667_, _05138_, _03187_);
  and (_08668_, _08667_, _07830_);
  and (_08669_, _08668_, _08666_);
  nor (_08670_, _08639_, _05606_);
  not (_08671_, _08670_);
  and (_08672_, _08642_, _08671_);
  and (_08673_, _08672_, _07306_);
  or (_08674_, _08673_, _08669_);
  and (_08675_, _08674_, _02000_);
  nor (_08676_, _02108_, _02000_);
  and (_08677_, _03118_, _01927_);
  nor (_08678_, _08677_, _08676_);
  nand (_08679_, _08678_, _07517_);
  or (_08680_, _08679_, _08675_);
  and (_08681_, _04120_, _02204_);
  nand (_08682_, _05137_, _03119_);
  or (_08683_, _08682_, _08681_);
  nand (_08684_, _05138_, _03200_);
  and (_08685_, _08684_, _07792_);
  and (_08686_, _08685_, _08683_);
  and (_08687_, _08686_, _08680_);
  or (_08688_, _08687_, _08628_);
  and (_08689_, _08688_, _07791_);
  and (_08690_, _02107_, _02025_);
  or (_08691_, _07255_, _08690_);
  or (_08692_, _08691_, _08689_);
  and (_08693_, _08692_, _08624_);
  or (_08694_, _08693_, _07256_);
  or (_08695_, _07856_, _04120_);
  and (_08696_, _08695_, _07259_);
  and (_08697_, _08696_, _08694_);
  nor (_08698_, _03859_, _05889_);
  and (_08699_, _05994_, \oc8051_golden_model_1.TCON [3]);
  not (_08700_, _08699_);
  and (_08701_, _05982_, \oc8051_golden_model_1.P0INREG [3]);
  and (_08702_, _05999_, \oc8051_golden_model_1.TMOD [3]);
  nor (_08703_, _08702_, _08701_);
  and (_08704_, _08703_, _08700_);
  and (_08705_, _05989_, \oc8051_golden_model_1.TL0 [3]);
  and (_08706_, _06002_, \oc8051_golden_model_1.SCON [3]);
  nor (_08707_, _08706_, _08705_);
  and (_08708_, _05977_, \oc8051_golden_model_1.P1INREG [3]);
  and (_08709_, _06004_, \oc8051_golden_model_1.SBUF [3]);
  nor (_08710_, _08709_, _08708_);
  and (_08711_, _08710_, _08707_);
  and (_08712_, _08711_, _08704_);
  and (_08713_, _06013_, \oc8051_golden_model_1.PCON [3]);
  and (_08714_, _06015_, \oc8051_golden_model_1.DPH [3]);
  nor (_08715_, _08714_, _08713_);
  and (_08716_, _08715_, _08712_);
  and (_08717_, _06063_, \oc8051_golden_model_1.TH0 [3]);
  not (_08718_, _08717_);
  and (_08719_, _06061_, \oc8051_golden_model_1.DPL [3]);
  and (_08720_, _06020_, \oc8051_golden_model_1.SP [3]);
  nor (_08721_, _08720_, _08719_);
  and (_08722_, _08721_, _08718_);
  and (_08723_, _06041_, \oc8051_golden_model_1.IP [3]);
  not (_08724_, _08723_);
  and (_08725_, _06053_, \oc8051_golden_model_1.IE [3]);
  and (_08726_, _06056_, \oc8051_golden_model_1.PSW [3]);
  nor (_08727_, _08726_, _08725_);
  and (_08728_, _08727_, _08724_);
  and (_08729_, _06047_, \oc8051_golden_model_1.ACC [3]);
  and (_08730_, _06050_, \oc8051_golden_model_1.B [3]);
  nor (_08731_, _08730_, _08729_);
  and (_08732_, _06039_, \oc8051_golden_model_1.P2INREG [3]);
  and (_08733_, _06033_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_08734_, _08733_, _08732_);
  and (_08735_, _08734_, _08731_);
  and (_08736_, _08735_, _08728_);
  and (_08737_, _06025_, \oc8051_golden_model_1.TH1 [3]);
  and (_08738_, _06027_, \oc8051_golden_model_1.TL1 [3]);
  nor (_08739_, _08738_, _08737_);
  and (_08740_, _08739_, _08736_);
  and (_08741_, _08740_, _08722_);
  and (_08742_, _08741_, _08716_);
  not (_08743_, _08742_);
  nor (_08744_, _08743_, _08698_);
  nor (_08745_, _08744_, _07259_);
  or (_08746_, _08745_, _02577_);
  or (_08747_, _08746_, _08697_);
  not (_08748_, _02577_);
  nor (_08749_, _08748_, _02405_);
  nor (_08750_, _08749_, _07326_);
  and (_08751_, _08750_, _08747_);
  and (_08752_, _07326_, _05986_);
  or (_08753_, _08752_, _01967_);
  or (_08754_, _08753_, _08751_);
  and (_08755_, _02108_, _01967_);
  nor (_08756_, _08755_, _07333_);
  and (_08757_, _08756_, _08754_);
  or (_08758_, _08757_, _08623_);
  and (_08759_, _08758_, _07876_);
  or (_08760_, _08759_, _08619_);
  and (_08761_, _08760_, _07875_);
  and (_08762_, _08620_, _07336_);
  or (_08763_, _08762_, _07335_);
  or (_08764_, _08763_, _08761_);
  or (_08765_, _08616_, _07789_);
  and (_08766_, _08765_, _08764_);
  or (_08767_, _08766_, _01965_);
  and (_08768_, _02108_, _01965_);
  nor (_08769_, _08768_, _07885_);
  and (_08770_, _08769_, _08767_);
  and (_08771_, _08621_, _07890_);
  nor (_08772_, _08771_, _07345_);
  or (_08773_, _08772_, _08770_);
  nand (_08774_, _08617_, _07889_);
  and (_08775_, _08774_, _05408_);
  and (_08776_, _08775_, _08773_);
  and (_08777_, _02107_, _01936_);
  or (_08778_, _07899_, _08777_);
  or (_08779_, _08778_, _08776_);
  and (_08780_, _08779_, _08615_);
  or (_08781_, _08780_, _07353_);
  nor (_08782_, _07908_, _04118_);
  or (_08783_, _07909_, _07906_);
  or (_08784_, _08783_, _08782_);
  and (_08785_, _08784_, _07905_);
  and (_08786_, _08785_, _08781_);
  nor (_08787_, _08646_, _07905_);
  or (_08788_, _08787_, _02646_);
  or (_08789_, _08788_, _08786_);
  nand (_08790_, _02948_, _02646_);
  and (_08791_, _08790_, _08789_);
  or (_08792_, _08791_, _01971_);
  and (_08793_, _02108_, _01971_);
  nor (_08794_, _08793_, _03287_);
  and (_08795_, _08794_, _08792_);
  and (_08796_, _08625_, _03287_);
  or (_08797_, _08796_, _08795_);
  and (_08798_, _08797_, _05822_);
  or (_08799_, _07938_, _07936_);
  nor (_08800_, _07939_, _05822_);
  and (_08801_, _08800_, _08799_);
  or (_08802_, _08801_, _05812_);
  or (_08803_, _08802_, _08798_);
  and (_08804_, _08803_, _08612_);
  or (_08805_, _08804_, _07365_);
  nor (_08806_, _06124_, _06120_);
  nor (_08807_, _08806_, _06125_);
  or (_08808_, _08807_, _08374_);
  and (_08809_, _08808_, _07544_);
  and (_08810_, _08809_, _08805_);
  or (_08811_, _08810_, _07964_);
  and (_08812_, _08811_, _08609_);
  and (_08813_, _05786_, _02243_);
  and (_08814_, _02784_, _02646_);
  or (_08815_, _08814_, _08813_);
  and (_08816_, _08815_, _08162_);
  or (_30705_, _08816_, _08812_);
  or (_08817_, _07963_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_08818_, _08817_, _08163_);
  nor (_08819_, _07781_, _04012_);
  nor (_08820_, _08819_, _07782_);
  or (_08821_, _08820_, _05814_);
  nor (_08822_, _07909_, _04014_);
  or (_08823_, _08822_, _07910_);
  and (_08824_, _08823_, _07353_);
  and (_08825_, _02372_, _01936_);
  not (_08826_, \oc8051_golden_model_1.ACC [4]);
  nor (_08827_, _04741_, _08826_);
  and (_08828_, _04741_, _08826_);
  nor (_08830_, _08828_, _08827_);
  and (_08831_, _08830_, _07332_);
  and (_08832_, _02372_, _02025_);
  and (_08833_, _04012_, _02204_);
  nand (_08834_, _05123_, _03119_);
  or (_08835_, _08834_, _08833_);
  nor (_08836_, _08644_, _04741_);
  and (_08837_, _08644_, _04741_);
  nor (_08838_, _08837_, _08836_);
  nor (_08839_, _08838_, _07379_);
  or (_08841_, _07798_, _04012_);
  and (_08842_, _07802_, _04325_);
  nor (_08843_, _07802_, _04325_);
  or (_08844_, _08843_, _08842_);
  and (_08845_, _08844_, _03406_);
  or (_08846_, _02372_, _01988_);
  nand (_08847_, _01988_, _08826_);
  and (_08848_, _08847_, _08846_);
  and (_08849_, _08848_, _04539_);
  or (_08850_, _08849_, _04545_);
  or (_08852_, _08850_, _08845_);
  and (_08853_, _08852_, _07379_);
  and (_08854_, _08853_, _08841_);
  or (_08855_, _08854_, _08839_);
  and (_08856_, _08855_, _07796_);
  and (_08857_, _05444_, \oc8051_golden_model_1.P1 [4]);
  not (_08858_, _08857_);
  and (_08859_, _04552_, \oc8051_golden_model_1.P0 [4]);
  nor (_08860_, _08859_, _05497_);
  and (_08861_, _08860_, _08858_);
  and (_08863_, _05436_, \oc8051_golden_model_1.P2 [4]);
  and (_08864_, _05446_, \oc8051_golden_model_1.P3 [4]);
  nor (_08865_, _08864_, _08863_);
  and (_08866_, _08865_, _08861_);
  and (_08867_, _08866_, _05490_);
  and (_08868_, _08867_, _04697_);
  nand (_08869_, _08868_, _05504_);
  and (_08870_, _08869_, _03288_);
  or (_08871_, _08870_, _07558_);
  or (_08872_, _08871_, _08856_);
  nor (_08874_, _02372_, _01995_);
  nor (_08875_, _08874_, _07290_);
  and (_08876_, _08875_, _08872_);
  and (_08877_, _07290_, _07935_);
  or (_08878_, _08877_, _07265_);
  or (_08879_, _08878_, _08876_);
  nor (_08880_, _08868_, _05503_);
  or (_08881_, _08880_, _07794_);
  and (_08882_, _08881_, _08879_);
  or (_08883_, _08882_, _03187_);
  nand (_08885_, _05124_, _03187_);
  and (_08886_, _08885_, _07830_);
  and (_08887_, _08886_, _08883_);
  nor (_08888_, _08868_, _05504_);
  not (_08889_, _08888_);
  and (_08890_, _08869_, _08889_);
  and (_08891_, _08890_, _07306_);
  or (_08892_, _08891_, _08887_);
  and (_08893_, _08892_, _02000_);
  nor (_08894_, _02373_, _02000_);
  or (_08896_, _08894_, _08019_);
  or (_08897_, _08896_, _08893_);
  nand (_08898_, _08019_, _05124_);
  and (_08899_, _08898_, _08023_);
  and (_08900_, _08899_, _08897_);
  nor (_08901_, _05124_, _08023_);
  or (_08902_, _08901_, _03119_);
  or (_08903_, _08902_, _08900_);
  and (_08904_, _08903_, _08835_);
  or (_08905_, _08904_, _03300_);
  nor (_08906_, _05503_, _05502_);
  and (_08907_, _08033_, _04123_);
  nor (_08908_, _08907_, _08906_);
  nand (_08909_, _08908_, _03300_);
  and (_08910_, _08909_, _07791_);
  and (_08911_, _08910_, _08905_);
  or (_08912_, _08911_, _08832_);
  and (_08913_, _08912_, _07970_);
  nor (_08914_, _07970_, _04325_);
  or (_08915_, _08914_, _07256_);
  or (_08916_, _08915_, _08913_);
  not (_08917_, _07475_);
  or (_08918_, _07856_, _04012_);
  and (_08919_, _08918_, _08917_);
  and (_08920_, _08919_, _08916_);
  nor (_08921_, _04325_, _05889_);
  and (_08922_, _06013_, \oc8051_golden_model_1.PCON [4]);
  and (_08923_, _06015_, \oc8051_golden_model_1.DPH [4]);
  nor (_08924_, _08923_, _08922_);
  and (_08925_, _05982_, \oc8051_golden_model_1.P0INREG [4]);
  not (_08926_, _08925_);
  and (_08927_, _05999_, \oc8051_golden_model_1.TMOD [4]);
  and (_08928_, _06004_, \oc8051_golden_model_1.SBUF [4]);
  nor (_08929_, _08928_, _08927_);
  and (_08930_, _08929_, _08926_);
  and (_08931_, _05989_, \oc8051_golden_model_1.TL0 [4]);
  and (_08932_, _05977_, \oc8051_golden_model_1.P1INREG [4]);
  nor (_08933_, _08932_, _08931_);
  and (_08934_, _05994_, \oc8051_golden_model_1.TCON [4]);
  and (_08935_, _06002_, \oc8051_golden_model_1.SCON [4]);
  nor (_08936_, _08935_, _08934_);
  and (_08937_, _08936_, _08933_);
  and (_08938_, _08937_, _08930_);
  and (_08939_, _08938_, _08924_);
  and (_08940_, _06020_, \oc8051_golden_model_1.SP [4]);
  not (_08941_, _08940_);
  and (_08942_, _06061_, \oc8051_golden_model_1.DPL [4]);
  and (_08943_, _06063_, \oc8051_golden_model_1.TH0 [4]);
  nor (_08944_, _08943_, _08942_);
  and (_08945_, _08944_, _08941_);
  and (_08946_, _06056_, \oc8051_golden_model_1.PSW [4]);
  and (_08947_, _06047_, \oc8051_golden_model_1.ACC [4]);
  nor (_08948_, _08947_, _08946_);
  and (_08949_, _06041_, \oc8051_golden_model_1.IP [4]);
  and (_08950_, _06050_, \oc8051_golden_model_1.B [4]);
  nor (_08951_, _08950_, _08949_);
  and (_08952_, _08951_, _08948_);
  and (_08953_, _06053_, \oc8051_golden_model_1.IE [4]);
  not (_08954_, _08953_);
  and (_08955_, _06039_, \oc8051_golden_model_1.P2INREG [4]);
  and (_08956_, _06033_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_08957_, _08956_, _08955_);
  and (_08958_, _08957_, _08954_);
  and (_08959_, _08958_, _08952_);
  and (_08960_, _06025_, \oc8051_golden_model_1.TH1 [4]);
  and (_08961_, _06027_, \oc8051_golden_model_1.TL1 [4]);
  nor (_08962_, _08961_, _08960_);
  and (_08963_, _08962_, _08959_);
  and (_08964_, _08963_, _08945_);
  and (_08965_, _08964_, _08939_);
  not (_08966_, _08965_);
  nor (_08967_, _08966_, _08921_);
  nor (_08968_, _08967_, _07259_);
  or (_08969_, _08968_, _02577_);
  or (_08970_, _08969_, _08920_);
  and (_08971_, _02577_, _02370_);
  nor (_08972_, _08971_, _07326_);
  and (_08973_, _08972_, _08970_);
  and (_08974_, _07326_, _05974_);
  or (_08975_, _08974_, _01967_);
  or (_08976_, _08975_, _08973_);
  and (_08977_, _02373_, _01967_);
  nor (_08978_, _08977_, _07333_);
  and (_08979_, _08978_, _08976_);
  nor (_08980_, _04741_, _02910_);
  and (_08981_, _04741_, _02910_);
  nor (_08982_, _08981_, _08980_);
  and (_08983_, _08982_, _07333_);
  or (_08984_, _08983_, _08979_);
  and (_08985_, _08984_, _07876_);
  or (_08986_, _08985_, _08831_);
  and (_08987_, _08986_, _07875_);
  and (_08988_, _08980_, _07336_);
  or (_08989_, _08988_, _08987_);
  and (_08990_, _08989_, _07789_);
  and (_08991_, _08827_, _07335_);
  or (_08992_, _08991_, _01965_);
  or (_08993_, _08992_, _08990_);
  and (_08994_, _02373_, _01965_);
  nor (_08995_, _08994_, _07885_);
  and (_08996_, _08995_, _08993_);
  and (_08997_, _08981_, _07890_);
  nor (_08998_, _08997_, _07345_);
  or (_08999_, _08998_, _08996_);
  nand (_09000_, _08828_, _07889_);
  and (_09001_, _09000_, _05408_);
  and (_09002_, _09001_, _08999_);
  or (_09003_, _09002_, _08825_);
  and (_09004_, _09003_, _08179_);
  nor (_09005_, _03547_, _03350_);
  not (_09006_, _09005_);
  and (_09007_, _08844_, _08178_);
  or (_09008_, _09007_, _09006_);
  or (_09009_, _09008_, _09004_);
  or (_09010_, _08844_, _09005_);
  and (_09011_, _09010_, _07906_);
  and (_09012_, _09011_, _09009_);
  or (_09013_, _09012_, _08824_);
  and (_09014_, _09013_, _07905_);
  nor (_09015_, _08838_, _07905_);
  or (_09016_, _09015_, _02646_);
  or (_09017_, _09016_, _09014_);
  nand (_09018_, _02913_, _02646_);
  and (_09019_, _09018_, _05802_);
  and (_09020_, _09019_, _09017_);
  and (_09021_, _02372_, _01971_);
  or (_09022_, _09021_, _03287_);
  or (_09023_, _09022_, _09020_);
  or (_09024_, _08906_, _07253_);
  and (_09025_, _09024_, _05822_);
  and (_09026_, _09025_, _09023_);
  nor (_09027_, _07939_, _07935_);
  nor (_09028_, _09027_, _07940_);
  and (_09029_, _09028_, _07928_);
  or (_09030_, _09029_, _05812_);
  or (_09031_, _09030_, _09026_);
  and (_09032_, _09031_, _08821_);
  or (_09033_, _09032_, _07365_);
  not (_09034_, _04741_);
  and (_09035_, _06125_, _09034_);
  nor (_09036_, _06125_, _09034_);
  nor (_09037_, _09036_, _09035_);
  or (_09038_, _09037_, _08374_);
  and (_09039_, _09038_, _07544_);
  and (_09040_, _09039_, _09033_);
  or (_09041_, _09040_, _07964_);
  and (_09042_, _09041_, _08818_);
  nor (_09043_, _02646_, _02235_);
  and (_09044_, _02773_, _02646_);
  or (_09045_, _09044_, _09043_);
  and (_09046_, _09045_, _08162_);
  or (_30706_, _09046_, _09042_);
  or (_09047_, _07963_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_09048_, _09047_, _08163_);
  nor (_09049_, _07940_, _07934_);
  nor (_09050_, _09049_, _07941_);
  and (_09051_, _09050_, _07928_);
  not (_09052_, \oc8051_golden_model_1.ACC [5]);
  nor (_09053_, _04787_, _09052_);
  and (_09054_, _04787_, _09052_);
  nor (_09055_, _09054_, _09053_);
  and (_09056_, _09055_, _07332_);
  nor (_09057_, _05692_, _05690_);
  and (_09058_, _08244_, _04123_);
  nor (_09059_, _09058_, _09057_);
  nor (_09060_, _09059_, _07792_);
  and (_09061_, _05446_, \oc8051_golden_model_1.P3 [5]);
  nor (_09062_, _09061_, _05678_);
  and (_09063_, _09062_, _05664_);
  and (_09064_, _05444_, \oc8051_golden_model_1.P1 [5]);
  and (_09065_, _05436_, \oc8051_golden_model_1.P2 [5]);
  and (_09066_, _04552_, \oc8051_golden_model_1.P0 [5]);
  or (_09067_, _09066_, _09065_);
  nor (_09068_, _09067_, _09064_);
  and (_09069_, _09068_, _05658_);
  and (_09070_, _09069_, _09063_);
  and (_09071_, _09070_, _04742_);
  nand (_09072_, _09071_, _05694_);
  or (_09073_, _09072_, _07796_);
  or (_09074_, _07798_, _03904_);
  nor (_09075_, _08842_, _04480_);
  or (_09076_, _09075_, _07803_);
  and (_09077_, _09076_, _03406_);
  and (_09078_, _01988_, \oc8051_golden_model_1.ACC [5]);
  nor (_09079_, _02337_, _01988_);
  or (_09080_, _09079_, _09078_);
  and (_09081_, _09080_, _04539_);
  or (_09082_, _09081_, _04545_);
  or (_09083_, _09082_, _09077_);
  and (_09084_, _09083_, _09074_);
  or (_09085_, _09084_, _07283_);
  nor (_09086_, _08837_, _04787_);
  nor (_09087_, _09086_, _05919_);
  nand (_09088_, _09087_, _07283_);
  and (_09089_, _09088_, _09085_);
  or (_09090_, _09089_, _03288_);
  and (_09091_, _09090_, _09073_);
  or (_09092_, _09091_, _07558_);
  nor (_09093_, _02336_, _01995_);
  nor (_09094_, _09093_, _07290_);
  and (_09095_, _09094_, _09092_);
  and (_09096_, _07290_, _07934_);
  or (_09097_, _09096_, _07265_);
  or (_09098_, _09097_, _09095_);
  nor (_09099_, _09071_, _05692_);
  or (_09100_, _09099_, _07794_);
  and (_09101_, _09100_, _09098_);
  or (_09102_, _09101_, _03187_);
  nand (_09103_, _05151_, _03187_);
  and (_09104_, _09103_, _07830_);
  and (_09105_, _09104_, _09102_);
  nor (_09106_, _09071_, _05694_);
  not (_09107_, _09106_);
  and (_09108_, _09072_, _09107_);
  and (_09109_, _09108_, _07306_);
  or (_09110_, _09109_, _09105_);
  and (_09111_, _09110_, _02000_);
  nor (_09112_, _02337_, _02000_);
  or (_09113_, _09112_, _03200_);
  or (_09114_, _09113_, _09111_);
  nand (_09115_, _05151_, _03200_);
  and (_09116_, _09115_, _09114_);
  or (_09117_, _09116_, _03119_);
  and (_09118_, _03904_, _02204_);
  nand (_09119_, _05150_, _03119_);
  or (_09120_, _09119_, _09118_);
  and (_09121_, _09120_, _07792_);
  and (_09122_, _09121_, _09117_);
  or (_09123_, _09122_, _09060_);
  and (_09124_, _09123_, _07791_);
  and (_09125_, _02336_, _02025_);
  or (_09126_, _09125_, _07255_);
  or (_09127_, _09126_, _09124_);
  nand (_09128_, _07255_, _04480_);
  and (_09129_, _09128_, _09127_);
  or (_09130_, _09129_, _07256_);
  or (_09131_, _07856_, _03904_);
  and (_09132_, _09131_, _07259_);
  and (_09133_, _09132_, _09130_);
  nor (_09134_, _04480_, _05889_);
  and (_09135_, _06002_, \oc8051_golden_model_1.SCON [5]);
  not (_09136_, _09135_);
  and (_09137_, _05994_, \oc8051_golden_model_1.TCON [5]);
  and (_09138_, _06004_, \oc8051_golden_model_1.SBUF [5]);
  nor (_09139_, _09138_, _09137_);
  and (_09140_, _09139_, _09136_);
  and (_09141_, _05989_, \oc8051_golden_model_1.TL0 [5]);
  and (_09142_, _05977_, \oc8051_golden_model_1.P1INREG [5]);
  nor (_09143_, _09142_, _09141_);
  and (_09144_, _05982_, \oc8051_golden_model_1.P0INREG [5]);
  and (_09145_, _05999_, \oc8051_golden_model_1.TMOD [5]);
  nor (_09146_, _09145_, _09144_);
  and (_09147_, _09146_, _09143_);
  and (_09148_, _09147_, _09140_);
  and (_09149_, _06013_, \oc8051_golden_model_1.PCON [5]);
  and (_09150_, _06015_, \oc8051_golden_model_1.DPH [5]);
  nor (_09151_, _09150_, _09149_);
  and (_09152_, _09151_, _09148_);
  and (_09153_, _06025_, \oc8051_golden_model_1.TH1 [5]);
  not (_09154_, _09153_);
  and (_09155_, _06061_, \oc8051_golden_model_1.DPL [5]);
  and (_09156_, _06020_, \oc8051_golden_model_1.SP [5]);
  nor (_09157_, _09156_, _09155_);
  and (_09158_, _09157_, _09154_);
  and (_09159_, _06039_, \oc8051_golden_model_1.P2INREG [5]);
  not (_09160_, _09159_);
  and (_09161_, _06033_, \oc8051_golden_model_1.P3INREG [5]);
  and (_09162_, _06050_, \oc8051_golden_model_1.B [5]);
  nor (_09163_, _09162_, _09161_);
  and (_09164_, _09163_, _09160_);
  and (_09165_, _06041_, \oc8051_golden_model_1.IP [5]);
  and (_09166_, _06056_, \oc8051_golden_model_1.PSW [5]);
  nor (_09167_, _09166_, _09165_);
  and (_09168_, _06053_, \oc8051_golden_model_1.IE [5]);
  and (_09169_, _06047_, \oc8051_golden_model_1.ACC [5]);
  nor (_09170_, _09169_, _09168_);
  and (_09171_, _09170_, _09167_);
  and (_09172_, _09171_, _09164_);
  and (_09173_, _06063_, \oc8051_golden_model_1.TH0 [5]);
  and (_09174_, _06027_, \oc8051_golden_model_1.TL1 [5]);
  nor (_09175_, _09174_, _09173_);
  and (_09176_, _09175_, _09172_);
  and (_09177_, _09176_, _09158_);
  and (_09178_, _09177_, _09152_);
  not (_09179_, _09178_);
  nor (_09180_, _09179_, _09134_);
  nor (_09181_, _09180_, _07259_);
  or (_09182_, _09181_, _02577_);
  or (_09183_, _09182_, _09133_);
  and (_09184_, _02577_, _02333_);
  nor (_09185_, _09184_, _07326_);
  and (_09186_, _09185_, _09183_);
  and (_09187_, _07326_, _06036_);
  or (_09188_, _09187_, _01967_);
  or (_09189_, _09188_, _09186_);
  and (_09190_, _02337_, _01967_);
  nor (_09191_, _09190_, _07333_);
  and (_09192_, _09191_, _09189_);
  nor (_09193_, _04787_, _02873_);
  and (_09194_, _04787_, _02873_);
  nor (_09195_, _09194_, _09193_);
  and (_09196_, _09195_, _07333_);
  or (_09197_, _09196_, _09192_);
  and (_09198_, _09197_, _07876_);
  or (_09199_, _09198_, _09056_);
  and (_09200_, _09199_, _07875_);
  and (_09201_, _09193_, _07336_);
  or (_09202_, _09201_, _07335_);
  or (_09203_, _09202_, _09200_);
  or (_09204_, _09053_, _07789_);
  and (_09205_, _09204_, _09203_);
  or (_09206_, _09205_, _01965_);
  and (_09207_, _02337_, _01965_);
  nor (_09208_, _09207_, _07885_);
  and (_09209_, _09208_, _09206_);
  and (_09210_, _09194_, _07890_);
  nor (_09211_, _09210_, _07345_);
  or (_09212_, _09211_, _09209_);
  nand (_09213_, _09054_, _07889_);
  and (_09214_, _09213_, _05408_);
  and (_09215_, _09214_, _09212_);
  and (_09216_, _02336_, _01936_);
  or (_09217_, _09216_, _07899_);
  or (_09218_, _09217_, _09215_);
  or (_09219_, _09076_, _07898_);
  and (_09220_, _09219_, _07906_);
  and (_09221_, _09220_, _09218_);
  nor (_09222_, _07910_, _03906_);
  or (_09223_, _09222_, _07911_);
  and (_09224_, _09223_, _07353_);
  or (_09225_, _09224_, _09221_);
  and (_09226_, _09225_, _07905_);
  nor (_09227_, _09087_, _07905_);
  or (_09228_, _09227_, _02646_);
  or (_09229_, _09228_, _09226_);
  nand (_09230_, _02877_, _02646_);
  and (_09231_, _09230_, _05802_);
  and (_09232_, _09231_, _09229_);
  and (_09233_, _02336_, _01971_);
  or (_09234_, _09233_, _03287_);
  or (_09235_, _09234_, _09232_);
  or (_09236_, _09057_, _07253_);
  and (_09237_, _09236_, _05822_);
  and (_09238_, _09237_, _09235_);
  or (_09239_, _09238_, _09051_);
  and (_09240_, _09239_, _05814_);
  or (_09241_, _07782_, _03904_);
  nor (_09242_, _07783_, _05814_);
  and (_09243_, _09242_, _09241_);
  or (_09244_, _09243_, _07365_);
  or (_09245_, _09244_, _09240_);
  and (_09246_, _09035_, _04787_);
  nor (_09247_, _09035_, _04787_);
  or (_09248_, _09247_, _09246_);
  or (_09249_, _09248_, _08374_);
  and (_09250_, _09249_, _07544_);
  and (_09251_, _09250_, _09245_);
  or (_09252_, _09251_, _07964_);
  and (_09253_, _09252_, _09048_);
  and (_09254_, _05786_, _02230_);
  and (_09255_, _02768_, _02646_);
  or (_09256_, _09255_, _09254_);
  and (_09257_, _09256_, _08162_);
  or (_30707_, _09257_, _09253_);
  nor (_09258_, _07783_, _03960_);
  nor (_09259_, _09258_, _07784_);
  or (_09260_, _09259_, _05814_);
  nor (_09261_, _07911_, _03958_);
  or (_09262_, _09261_, _07912_);
  and (_09263_, _09262_, _07353_);
  and (_09264_, _02298_, _01936_);
  not (_09265_, \oc8051_golden_model_1.ACC [6]);
  nor (_09266_, _04937_, _09265_);
  and (_09267_, _04937_, _09265_);
  nor (_09268_, _09267_, _09266_);
  and (_09269_, _09268_, _07332_);
  nor (_09270_, _05598_, _05596_);
  and (_09271_, _08463_, _04123_);
  nor (_09272_, _09271_, _09270_);
  nor (_09273_, _09272_, _07792_);
  nand (_09274_, _05087_, _03200_);
  and (_09275_, _05444_, \oc8051_golden_model_1.P1 [6]);
  not (_09276_, _09275_);
  and (_09277_, _04552_, \oc8051_golden_model_1.P0 [6]);
  nor (_09278_, _09277_, _05586_);
  and (_09279_, _09278_, _09276_);
  and (_09280_, _05436_, \oc8051_golden_model_1.P2 [6]);
  and (_09281_, _05446_, \oc8051_golden_model_1.P3 [6]);
  nor (_09282_, _09281_, _09280_);
  and (_09283_, _09282_, _09279_);
  and (_09284_, _09283_, _05572_);
  and (_09285_, _09284_, _04890_);
  nor (_09286_, _09285_, _05598_);
  or (_09287_, _09286_, _07794_);
  or (_09288_, _07798_, _03960_);
  nor (_09289_, _07803_, _04373_);
  or (_09290_, _09289_, _07804_);
  and (_09291_, _09290_, _03406_);
  or (_09292_, _02298_, _01988_);
  nand (_09293_, _01988_, _09265_);
  and (_09294_, _09293_, _09292_);
  and (_09295_, _09294_, _04539_);
  or (_09296_, _09295_, _04545_);
  or (_09297_, _09296_, _09291_);
  and (_09298_, _09297_, _07379_);
  and (_09299_, _09298_, _09288_);
  nor (_09300_, _05919_, _04937_);
  nor (_09301_, _09300_, _05921_);
  nor (_09302_, _09301_, _07379_);
  or (_09303_, _09302_, _03288_);
  or (_09304_, _09303_, _09299_);
  nand (_09305_, _09285_, _05600_);
  or (_09306_, _09305_, _07796_);
  and (_09307_, _09306_, _09304_);
  or (_09308_, _09307_, _07558_);
  nor (_09309_, _02298_, _01995_);
  nor (_09310_, _09309_, _07290_);
  and (_09311_, _09310_, _09308_);
  and (_09312_, _07290_, _07933_);
  or (_09313_, _09312_, _07265_);
  or (_09314_, _09313_, _09311_);
  and (_09315_, _09314_, _09287_);
  or (_09316_, _09315_, _03187_);
  nand (_09317_, _05087_, _03187_);
  and (_09318_, _09317_, _07830_);
  nand (_09319_, _09318_, _09316_);
  nor (_09320_, _09285_, _05600_);
  nand (_09321_, _09305_, _07306_);
  or (_09322_, _09321_, _09320_);
  nand (_09323_, _09322_, _09319_);
  and (_09324_, _09323_, _02000_);
  nor (_09325_, _02299_, _02000_);
  or (_09326_, _09325_, _03200_);
  or (_09327_, _09326_, _09324_);
  and (_09328_, _09327_, _09274_);
  or (_09329_, _09328_, _03119_);
  and (_09330_, _03960_, _02204_);
  nand (_09331_, _05086_, _03119_);
  or (_09332_, _09331_, _09330_);
  and (_09333_, _09332_, _07792_);
  and (_09334_, _09333_, _09329_);
  or (_09335_, _09334_, _09273_);
  and (_09336_, _09335_, _07791_);
  and (_09337_, _02298_, _02025_);
  or (_09338_, _09337_, _07255_);
  or (_09339_, _09338_, _09336_);
  nand (_09340_, _07255_, _04373_);
  and (_09341_, _09340_, _09339_);
  or (_09342_, _09341_, _07256_);
  or (_09343_, _07856_, _03960_);
  and (_09344_, _09343_, _08917_);
  and (_09345_, _09344_, _09342_);
  nor (_09346_, _04373_, _05889_);
  and (_09347_, _05999_, \oc8051_golden_model_1.TMOD [6]);
  and (_09348_, _06002_, \oc8051_golden_model_1.SCON [6]);
  and (_09349_, _06004_, \oc8051_golden_model_1.SBUF [6]);
  or (_09350_, _09349_, _09348_);
  or (_09351_, _09350_, _09347_);
  and (_09352_, _05982_, \oc8051_golden_model_1.P0INREG [6]);
  and (_09353_, _05977_, \oc8051_golden_model_1.P1INREG [6]);
  or (_09354_, _09353_, _09352_);
  and (_09355_, _05994_, \oc8051_golden_model_1.TCON [6]);
  and (_09356_, _05989_, \oc8051_golden_model_1.TL0 [6]);
  or (_09357_, _09356_, _09355_);
  or (_09358_, _09357_, _09354_);
  or (_09359_, _09358_, _09351_);
  and (_09360_, _06013_, \oc8051_golden_model_1.PCON [6]);
  and (_09361_, _06015_, \oc8051_golden_model_1.DPH [6]);
  or (_09362_, _09361_, _09360_);
  or (_09363_, _09362_, _09359_);
  and (_09364_, _06061_, \oc8051_golden_model_1.DPL [6]);
  and (_09365_, _06027_, \oc8051_golden_model_1.TL1 [6]);
  and (_09366_, _06020_, \oc8051_golden_model_1.SP [6]);
  or (_09367_, _09366_, _09365_);
  or (_09368_, _09367_, _09364_);
  and (_09369_, _06033_, \oc8051_golden_model_1.P3INREG [6]);
  and (_09370_, _06039_, \oc8051_golden_model_1.P2INREG [6]);
  and (_09371_, _06047_, \oc8051_golden_model_1.ACC [6]);
  or (_09372_, _09371_, _09370_);
  or (_09373_, _09372_, _09369_);
  and (_09374_, _06053_, \oc8051_golden_model_1.IE [6]);
  and (_09375_, _06056_, \oc8051_golden_model_1.PSW [6]);
  or (_09376_, _09375_, _09374_);
  and (_09377_, _06041_, \oc8051_golden_model_1.IP [6]);
  and (_09378_, _06050_, \oc8051_golden_model_1.B [6]);
  or (_09379_, _09378_, _09377_);
  or (_09380_, _09379_, _09376_);
  or (_09381_, _09380_, _09373_);
  and (_09382_, _06025_, \oc8051_golden_model_1.TH1 [6]);
  and (_09383_, _06063_, \oc8051_golden_model_1.TH0 [6]);
  or (_09384_, _09383_, _09382_);
  or (_09385_, _09384_, _09381_);
  or (_09386_, _09385_, _09368_);
  or (_09387_, _09386_, _09363_);
  or (_09388_, _09387_, _09346_);
  and (_09389_, _09388_, _07258_);
  or (_09390_, _09389_, _02577_);
  or (_09391_, _09390_, _09345_);
  and (_09392_, _02577_, _02295_);
  nor (_09393_, _09392_, _07326_);
  and (_09394_, _09393_, _09391_);
  not (_09395_, _02834_);
  and (_09396_, _07326_, _09395_);
  or (_09397_, _09396_, _01967_);
  or (_09398_, _09397_, _09394_);
  and (_09399_, _02299_, _01967_);
  nor (_09400_, _09399_, _07333_);
  and (_09401_, _09400_, _09398_);
  nor (_09402_, _04937_, _02834_);
  and (_09403_, _04937_, _02834_);
  nor (_09404_, _09403_, _09402_);
  and (_09405_, _09404_, _07333_);
  or (_09406_, _09405_, _09401_);
  and (_09407_, _09406_, _07876_);
  or (_09408_, _09407_, _09269_);
  and (_09409_, _09408_, _07875_);
  and (_09410_, _09402_, _07336_);
  or (_09411_, _09410_, _07335_);
  or (_09412_, _09411_, _09409_);
  or (_09413_, _09266_, _07789_);
  and (_09414_, _09413_, _09412_);
  or (_09415_, _09414_, _01965_);
  and (_09416_, _02299_, _01965_);
  nor (_09417_, _09416_, _07885_);
  and (_09418_, _09417_, _09415_);
  and (_09419_, _09403_, _07890_);
  nor (_09420_, _09419_, _07345_);
  or (_09421_, _09420_, _09418_);
  nand (_09422_, _09267_, _07889_);
  and (_09423_, _09422_, _05408_);
  and (_09424_, _09423_, _09421_);
  or (_09425_, _09424_, _09264_);
  and (_09426_, _09425_, _08179_);
  and (_09427_, _09290_, _08178_);
  or (_09428_, _09427_, _09006_);
  or (_09429_, _09428_, _09426_);
  or (_09430_, _09290_, _09005_);
  and (_09431_, _09430_, _07906_);
  and (_09432_, _09431_, _09429_);
  or (_09433_, _09432_, _09263_);
  and (_09434_, _09433_, _07905_);
  nor (_09435_, _09301_, _07905_);
  or (_09436_, _09435_, _02646_);
  or (_09437_, _09436_, _09434_);
  nand (_09438_, _02838_, _02646_);
  and (_09439_, _09438_, _05802_);
  and (_09440_, _09439_, _09437_);
  and (_09441_, _02298_, _01971_);
  or (_09442_, _09441_, _03287_);
  or (_09443_, _09442_, _09440_);
  or (_09444_, _09270_, _07253_);
  and (_09445_, _09444_, _05822_);
  and (_09446_, _09445_, _09443_);
  nor (_09447_, _07941_, _07933_);
  nor (_09448_, _09447_, _07942_);
  and (_09449_, _09448_, _07928_);
  or (_09450_, _09449_, _05812_);
  or (_09451_, _09450_, _09446_);
  and (_09452_, _09451_, _09260_);
  or (_09453_, _09452_, _07365_);
  and (_09454_, _06127_, _04937_);
  nor (_09455_, _06127_, _04937_);
  or (_09456_, _09455_, _09454_);
  or (_09457_, _09456_, _08374_);
  and (_09458_, _09457_, _07544_);
  and (_09459_, _09458_, _09453_);
  or (_09460_, _09459_, _07964_);
  or (_09461_, _07963_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_09462_, _09461_, _08163_);
  and (_09463_, _09462_, _09460_);
  nor (_09464_, _02646_, _02217_);
  and (_09465_, _02755_, _02646_);
  or (_09466_, _09465_, _09464_);
  and (_09467_, _09466_, _08162_);
  or (_30708_, _09467_, _09463_);
  nand (_09468_, _07963_, _07951_);
  or (_09469_, _07963_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_09470_, _09469_, _08163_);
  and (_09471_, _09470_, _09468_);
  and (_09472_, _08162_, _07957_);
  or (_30709_, _09472_, _09471_);
  and (_09473_, _07772_, _07465_);
  and (_09474_, _09473_, _07961_);
  not (_09475_, _09474_);
  or (_09476_, _09475_, _08157_);
  and (_09477_, _08161_, _03782_);
  not (_09478_, _09477_);
  or (_09479_, _09474_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_09480_, _09479_, _09478_);
  and (_09481_, _09480_, _09476_);
  and (_09482_, _09477_, _08169_);
  or (_30713_, _09482_, _09481_);
  or (_09483_, _09475_, _08377_);
  or (_09484_, _09474_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_09485_, _09484_, _09478_);
  and (_09486_, _09485_, _09483_);
  and (_09487_, _09477_, _08382_);
  or (_30714_, _09487_, _09486_);
  or (_09488_, _09475_, _08599_);
  or (_09489_, _09474_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_09490_, _09489_, _09478_);
  and (_09491_, _09490_, _09488_);
  and (_09492_, _09477_, _08606_);
  or (_30715_, _09492_, _09491_);
  or (_09493_, _09475_, _08810_);
  or (_09494_, _09474_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_09495_, _09494_, _09478_);
  and (_09496_, _09495_, _09493_);
  and (_09497_, _09477_, _08815_);
  or (_30716_, _09497_, _09496_);
  or (_09498_, _09475_, _09040_);
  or (_09499_, _09474_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_09500_, _09499_, _09478_);
  and (_09501_, _09500_, _09498_);
  and (_09502_, _09477_, _09045_);
  or (_30717_, _09502_, _09501_);
  or (_09503_, _09475_, _09251_);
  or (_09504_, _09474_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_09505_, _09504_, _09478_);
  and (_09506_, _09505_, _09503_);
  and (_09507_, _09477_, _09256_);
  or (_30718_, _09507_, _09506_);
  or (_09508_, _09475_, _09459_);
  or (_09509_, _09474_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_09510_, _09509_, _09478_);
  and (_09511_, _09510_, _09508_);
  and (_09512_, _09477_, _09466_);
  or (_30719_, _09512_, _09511_);
  or (_09513_, _09475_, _07952_);
  or (_09514_, _09474_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_09515_, _09514_, _09478_);
  and (_09516_, _09515_, _09513_);
  and (_09517_, _09477_, _07957_);
  or (_30720_, _09517_, _09516_);
  and (_09518_, _07546_, _07370_);
  and (_09519_, _09518_, _07961_);
  or (_09520_, _09519_, \oc8051_golden_model_1.IRAM[2] [0]);
  not (_09521_, _09519_);
  or (_09522_, _09521_, _08157_);
  and (_09523_, _09522_, _09520_);
  and (_09524_, _08161_, _03112_);
  or (_09525_, _09524_, _09523_);
  not (_09526_, _09524_);
  and (_09527_, _08169_, _07756_);
  or (_09528_, _09527_, _09526_);
  and (_30759_[0], _09528_, _09525_);
  or (_09529_, _09521_, _08377_);
  or (_09530_, _09519_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_09531_, _09530_, _09526_);
  and (_09532_, _09531_, _09529_);
  and (_09533_, _08382_, _07756_);
  and (_09534_, _09533_, _09524_);
  or (_30759_[1], _09534_, _09532_);
  or (_09535_, _09521_, _08599_);
  or (_09536_, _09519_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_09537_, _09536_, _09526_);
  and (_09538_, _09537_, _09535_);
  and (_09539_, _08606_, _07756_);
  and (_09540_, _09539_, _09524_);
  or (_30759_[2], _09540_, _09538_);
  or (_09541_, _09521_, _08810_);
  or (_09542_, _09519_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_09543_, _09542_, _09526_);
  and (_09544_, _09543_, _09541_);
  and (_09545_, _08815_, _07756_);
  and (_09546_, _09545_, _09524_);
  or (_30759_[3], _09546_, _09544_);
  or (_09547_, _09521_, _09040_);
  or (_09548_, _09519_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_09549_, _09548_, _09526_);
  and (_09550_, _09549_, _09547_);
  and (_09551_, _09045_, _07756_);
  and (_09552_, _09551_, _09524_);
  or (_30759_[4], _09552_, _09550_);
  or (_09553_, _09521_, _09251_);
  or (_09554_, _09519_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_09555_, _09554_, _09526_);
  and (_09556_, _09555_, _09553_);
  and (_09557_, _09256_, _07756_);
  and (_09558_, _09557_, _09524_);
  or (_30759_[5], _09558_, _09556_);
  or (_09559_, _09521_, _09459_);
  or (_09560_, _09519_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_09561_, _09560_, _09526_);
  and (_09562_, _09561_, _09559_);
  and (_09563_, _09466_, _07756_);
  and (_09564_, _09563_, _09524_);
  or (_30759_[6], _09564_, _09562_);
  or (_09565_, _09521_, _07952_);
  or (_09566_, _09519_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_09567_, _09566_, _09526_);
  and (_09568_, _09567_, _09565_);
  and (_09569_, _09524_, _07958_);
  or (_30759_[7], _09569_, _09568_);
  and (_09570_, _07961_, _07547_);
  not (_09571_, _09570_);
  and (_09572_, _09571_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_09573_, _09570_, _08157_);
  or (_09574_, _09573_, _09572_);
  and (_09575_, _08160_, _07758_);
  not (_09576_, _09575_);
  and (_09577_, _09576_, _09574_);
  and (_09578_, _09575_, _09527_);
  or (_30760_[0], _09578_, _09577_);
  or (_09579_, _09570_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_09580_, _09579_, _09576_);
  or (_09581_, _09571_, _08377_);
  and (_09582_, _09581_, _09580_);
  and (_09583_, _09575_, _09533_);
  or (_30760_[1], _09583_, _09582_);
  or (_09584_, _09570_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_09585_, _09584_, _09576_);
  or (_09586_, _09571_, _08599_);
  and (_09587_, _09586_, _09585_);
  and (_09588_, _09575_, _09539_);
  or (_30760_[2], _09588_, _09587_);
  or (_09589_, _09570_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_09590_, _09589_, _09576_);
  or (_09591_, _09571_, _08810_);
  and (_09592_, _09591_, _09590_);
  and (_09593_, _09575_, _09545_);
  or (_30760_[3], _09593_, _09592_);
  or (_09594_, _09570_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_09595_, _09594_, _09576_);
  or (_09596_, _09571_, _09040_);
  and (_09597_, _09596_, _09595_);
  and (_09598_, _09575_, _09551_);
  or (_30760_[4], _09598_, _09597_);
  or (_09599_, _09570_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_09600_, _09599_, _09576_);
  or (_09601_, _09571_, _09251_);
  and (_09602_, _09601_, _09600_);
  and (_09603_, _09575_, _09557_);
  or (_30760_[5], _09603_, _09602_);
  or (_09604_, _09570_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_09605_, _09604_, _09576_);
  or (_09606_, _09571_, _09459_);
  and (_09607_, _09606_, _09605_);
  and (_09608_, _09575_, _09563_);
  or (_30760_[6], _09608_, _09607_);
  or (_09609_, _09570_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_09610_, _09609_, _09576_);
  or (_09611_, _09571_, _07952_);
  and (_09612_, _09611_, _09610_);
  and (_09613_, _09575_, _07958_);
  or (_30760_[7], _09613_, _09612_);
  and (_09614_, _07748_, _07658_);
  and (_09615_, _09614_, _07960_);
  not (_09616_, _09615_);
  or (_09617_, _09616_, _08157_);
  not (_09618_, _07765_);
  and (_09619_, _08159_, _09618_);
  and (_09620_, _09619_, _07759_);
  not (_09621_, _09620_);
  or (_09622_, _09615_, \oc8051_golden_model_1.IRAM[4] [0]);
  and (_09623_, _09622_, _09621_);
  and (_09624_, _09623_, _09617_);
  and (_09625_, _09620_, _09527_);
  or (_30761_[0], _09625_, _09624_);
  or (_09626_, _09616_, _08377_);
  or (_09627_, _09615_, \oc8051_golden_model_1.IRAM[4] [1]);
  and (_09628_, _09627_, _09621_);
  and (_09629_, _09628_, _09626_);
  and (_09630_, _09620_, _09533_);
  or (_30761_[1], _09630_, _09629_);
  or (_09631_, _09616_, _08599_);
  or (_09632_, _09615_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_09633_, _09632_, _09621_);
  and (_09634_, _09633_, _09631_);
  and (_09635_, _09620_, _09539_);
  or (_30761_[2], _09635_, _09634_);
  or (_09636_, _09616_, _08810_);
  or (_09637_, _09615_, \oc8051_golden_model_1.IRAM[4] [3]);
  and (_09638_, _09637_, _09621_);
  and (_09639_, _09638_, _09636_);
  and (_09640_, _09620_, _09545_);
  or (_30761_[3], _09640_, _09639_);
  or (_09641_, _09616_, _09040_);
  or (_09642_, _09615_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_09643_, _09642_, _09621_);
  and (_09644_, _09643_, _09641_);
  and (_09645_, _09620_, _09551_);
  or (_30761_[4], _09645_, _09644_);
  or (_09646_, _09616_, _09251_);
  or (_09647_, _09615_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_09648_, _09647_, _09621_);
  and (_09649_, _09648_, _09646_);
  and (_09650_, _09620_, _09557_);
  or (_30761_[5], _09650_, _09649_);
  or (_09651_, _09616_, _09459_);
  or (_09652_, _09615_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_09653_, _09652_, _09621_);
  and (_09654_, _09653_, _09651_);
  and (_09655_, _09620_, _09563_);
  or (_30761_[6], _09655_, _09654_);
  or (_09656_, _09616_, _07952_);
  or (_09657_, _09615_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_09658_, _09657_, _09621_);
  and (_09659_, _09658_, _09656_);
  and (_09660_, _09620_, _07958_);
  or (_30761_[7], _09660_, _09659_);
  and (_09661_, _09614_, _09473_);
  not (_09662_, _09661_);
  or (_09663_, _09662_, _08157_);
  and (_09664_, _09619_, _03782_);
  not (_09665_, _09664_);
  or (_09666_, _09661_, \oc8051_golden_model_1.IRAM[5] [0]);
  and (_09667_, _09666_, _09665_);
  and (_09668_, _09667_, _09663_);
  and (_09669_, _09664_, _09527_);
  or (_30762_[0], _09669_, _09668_);
  or (_09670_, _09662_, _08377_);
  or (_09671_, _09661_, \oc8051_golden_model_1.IRAM[5] [1]);
  and (_09672_, _09671_, _09665_);
  and (_09673_, _09672_, _09670_);
  and (_09674_, _09664_, _09533_);
  or (_30762_[1], _09674_, _09673_);
  or (_09675_, _09662_, _08599_);
  or (_09676_, _09661_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_09677_, _09676_, _09665_);
  and (_09678_, _09677_, _09675_);
  and (_09679_, _09664_, _09539_);
  or (_30762_[2], _09679_, _09678_);
  or (_09680_, _09662_, _08810_);
  or (_09681_, _09661_, \oc8051_golden_model_1.IRAM[5] [3]);
  and (_09682_, _09681_, _09665_);
  and (_09683_, _09682_, _09680_);
  and (_09684_, _09664_, _09545_);
  or (_30762_[3], _09684_, _09683_);
  or (_09685_, _09662_, _09040_);
  or (_09686_, _09661_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_09687_, _09686_, _09665_);
  and (_09688_, _09687_, _09685_);
  and (_09689_, _09664_, _09551_);
  or (_30762_[4], _09689_, _09688_);
  or (_09690_, _09662_, _09251_);
  or (_09691_, _09661_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_09692_, _09691_, _09665_);
  and (_09693_, _09692_, _09690_);
  and (_09694_, _09664_, _09557_);
  or (_30762_[5], _09694_, _09693_);
  or (_09695_, _09662_, _09459_);
  or (_09696_, _09661_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_09697_, _09696_, _09665_);
  and (_09698_, _09697_, _09695_);
  and (_09699_, _09664_, _09563_);
  or (_30762_[6], _09699_, _09698_);
  or (_09700_, _09662_, _07952_);
  or (_09701_, _09661_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_09702_, _09701_, _09665_);
  and (_09703_, _09702_, _09700_);
  and (_09704_, _09664_, _07958_);
  or (_30762_[7], _09704_, _09703_);
  and (_09705_, _09614_, _09518_);
  not (_09706_, _09705_);
  or (_09707_, _09706_, _08157_);
  and (_09708_, _09619_, _03112_);
  not (_09709_, _09708_);
  or (_09710_, _09705_, \oc8051_golden_model_1.IRAM[6] [0]);
  and (_09711_, _09710_, _09709_);
  and (_09712_, _09711_, _09707_);
  and (_09713_, _09708_, _09527_);
  or (_30721_, _09713_, _09712_);
  or (_09714_, _09706_, _08377_);
  or (_09715_, _09705_, \oc8051_golden_model_1.IRAM[6] [1]);
  and (_09716_, _09715_, _09709_);
  and (_09717_, _09716_, _09714_);
  and (_09718_, _09708_, _09533_);
  or (_30722_, _09718_, _09717_);
  or (_09719_, _09706_, _08599_);
  or (_09720_, _09705_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_09721_, _09720_, _09709_);
  and (_09722_, _09721_, _09719_);
  and (_09723_, _09708_, _09539_);
  or (_30723_, _09723_, _09722_);
  or (_09724_, _09706_, _08810_);
  or (_09725_, _09705_, \oc8051_golden_model_1.IRAM[6] [3]);
  and (_09726_, _09725_, _09709_);
  and (_09727_, _09726_, _09724_);
  and (_09728_, _09708_, _09545_);
  or (_30724_, _09728_, _09727_);
  or (_09729_, _09706_, _09040_);
  or (_09730_, _09705_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_09731_, _09730_, _09709_);
  and (_09732_, _09731_, _09729_);
  and (_09733_, _09708_, _09551_);
  or (_30725_, _09733_, _09732_);
  or (_09734_, _09706_, _09251_);
  or (_09735_, _09705_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_09736_, _09735_, _09709_);
  and (_09737_, _09736_, _09734_);
  and (_09738_, _09708_, _09557_);
  or (_30726_, _09738_, _09737_);
  or (_09739_, _09706_, _09459_);
  or (_09740_, _09705_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_09741_, _09740_, _09709_);
  and (_09742_, _09741_, _09739_);
  and (_09743_, _09708_, _09563_);
  or (_30727_, _09743_, _09742_);
  or (_09744_, _09706_, _07952_);
  or (_09745_, _09705_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_09746_, _09745_, _09709_);
  and (_09747_, _09746_, _09744_);
  and (_09748_, _09708_, _07958_);
  or (_30728_, _09748_, _09747_);
  and (_09749_, _09614_, _07773_);
  not (_09750_, _09749_);
  or (_09751_, _09750_, _08157_);
  and (_09752_, _09619_, _07758_);
  not (_09753_, _09752_);
  or (_09754_, _09749_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_09755_, _09754_, _09753_);
  and (_09756_, _09755_, _09751_);
  and (_09757_, _09752_, _09527_);
  or (_30729_, _09757_, _09756_);
  or (_09758_, _09749_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_09759_, _09758_, _09753_);
  or (_09760_, _09750_, _08377_);
  and (_09761_, _09760_, _09759_);
  and (_09762_, _09752_, _09533_);
  or (_30730_, _09762_, _09761_);
  or (_09763_, _09749_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_09764_, _09763_, _09753_);
  or (_09765_, _09750_, _08599_);
  and (_09766_, _09765_, _09764_);
  and (_09767_, _09752_, _09539_);
  or (_30731_, _09767_, _09766_);
  or (_09768_, _09749_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_09769_, _09768_, _09753_);
  or (_09770_, _09750_, _08810_);
  and (_09771_, _09770_, _09769_);
  and (_09772_, _09752_, _09545_);
  or (_30732_, _09772_, _09771_);
  or (_09773_, _09750_, _09040_);
  or (_09774_, _09749_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_09775_, _09774_, _09753_);
  and (_09776_, _09775_, _09773_);
  and (_09777_, _09752_, _09551_);
  or (_30733_, _09777_, _09776_);
  or (_09778_, _09749_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_09779_, _09778_, _09753_);
  or (_09780_, _09750_, _09251_);
  and (_09781_, _09780_, _09779_);
  and (_09782_, _09752_, _09557_);
  or (_30734_, _09782_, _09781_);
  or (_09783_, _09749_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_09784_, _09783_, _09753_);
  or (_09785_, _09750_, _09459_);
  and (_09786_, _09785_, _09784_);
  and (_09787_, _09752_, _09563_);
  or (_30735_, _09787_, _09786_);
  or (_09788_, _09750_, _07952_);
  or (_09789_, _09749_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_09790_, _09789_, _09753_);
  and (_09791_, _09790_, _09788_);
  and (_09792_, _09752_, _07958_);
  or (_30736_, _09792_, _09791_);
  and (_09793_, _07775_, _07747_);
  and (_09794_, _09793_, _07960_);
  nor (_09795_, _09794_, _03683_);
  and (_09796_, _09794_, _08157_);
  or (_09797_, _09796_, _09795_);
  nand (_09798_, _07766_, _07760_);
  and (_09799_, _09798_, _09797_);
  not (_09800_, _07762_);
  and (_09801_, _07766_, _09800_);
  and (_09802_, _09801_, _07759_);
  and (_09803_, _09802_, _09527_);
  or (_30737_, _09803_, _09799_);
  not (_09804_, _09794_);
  or (_09805_, _09804_, _08377_);
  or (_09806_, _09794_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_09807_, _09806_, _09798_);
  and (_09808_, _09807_, _09805_);
  and (_09809_, _09802_, _09533_);
  or (_30738_, _09809_, _09808_);
  or (_09810_, _09804_, _08599_);
  or (_09811_, _09794_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_09812_, _09811_, _09798_);
  and (_09813_, _09812_, _09810_);
  and (_09814_, _09802_, _09539_);
  or (_30739_, _09814_, _09813_);
  or (_09815_, _09804_, _08810_);
  or (_09816_, _09794_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_09817_, _09816_, _09798_);
  and (_09818_, _09817_, _09815_);
  and (_09819_, _09802_, _09545_);
  or (_30740_, _09819_, _09818_);
  or (_09820_, _09804_, _09040_);
  or (_09821_, _09794_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_09822_, _09821_, _09798_);
  and (_09823_, _09822_, _09820_);
  and (_09824_, _09802_, _09551_);
  or (_30741_, _09824_, _09823_);
  or (_09825_, _09804_, _09251_);
  or (_09826_, _09794_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_09827_, _09826_, _09798_);
  and (_09828_, _09827_, _09825_);
  and (_09829_, _09802_, _09557_);
  or (_30742_, _09829_, _09828_);
  or (_09830_, _09804_, _09459_);
  or (_09831_, _09794_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_09832_, _09831_, _09798_);
  and (_09833_, _09832_, _09830_);
  and (_09834_, _09802_, _09563_);
  or (_30743_, _09834_, _09833_);
  or (_09835_, _09804_, _07952_);
  or (_09836_, _09794_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_09837_, _09836_, _09798_);
  and (_09838_, _09837_, _09835_);
  and (_09839_, _09802_, _07958_);
  or (_30744_, _09839_, _09838_);
  and (_09840_, _09793_, _09473_);
  nor (_09841_, _09840_, _03687_);
  and (_09842_, _09840_, _08157_);
  or (_09843_, _09842_, _09841_);
  nand (_09844_, _07766_, _07552_);
  and (_09845_, _09844_, _09843_);
  and (_09846_, _09801_, _03782_);
  and (_09847_, _09846_, _09527_);
  or (_30745_, _09847_, _09845_);
  not (_09848_, _09840_);
  or (_09849_, _09848_, _08377_);
  or (_09850_, _09840_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_09851_, _09850_, _09844_);
  and (_09852_, _09851_, _09849_);
  and (_09853_, _09846_, _09533_);
  or (_30746_, _09853_, _09852_);
  or (_09854_, _09848_, _08599_);
  or (_09855_, _09840_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_09856_, _09855_, _09844_);
  and (_09857_, _09856_, _09854_);
  and (_09858_, _09846_, _09539_);
  or (_30747_, _09858_, _09857_);
  or (_09859_, _09848_, _08810_);
  or (_09860_, _09840_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_09861_, _09860_, _09844_);
  and (_09862_, _09861_, _09859_);
  and (_09863_, _09846_, _09545_);
  or (_30748_, _09863_, _09862_);
  or (_09864_, _09848_, _09040_);
  or (_09865_, _09840_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_09866_, _09865_, _09844_);
  and (_09867_, _09866_, _09864_);
  and (_09868_, _09846_, _09551_);
  or (_30749_, _09868_, _09867_);
  or (_09869_, _09848_, _09251_);
  or (_09870_, _09840_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_09871_, _09870_, _09844_);
  and (_09872_, _09871_, _09869_);
  and (_09873_, _09846_, _09557_);
  or (_30750_, _09873_, _09872_);
  or (_09874_, _09848_, _09459_);
  or (_09875_, _09840_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_09876_, _09875_, _09844_);
  and (_09877_, _09876_, _09874_);
  and (_09878_, _09846_, _09563_);
  or (_30751_, _09878_, _09877_);
  or (_09879_, _09848_, _07952_);
  or (_09880_, _09840_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_09881_, _09880_, _09844_);
  and (_09882_, _09881_, _09879_);
  and (_09883_, _09846_, _07958_);
  or (_30752_, _09883_, _09882_);
  and (_09884_, _09793_, _09518_);
  not (_09885_, _09884_);
  or (_09886_, _09885_, _08157_);
  and (_09887_, _09801_, _03112_);
  not (_09888_, _09887_);
  or (_09889_, _09884_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_09890_, _09889_, _09888_);
  and (_09891_, _09890_, _09886_);
  and (_09892_, _09887_, _09527_);
  or (_30710_, _09892_, _09891_);
  or (_09893_, _09885_, _08377_);
  or (_09894_, _09884_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_09895_, _09894_, _09888_);
  and (_09896_, _09895_, _09893_);
  and (_09897_, _09887_, _09533_);
  or (_30711_, _09897_, _09896_);
  or (_09898_, _09885_, _08599_);
  or (_09899_, _09884_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_09900_, _09899_, _09888_);
  and (_09901_, _09900_, _09898_);
  and (_09902_, _09887_, _09539_);
  or (_30712_, _09902_, _09901_);
  or (_09903_, _09885_, _08810_);
  or (_09904_, _09884_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_09905_, _09904_, _09888_);
  and (_09906_, _09905_, _09903_);
  and (_09907_, _09887_, _09545_);
  or (_30753_[3], _09907_, _09906_);
  or (_09908_, _09885_, _09040_);
  or (_09909_, _09884_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_09910_, _09909_, _09888_);
  and (_09911_, _09910_, _09908_);
  and (_09912_, _09887_, _09551_);
  or (_30753_[4], _09912_, _09911_);
  or (_09913_, _09885_, _09251_);
  or (_09914_, _09884_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_09915_, _09914_, _09888_);
  and (_09916_, _09915_, _09913_);
  and (_09917_, _09887_, _09557_);
  or (_30753_[5], _09917_, _09916_);
  or (_09918_, _09885_, _09459_);
  or (_09919_, _09884_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_09920_, _09919_, _09888_);
  and (_09921_, _09920_, _09918_);
  and (_09922_, _09887_, _09563_);
  or (_30753_[6], _09922_, _09921_);
  or (_09923_, _09885_, _07952_);
  or (_09924_, _09884_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_09925_, _09924_, _09888_);
  and (_09926_, _09925_, _09923_);
  and (_09927_, _09887_, _07958_);
  or (_30753_[7], _09927_, _09926_);
  nand (_09928_, _09793_, _07773_);
  nor (_09929_, _09928_, _08157_);
  and (_09930_, _09801_, _07758_);
  and (_09931_, _09928_, _03694_);
  or (_09932_, _09931_, _09930_);
  nor (_09933_, _09932_, _09929_);
  and (_09934_, _09930_, _09527_);
  or (_30754_[0], _09934_, _09933_);
  not (_09935_, _09930_);
  and (_09936_, _09793_, _07547_);
  or (_09937_, _09936_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_09938_, _09937_, _09935_);
  not (_09939_, _09936_);
  or (_09940_, _09939_, _08377_);
  and (_09941_, _09940_, _09938_);
  and (_09942_, _09930_, _09533_);
  or (_30754_[1], _09942_, _09941_);
  or (_09943_, _09936_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_09944_, _09943_, _09935_);
  or (_09945_, _09939_, _08599_);
  and (_09946_, _09945_, _09944_);
  and (_09947_, _09930_, _09539_);
  or (_30754_[2], _09947_, _09946_);
  or (_09948_, _09936_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_09949_, _09948_, _09935_);
  or (_09950_, _09939_, _08810_);
  and (_09951_, _09950_, _09949_);
  and (_09952_, _09930_, _09545_);
  or (_30754_[3], _09952_, _09951_);
  or (_09953_, _09936_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_09954_, _09953_, _09935_);
  or (_09955_, _09939_, _09040_);
  and (_09956_, _09955_, _09954_);
  and (_09957_, _09930_, _09551_);
  or (_30754_[4], _09957_, _09956_);
  or (_09958_, _09936_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_09959_, _09958_, _09935_);
  or (_09960_, _09939_, _09251_);
  and (_09961_, _09960_, _09959_);
  and (_09962_, _09930_, _09557_);
  or (_30754_[5], _09962_, _09961_);
  or (_09963_, _09936_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_09964_, _09963_, _09935_);
  or (_09965_, _09939_, _09459_);
  and (_09966_, _09965_, _09964_);
  and (_09967_, _09930_, _09563_);
  or (_30754_[6], _09967_, _09966_);
  or (_09968_, _09936_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_09969_, _09968_, _09935_);
  or (_09970_, _09939_, _07952_);
  and (_09971_, _09970_, _09969_);
  and (_09972_, _09930_, _07958_);
  or (_30754_[7], _09972_, _09971_);
  and (_09973_, _07960_, _07750_);
  nor (_09974_, _09973_, _03706_);
  and (_09975_, _09973_, _08157_);
  or (_09976_, _09975_, _09974_);
  and (_09977_, _07767_, _07759_);
  not (_09978_, _09977_);
  and (_09979_, _09978_, _09976_);
  and (_09980_, _09977_, _09527_);
  or (_30755_[0], _09980_, _09979_);
  or (_09981_, _09973_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_09982_, _09981_, _09978_);
  nand (_09983_, _07960_, _07776_);
  or (_09984_, _09983_, _08377_);
  and (_09985_, _09984_, _09982_);
  and (_09986_, _09977_, _09533_);
  or (_30755_[1], _09986_, _09985_);
  or (_09987_, _09973_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_09988_, _09987_, _09978_);
  or (_09989_, _09983_, _08599_);
  and (_09990_, _09989_, _09988_);
  and (_09991_, _09977_, _09539_);
  or (_30755_[2], _09991_, _09990_);
  or (_09992_, _09983_, _08810_);
  or (_09993_, _09973_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_09994_, _09993_, _09978_);
  and (_09995_, _09994_, _09992_);
  and (_09996_, _09977_, _09545_);
  or (_30755_[3], _09996_, _09995_);
  or (_09997_, _09973_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_09998_, _09997_, _09978_);
  or (_09999_, _09983_, _09040_);
  and (_10000_, _09999_, _09998_);
  and (_10001_, _09977_, _09551_);
  or (_30755_[4], _10001_, _10000_);
  or (_10002_, _09973_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_10003_, _10002_, _09978_);
  or (_10004_, _09983_, _09251_);
  and (_10005_, _10004_, _10003_);
  and (_10006_, _09977_, _09557_);
  or (_30755_[5], _10006_, _10005_);
  or (_10007_, _09973_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_10008_, _10007_, _09978_);
  or (_10009_, _09983_, _09459_);
  and (_10010_, _10009_, _10008_);
  and (_10011_, _09977_, _09563_);
  or (_30755_[6], _10011_, _10010_);
  or (_10012_, _09973_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_10013_, _10012_, _09978_);
  or (_10014_, _09983_, _07952_);
  and (_10015_, _10014_, _10013_);
  and (_10016_, _09977_, _07958_);
  or (_30755_[7], _10016_, _10015_);
  nand (_10017_, _09473_, _07776_);
  or (_10018_, _10017_, _08157_);
  and (_10019_, _07767_, _03782_);
  not (_10020_, _10019_);
  nand (_10021_, _10017_, _03708_);
  and (_10022_, _10021_, _10020_);
  and (_10023_, _10022_, _10018_);
  and (_10024_, _10019_, _09527_);
  or (_30756_[0], _10024_, _10023_);
  and (_10025_, _09473_, _07750_);
  or (_10026_, _10025_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_10027_, _10026_, _10020_);
  or (_10028_, _10017_, _08377_);
  and (_10029_, _10028_, _10027_);
  and (_10030_, _10019_, _09533_);
  or (_30756_[1], _10030_, _10029_);
  or (_10031_, _10025_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_10032_, _10031_, _10020_);
  or (_10033_, _10017_, _08599_);
  and (_10034_, _10033_, _10032_);
  and (_10035_, _10019_, _09539_);
  or (_30756_[2], _10035_, _10034_);
  or (_10036_, _10025_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_10037_, _10036_, _10020_);
  or (_10038_, _10017_, _08810_);
  and (_10039_, _10038_, _10037_);
  and (_10040_, _10019_, _09545_);
  or (_30756_[3], _10040_, _10039_);
  or (_10041_, _10025_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_10042_, _10041_, _10020_);
  or (_10043_, _10017_, _09040_);
  and (_10044_, _10043_, _10042_);
  and (_10045_, _10019_, _09551_);
  or (_30756_[4], _10045_, _10044_);
  or (_10046_, _10025_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_10047_, _10046_, _10020_);
  or (_10048_, _10017_, _09251_);
  and (_10049_, _10048_, _10047_);
  and (_10050_, _10019_, _09557_);
  or (_30756_[5], _10050_, _10049_);
  or (_10051_, _10025_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_10052_, _10051_, _10020_);
  or (_10053_, _10017_, _09459_);
  and (_10054_, _10053_, _10052_);
  and (_10055_, _10019_, _09563_);
  or (_30756_[6], _10055_, _10054_);
  or (_10056_, _10025_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_10057_, _10056_, _10020_);
  or (_10058_, _10017_, _07952_);
  and (_10059_, _10058_, _10057_);
  and (_10060_, _10019_, _07958_);
  or (_30756_[7], _10060_, _10059_);
  and (_10061_, _09518_, _07776_);
  not (_10062_, _10061_);
  or (_10063_, _10062_, _08157_);
  and (_10064_, _07767_, _03112_);
  not (_10065_, _10064_);
  or (_10066_, _10061_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_10067_, _10066_, _10065_);
  and (_10068_, _10067_, _10063_);
  and (_10069_, _10064_, _09527_);
  or (_30757_[0], _10069_, _10068_);
  and (_10070_, _09518_, _07750_);
  or (_10071_, _10070_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_10072_, _10071_, _10065_);
  or (_10073_, _10062_, _08377_);
  and (_10074_, _10073_, _10072_);
  and (_10075_, _10064_, _09533_);
  or (_30757_[1], _10075_, _10074_);
  or (_10076_, _10070_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_10077_, _10076_, _10065_);
  or (_10078_, _10062_, _08599_);
  and (_10079_, _10078_, _10077_);
  and (_10080_, _10064_, _09539_);
  or (_30757_[2], _10080_, _10079_);
  or (_10081_, _10070_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_10082_, _10081_, _10065_);
  or (_10083_, _10062_, _08810_);
  and (_10084_, _10083_, _10082_);
  and (_10085_, _10064_, _09545_);
  or (_30757_[3], _10085_, _10084_);
  or (_10086_, _10070_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_10087_, _10086_, _10065_);
  or (_10088_, _10062_, _09040_);
  and (_10089_, _10088_, _10087_);
  and (_10090_, _10064_, _09551_);
  or (_30757_[4], _10090_, _10089_);
  or (_10091_, _10070_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_10092_, _10091_, _10065_);
  or (_10093_, _10062_, _09251_);
  and (_10094_, _10093_, _10092_);
  and (_10095_, _10064_, _09557_);
  or (_30757_[5], _10095_, _10094_);
  or (_10096_, _10070_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_10097_, _10096_, _10065_);
  or (_10098_, _10062_, _09459_);
  and (_10099_, _10098_, _10097_);
  and (_10100_, _10064_, _09563_);
  or (_30757_[6], _10100_, _10099_);
  nor (_10101_, _10061_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_10102_, _10062_, _07952_);
  or (_10103_, _10102_, _10101_);
  nand (_10104_, _10103_, _10065_);
  or (_10105_, _10065_, _07958_);
  and (_30757_[7], _10105_, _10104_);
  or (_10106_, _08157_, _07777_);
  nand (_10107_, _07777_, _03701_);
  and (_10108_, _10107_, _07769_);
  and (_10109_, _10108_, _10106_);
  and (_10110_, _09527_, _07768_);
  or (_30758_[0], _10110_, _10109_);
  or (_10111_, _07751_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_10112_, _10111_, _07769_);
  or (_10113_, _08377_, _07777_);
  and (_10114_, _10113_, _10112_);
  and (_10115_, _09533_, _07768_);
  or (_30758_[1], _10115_, _10114_);
  or (_10116_, _07751_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_10117_, _10116_, _07769_);
  or (_10118_, _08599_, _07777_);
  and (_10119_, _10118_, _10117_);
  and (_10120_, _09539_, _07768_);
  or (_30758_[2], _10120_, _10119_);
  or (_10121_, _07751_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_10122_, _10121_, _07769_);
  or (_10123_, _08810_, _07777_);
  and (_10124_, _10123_, _10122_);
  and (_10125_, _09545_, _07768_);
  or (_30758_[3], _10125_, _10124_);
  or (_10126_, _07751_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_10127_, _10126_, _07769_);
  or (_10128_, _09040_, _07777_);
  and (_10129_, _10128_, _10127_);
  and (_10130_, _09551_, _07768_);
  or (_30758_[4], _10130_, _10129_);
  or (_10131_, _07751_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_10132_, _10131_, _07769_);
  or (_10133_, _09251_, _07777_);
  and (_10134_, _10133_, _10132_);
  and (_10135_, _09557_, _07768_);
  or (_30758_[5], _10135_, _10134_);
  or (_10136_, _07751_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_10137_, _10136_, _07769_);
  or (_10138_, _09459_, _07777_);
  and (_10139_, _10138_, _10137_);
  and (_10140_, _09563_, _07768_);
  or (_30758_[6], _10140_, _10139_);
  not (_10141_, \oc8051_golden_model_1.B [0]);
  or (_10142_, _10141_, rst);
  nor (_28763_, _10142_, _27788_);
  nand (_10143_, \oc8051_golden_model_1.B [1], _27053_);
  nor (_28764_, _10143_, _27788_);
  not (_10144_, \oc8051_golden_model_1.B [2]);
  or (_10145_, _10144_, rst);
  nor (_28767_, _10145_, _27788_);
  nand (_10146_, \oc8051_golden_model_1.B [3], _27053_);
  nor (_28768_, _10146_, _27788_);
  not (_10147_, \oc8051_golden_model_1.B [4]);
  or (_10148_, _10147_, rst);
  nor (_28769_, _10148_, _27788_);
  nand (_10149_, \oc8051_golden_model_1.B [5], _27053_);
  nor (_28770_, _10149_, _27788_);
  not (_10150_, \oc8051_golden_model_1.B [6]);
  or (_10151_, _10150_, rst);
  nor (_28771_, _10151_, _27788_);
  or (_10152_, _02059_, rst);
  nor (_28773_, _10152_, _27788_);
  or (_10153_, _08322_, rst);
  nor (_28776_, _10153_, _27788_);
  or (_10154_, _08384_, rst);
  nor (_28777_, _10154_, _27788_);
  or (_10155_, _02129_, rst);
  nor (_28778_, _10155_, _27788_);
  or (_10156_, _08826_, rst);
  nor (_28779_, _10156_, _27788_);
  or (_10157_, _09052_, rst);
  nor (_28780_, _10157_, _27788_);
  or (_10158_, _09265_, rst);
  nor (_28781_, _10158_, _27788_);
  not (_10159_, \oc8051_golden_model_1.DPL [0]);
  or (_10160_, _10159_, rst);
  nor (_28783_, _10160_, _27788_);
  nand (_10161_, \oc8051_golden_model_1.DPL [1], _27053_);
  nor (_28784_, _10161_, _27788_);
  not (_10162_, \oc8051_golden_model_1.DPL [2]);
  or (_10163_, _10162_, rst);
  nor (_28785_, _10163_, _27788_);
  nand (_10164_, \oc8051_golden_model_1.DPL [3], _27053_);
  nor (_28786_, _10164_, _27788_);
  not (_10165_, \oc8051_golden_model_1.DPL [4]);
  or (_10166_, _10165_, rst);
  nor (_28787_, _10166_, _27788_);
  nand (_10167_, \oc8051_golden_model_1.DPL [5], _27053_);
  nor (_28788_, _10167_, _27788_);
  not (_10168_, \oc8051_golden_model_1.DPL [6]);
  or (_10169_, _10168_, rst);
  nor (_28789_, _10169_, _27788_);
  or (_10170_, _05254_, rst);
  nor (_28794_, _10170_, _27788_);
  nand (_10171_, \oc8051_golden_model_1.DPH [1], _27053_);
  nor (_28795_, _10171_, _27788_);
  not (_10172_, \oc8051_golden_model_1.DPH [2]);
  or (_10173_, _10172_, rst);
  nor (_28796_, _10173_, _27788_);
  nand (_10174_, \oc8051_golden_model_1.DPH [3], _27053_);
  nor (_28797_, _10174_, _27788_);
  not (_10175_, \oc8051_golden_model_1.DPH [4]);
  or (_10176_, _10175_, rst);
  nor (_28798_, _10176_, _27788_);
  nand (_10177_, \oc8051_golden_model_1.DPH [5], _27053_);
  nor (_28799_, _10177_, _27788_);
  not (_10178_, \oc8051_golden_model_1.DPH [6]);
  or (_10179_, _10178_, rst);
  nor (_28800_, _10179_, _27788_);
  not (_10180_, \oc8051_golden_model_1.IE [0]);
  nor (_10181_, _04629_, _10180_);
  nor (_10182_, _04888_, _07143_);
  nor (_10183_, _10182_, _10181_);
  nor (_10184_, _10183_, _03513_);
  and (_10185_, _04629_, _04268_);
  nor (_10186_, _10181_, _05963_);
  not (_10187_, _10186_);
  nor (_10188_, _10187_, _10185_);
  nor (_10189_, _05433_, _10180_);
  and (_10190_, _07997_, _05433_);
  nor (_10191_, _10190_, _10189_);
  nor (_10192_, _10191_, _03390_);
  and (_10193_, _10183_, _02661_);
  and (_10194_, _04629_, \oc8051_golden_model_1.ACC [0]);
  nor (_10195_, _10194_, _10181_);
  nor (_10196_, _10195_, _05903_);
  nor (_10197_, _04505_, _10180_);
  or (_10198_, _10197_, _02661_);
  nor (_10199_, _10198_, _10196_);
  or (_10200_, _10199_, _06504_);
  nor (_10201_, _10200_, _10193_);
  and (_10202_, _04629_, _03716_);
  nor (_10203_, _10202_, _10181_);
  nor (_10204_, _10203_, _03365_);
  or (_10205_, _10204_, _03168_);
  or (_10206_, _10205_, _10201_);
  nor (_10207_, _10206_, _10192_);
  and (_10208_, _10195_, _03168_);
  nor (_10209_, _10208_, _03176_);
  not (_10210_, _10209_);
  nor (_10211_, _10210_, _10207_);
  and (_10212_, _10181_, _03176_);
  or (_10213_, _10212_, _10211_);
  and (_10214_, _10213_, _05168_);
  nor (_10215_, _10183_, _05168_);
  or (_10216_, _10215_, _10214_);
  nor (_10217_, _10216_, _03140_);
  nor (_10218_, _08035_, _07180_);
  or (_10219_, _10189_, _03141_);
  nor (_10220_, _10219_, _10218_);
  or (_10221_, _10220_, _05949_);
  or (_10222_, _10221_, _10217_);
  or (_10223_, _10203_, _06673_);
  and (_10224_, _10223_, _05963_);
  and (_10225_, _10224_, _10222_);
  nor (_10226_, _10225_, _10188_);
  nor (_10227_, _10226_, _02024_);
  nor (_10228_, _08093_, _07143_);
  or (_10229_, _10181_, _03139_);
  nor (_10230_, _10229_, _10228_);
  or (_10231_, _10230_, _02575_);
  nor (_10232_, _10231_, _10227_);
  and (_10233_, _04629_, _05996_);
  nor (_10234_, _10233_, _10181_);
  nand (_10235_, _10234_, _05305_);
  and (_10236_, _10235_, _06549_);
  nor (_10237_, _10236_, _10232_);
  and (_10238_, _07968_, _04629_);
  nor (_10239_, _10238_, _10181_);
  and (_10240_, _10239_, _02656_);
  nor (_10241_, _10240_, _10237_);
  and (_10242_, _10241_, _03252_);
  and (_10243_, _08110_, _04629_);
  nor (_10244_, _10243_, _10181_);
  nor (_10245_, _10244_, _03252_);
  or (_10246_, _10245_, _10242_);
  and (_10247_, _10246_, _05332_);
  or (_10248_, _10234_, _05332_);
  nor (_10249_, _10248_, _10182_);
  nor (_10250_, _10249_, _10247_);
  nor (_10251_, _10250_, _03243_);
  nor (_10252_, _10181_, _04888_);
  or (_10253_, _10252_, _03244_);
  nor (_10254_, _10253_, _10195_);
  or (_10255_, _10254_, _02654_);
  nor (_10256_, _10255_, _10251_);
  nor (_10257_, _07967_, _07143_);
  nor (_10258_, _10257_, _10181_);
  and (_10259_, _10258_, _02654_);
  nor (_10260_, _10259_, _10256_);
  and (_10261_, _10260_, _05883_);
  nor (_10262_, _08109_, _07143_);
  nor (_10263_, _10262_, _10181_);
  nor (_10264_, _10263_, _05883_);
  or (_10265_, _10264_, _10261_);
  and (_10266_, _10265_, _03124_);
  nor (_10267_, _10183_, _03124_);
  nor (_10268_, _10267_, _02650_);
  not (_10269_, _10268_);
  nor (_10270_, _10269_, _10266_);
  nor (_10271_, _10181_, _03122_);
  nor (_10272_, _10271_, _10270_);
  and (_10273_, _10272_, _03513_);
  nor (_10274_, _10273_, _10184_);
  nand (_10275_, _10274_, _27788_);
  or (_10276_, _27788_, \oc8051_golden_model_1.IE [0]);
  and (_10277_, _10276_, _27053_);
  and (_28801_, _10277_, _10275_);
  not (_10278_, \oc8051_golden_model_1.IE [1]);
  nor (_10279_, _04629_, _10278_);
  and (_10280_, _04629_, _04218_);
  or (_10281_, _10280_, _10279_);
  and (_10282_, _10281_, _05959_);
  nor (_10283_, _08246_, _07180_);
  nor (_10284_, _05433_, _10278_);
  or (_10285_, _10284_, _03141_);
  or (_10286_, _10285_, _10283_);
  nor (_10287_, _04629_, \oc8051_golden_model_1.IE [1]);
  and (_10288_, _08209_, _04629_);
  nor (_10289_, _10288_, _10287_);
  nor (_10290_, _10289_, _02662_);
  and (_10291_, _04629_, _08322_);
  nor (_10292_, _10291_, _10287_);
  and (_10293_, _10292_, _04505_);
  nor (_10294_, _04505_, _10278_);
  or (_10295_, _10294_, _02661_);
  nor (_10296_, _10295_, _10293_);
  or (_10297_, _10296_, _06504_);
  nor (_10298_, _10297_, _10290_);
  nor (_10299_, _07143_, _03777_);
  nor (_10300_, _10299_, _10279_);
  nor (_10301_, _10300_, _03365_);
  and (_10302_, _08213_, _05433_);
  nor (_10303_, _10302_, _10284_);
  nor (_10304_, _10303_, _03390_);
  nor (_10305_, _10304_, _10301_);
  nand (_10306_, _10305_, _03179_);
  or (_10307_, _10306_, _10298_);
  or (_10308_, _10292_, _03179_);
  and (_10309_, _10308_, _10307_);
  and (_10310_, _10309_, _03177_);
  and (_10311_, _08200_, _05433_);
  nor (_10312_, _10311_, _10284_);
  nor (_10313_, _10312_, _03177_);
  or (_10314_, _10313_, _10310_);
  and (_10315_, _10314_, _05168_);
  nor (_10316_, _10284_, _08228_);
  or (_10317_, _10316_, _05168_);
  nor (_10318_, _10317_, _10303_);
  or (_10319_, _10318_, _03140_);
  or (_10320_, _10319_, _10315_);
  and (_10321_, _10320_, _10286_);
  nor (_10322_, _10321_, _05949_);
  and (_10323_, _10300_, _05949_);
  or (_10324_, _10323_, _05959_);
  nor (_10325_, _10324_, _10322_);
  or (_10326_, _10325_, _10282_);
  and (_10327_, _10326_, _03139_);
  nor (_10328_, _08307_, _07143_);
  nor (_10329_, _10328_, _10279_);
  nor (_10330_, _10329_, _03139_);
  nor (_10331_, _10330_, _10327_);
  nor (_10332_, _10331_, _06549_);
  and (_10333_, _04629_, _03016_);
  not (_10334_, _10333_);
  nor (_10335_, _10287_, _05245_);
  and (_10336_, _10335_, _10334_);
  nor (_10337_, _10336_, _10332_);
  not (_10338_, _10279_);
  nand (_10339_, _08185_, _04629_);
  and (_10340_, _10339_, _10338_);
  or (_10341_, _10340_, _05305_);
  and (_10342_, _10341_, _10337_);
  nor (_10343_, _10342_, _03251_);
  not (_10344_, _10287_);
  nor (_10345_, _08325_, _07143_);
  nor (_10346_, _10345_, _03252_);
  and (_10347_, _10346_, _10344_);
  nor (_10348_, _10347_, _10343_);
  nor (_10349_, _10348_, _02669_);
  nor (_10350_, _08184_, _07143_);
  nor (_10351_, _10350_, _05332_);
  and (_10352_, _10351_, _10344_);
  nor (_10353_, _10352_, _10349_);
  nor (_10354_, _10353_, _03243_);
  and (_10355_, _10338_, _04835_);
  nor (_10356_, _10355_, _03244_);
  and (_10357_, _10356_, _10292_);
  nor (_10358_, _10357_, _10354_);
  nor (_10359_, _10358_, _03241_);
  and (_10360_, _10333_, _04835_);
  nor (_10361_, _10360_, _05357_);
  nand (_10362_, _10291_, _04835_);
  and (_10363_, _10362_, _03239_);
  or (_10364_, _10363_, _10361_);
  and (_10365_, _10364_, _10344_);
  or (_10366_, _10365_, _03123_);
  nor (_10367_, _10366_, _10359_);
  nor (_10368_, _10289_, _03124_);
  or (_10369_, _10368_, _02650_);
  nor (_10370_, _10369_, _10367_);
  nor (_10371_, _10312_, _03122_);
  or (_10372_, _10371_, _03121_);
  nor (_10373_, _10372_, _10370_);
  nor (_10374_, _10288_, _10279_);
  and (_10375_, _10374_, _03121_);
  nor (_10376_, _10375_, _10373_);
  or (_10377_, _10376_, _27789_);
  or (_10378_, _27788_, \oc8051_golden_model_1.IE [1]);
  and (_10379_, _10378_, _27053_);
  and (_28802_, _10379_, _10377_);
  not (_10380_, \oc8051_golden_model_1.IE [2]);
  nor (_10381_, _04629_, _10380_);
  and (_10382_, _04629_, _06009_);
  nor (_10383_, _10382_, _10381_);
  and (_10384_, _10383_, _02575_);
  nor (_10385_, _07143_, _03644_);
  nor (_10386_, _10385_, _10381_);
  and (_10387_, _10386_, _05949_);
  nor (_10388_, _08420_, _07143_);
  nor (_10389_, _10388_, _10381_);
  and (_10390_, _10389_, _02661_);
  and (_10391_, _04629_, \oc8051_golden_model_1.ACC [2]);
  nor (_10392_, _10391_, _10381_);
  nor (_10393_, _10392_, _05903_);
  nor (_10394_, _04505_, _10380_);
  or (_10395_, _10394_, _02661_);
  nor (_10396_, _10395_, _10393_);
  or (_10397_, _10396_, _06504_);
  nor (_10398_, _10397_, _10390_);
  nor (_10399_, _10386_, _03365_);
  nor (_10400_, _05433_, _10380_);
  and (_10401_, _08406_, _05433_);
  nor (_10402_, _10401_, _10400_);
  nor (_10403_, _10402_, _03390_);
  nor (_10404_, _10403_, _10399_);
  nand (_10405_, _10404_, _03179_);
  or (_10406_, _10405_, _10398_);
  nand (_10407_, _10392_, _03168_);
  and (_10408_, _10407_, _10406_);
  nor (_10409_, _10408_, _03176_);
  and (_10410_, _08404_, _05433_);
  nor (_10411_, _10410_, _10400_);
  and (_10412_, _10411_, _03176_);
  or (_10413_, _10412_, _03144_);
  nor (_10414_, _10413_, _10409_);
  nor (_10415_, _10400_, _08446_);
  or (_10416_, _10415_, _05168_);
  nor (_10417_, _10416_, _10402_);
  or (_10418_, _10417_, _10414_);
  and (_10419_, _10418_, _03141_);
  nor (_10420_, _08465_, _07180_);
  nor (_10421_, _10400_, _10420_);
  nor (_10422_, _10421_, _03141_);
  or (_10423_, _10422_, _05949_);
  nor (_10424_, _10423_, _10419_);
  nor (_10425_, _10424_, _10387_);
  nor (_10426_, _10425_, _05959_);
  and (_10427_, _04629_, _04170_);
  nor (_10428_, _10381_, _05963_);
  not (_10429_, _10428_);
  nor (_10430_, _10429_, _10427_);
  or (_10431_, _10430_, _02024_);
  nor (_10432_, _10431_, _10426_);
  nor (_10433_, _08522_, _07143_);
  nor (_10434_, _10433_, _10381_);
  nor (_10435_, _10434_, _03139_);
  or (_10436_, _10435_, _02575_);
  nor (_10437_, _10436_, _10432_);
  nor (_10438_, _10437_, _10384_);
  or (_10439_, _10438_, _02656_);
  and (_10440_, _08537_, _04629_);
  or (_10441_, _10440_, _10381_);
  or (_10442_, _10441_, _05305_);
  and (_10443_, _10442_, _03252_);
  and (_10444_, _10443_, _10439_);
  and (_10445_, _08387_, _04629_);
  nor (_10446_, _10445_, _10381_);
  nor (_10447_, _10446_, _03252_);
  nor (_10448_, _10447_, _10444_);
  nor (_10449_, _10448_, _02669_);
  nor (_10450_, _10381_, _06121_);
  not (_10451_, _10450_);
  nor (_10452_, _10383_, _05332_);
  and (_10453_, _10452_, _10451_);
  nor (_10454_, _10453_, _10449_);
  nor (_10455_, _10454_, _03243_);
  or (_10456_, _10450_, _03244_);
  nor (_10457_, _10456_, _10392_);
  or (_10458_, _10457_, _02654_);
  nor (_10459_, _10458_, _10455_);
  nor (_10460_, _08536_, _07143_);
  nor (_10461_, _10460_, _10381_);
  and (_10462_, _10461_, _02654_);
  nor (_10463_, _10462_, _10459_);
  and (_10464_, _10463_, _05883_);
  nor (_10465_, _08386_, _07143_);
  nor (_10466_, _10465_, _10381_);
  nor (_10467_, _10466_, _05883_);
  or (_10468_, _10467_, _10464_);
  and (_10469_, _10468_, _03124_);
  nor (_10470_, _10389_, _03124_);
  or (_10471_, _10470_, _02650_);
  or (_10472_, _10471_, _10469_);
  nand (_10473_, _10411_, _02650_);
  and (_10474_, _10473_, _10472_);
  nor (_10475_, _10474_, _03121_);
  and (_10476_, _08596_, _04629_);
  nor (_10477_, _10476_, _10381_);
  and (_10478_, _10477_, _03121_);
  nor (_10479_, _10478_, _10475_);
  or (_10480_, _10479_, _27789_);
  or (_10481_, _27788_, \oc8051_golden_model_1.IE [2]);
  and (_10482_, _10481_, _27053_);
  and (_28803_, _10482_, _10480_);
  not (_10483_, \oc8051_golden_model_1.IE [3]);
  nor (_10484_, _04629_, _10483_);
  and (_10485_, _04629_, _05986_);
  nor (_10486_, _10485_, _10484_);
  and (_10487_, _10486_, _02575_);
  nor (_10488_, _07143_, _03859_);
  nor (_10489_, _10488_, _10484_);
  and (_10490_, _10489_, _05949_);
  nor (_10491_, _08627_, _07180_);
  nor (_10492_, _05433_, _10483_);
  or (_10493_, _10492_, _03141_);
  or (_10494_, _10493_, _10491_);
  nor (_10495_, _08646_, _07143_);
  nor (_10496_, _10495_, _10484_);
  and (_10497_, _10496_, _02661_);
  and (_10498_, _04629_, \oc8051_golden_model_1.ACC [3]);
  nor (_10499_, _10498_, _10484_);
  nor (_10500_, _10499_, _05903_);
  nor (_10501_, _04505_, _10483_);
  or (_10502_, _10501_, _02661_);
  nor (_10503_, _10502_, _10500_);
  or (_10504_, _10503_, _06504_);
  nor (_10505_, _10504_, _10497_);
  nor (_10506_, _10489_, _03365_);
  and (_10507_, _08642_, _05433_);
  nor (_10508_, _10507_, _10492_);
  nor (_10509_, _10508_, _03390_);
  nor (_10510_, _10509_, _10506_);
  nand (_10511_, _10510_, _03179_);
  or (_10512_, _10511_, _10505_);
  nand (_10513_, _10499_, _03168_);
  and (_10514_, _10513_, _10512_);
  and (_10515_, _10514_, _03177_);
  and (_10516_, _08640_, _05433_);
  nor (_10517_, _10516_, _10492_);
  nor (_10518_, _10517_, _03177_);
  or (_10519_, _10518_, _10515_);
  and (_10520_, _10519_, _05168_);
  nor (_10521_, _10492_, _08671_);
  or (_10522_, _10508_, _05168_);
  nor (_10523_, _10522_, _10521_);
  or (_10524_, _10523_, _03140_);
  or (_10525_, _10524_, _10520_);
  and (_10526_, _10525_, _10494_);
  nor (_10527_, _10526_, _05949_);
  nor (_10528_, _10527_, _10490_);
  nor (_10529_, _10528_, _05959_);
  and (_10530_, _04629_, _04120_);
  nor (_10531_, _10484_, _05963_);
  not (_10532_, _10531_);
  nor (_10533_, _10532_, _10530_);
  or (_10534_, _10533_, _02024_);
  nor (_10535_, _10534_, _10529_);
  nor (_10536_, _08744_, _07143_);
  nor (_10537_, _10536_, _10484_);
  nor (_10538_, _10537_, _03139_);
  or (_10539_, _10538_, _02575_);
  nor (_10540_, _10539_, _10535_);
  nor (_10541_, _10540_, _10487_);
  or (_10542_, _10541_, _02656_);
  and (_10543_, _08622_, _04629_);
  or (_10544_, _10543_, _10484_);
  or (_10545_, _10544_, _05305_);
  and (_10546_, _10545_, _03252_);
  and (_10547_, _10546_, _10542_);
  and (_10548_, _08618_, _04629_);
  nor (_10549_, _10548_, _10484_);
  nor (_10550_, _10549_, _03252_);
  nor (_10551_, _10550_, _10547_);
  nor (_10552_, _10551_, _02669_);
  nor (_10553_, _10484_, _06120_);
  not (_10554_, _10553_);
  nor (_10555_, _10486_, _05332_);
  and (_10556_, _10555_, _10554_);
  nor (_10557_, _10556_, _10552_);
  nor (_10558_, _10557_, _03243_);
  or (_10559_, _10553_, _03244_);
  nor (_10560_, _10559_, _10499_);
  or (_10561_, _10560_, _02654_);
  nor (_10562_, _10561_, _10558_);
  nor (_10563_, _08621_, _07143_);
  nor (_10564_, _10563_, _10484_);
  and (_10565_, _10564_, _02654_);
  nor (_10566_, _10565_, _10562_);
  and (_10567_, _10566_, _05883_);
  nor (_10568_, _08617_, _07143_);
  nor (_10569_, _10568_, _10484_);
  nor (_10570_, _10569_, _05883_);
  or (_10571_, _10570_, _10567_);
  and (_10572_, _10571_, _03124_);
  nor (_10573_, _10496_, _03124_);
  or (_10574_, _10573_, _02650_);
  or (_10575_, _10574_, _10572_);
  nand (_10576_, _10517_, _02650_);
  and (_10577_, _10576_, _10575_);
  nor (_10578_, _10577_, _03121_);
  and (_10579_, _08807_, _04629_);
  nor (_10580_, _10579_, _10484_);
  and (_10581_, _10580_, _03121_);
  nor (_10582_, _10581_, _10578_);
  or (_10583_, _10582_, _27789_);
  or (_10584_, _27788_, \oc8051_golden_model_1.IE [3]);
  and (_10585_, _10584_, _27053_);
  and (_28804_, _10585_, _10583_);
  not (_10586_, \oc8051_golden_model_1.IE [4]);
  nor (_10587_, _04629_, _10586_);
  and (_10588_, _04629_, _05974_);
  nor (_10589_, _10588_, _10587_);
  and (_10590_, _10589_, _02575_);
  nor (_10591_, _07143_, _04325_);
  nor (_10592_, _10591_, _10587_);
  and (_10593_, _10592_, _05949_);
  nor (_10594_, _05433_, _10586_);
  nor (_10595_, _10594_, _08889_);
  and (_10596_, _08869_, _05433_);
  nor (_10597_, _10596_, _10594_);
  or (_10598_, _10597_, _05168_);
  nor (_10599_, _10598_, _10595_);
  nor (_10600_, _08838_, _07143_);
  nor (_10601_, _10600_, _10587_);
  and (_10602_, _10601_, _02661_);
  and (_10603_, _04629_, \oc8051_golden_model_1.ACC [4]);
  nor (_10604_, _10603_, _10587_);
  nor (_10605_, _10604_, _05903_);
  nor (_10606_, _04505_, _10586_);
  or (_10607_, _10606_, _02661_);
  nor (_10608_, _10607_, _10605_);
  or (_10609_, _10608_, _06504_);
  nor (_10610_, _10609_, _10602_);
  nor (_10611_, _10592_, _03365_);
  nor (_10612_, _10597_, _03390_);
  nor (_10613_, _10612_, _10611_);
  nand (_10614_, _10613_, _03179_);
  or (_10615_, _10614_, _10610_);
  nand (_10616_, _10604_, _03168_);
  and (_10617_, _10616_, _10615_);
  and (_10618_, _10617_, _03177_);
  and (_10619_, _08880_, _05433_);
  nor (_10620_, _10619_, _10594_);
  nor (_10621_, _10620_, _03177_);
  or (_10622_, _10621_, _10618_);
  and (_10623_, _10622_, _05168_);
  nor (_10624_, _10623_, _10599_);
  nor (_10625_, _10624_, _03140_);
  nor (_10626_, _08908_, _07180_);
  nor (_10627_, _10626_, _10594_);
  nor (_10628_, _10627_, _03141_);
  nor (_10629_, _10628_, _05949_);
  not (_10630_, _10629_);
  nor (_10631_, _10630_, _10625_);
  nor (_10632_, _10631_, _10593_);
  nor (_10633_, _10632_, _05959_);
  and (_10634_, _04629_, _04012_);
  nor (_10635_, _10587_, _05963_);
  not (_10636_, _10635_);
  nor (_10637_, _10636_, _10634_);
  or (_10638_, _10637_, _02024_);
  nor (_10639_, _10638_, _10633_);
  nor (_10640_, _08967_, _07143_);
  nor (_10641_, _10640_, _10587_);
  nor (_10642_, _10641_, _03139_);
  or (_10643_, _10642_, _02575_);
  nor (_10644_, _10643_, _10639_);
  nor (_10645_, _10644_, _10590_);
  or (_10646_, _10645_, _02656_);
  and (_10647_, _08982_, _04629_);
  or (_10648_, _10647_, _10587_);
  or (_10649_, _10648_, _05305_);
  and (_10650_, _10649_, _03252_);
  and (_10651_, _10650_, _10646_);
  and (_10652_, _08830_, _04629_);
  nor (_10653_, _10652_, _10587_);
  nor (_10654_, _10653_, _03252_);
  nor (_10655_, _10654_, _10651_);
  nor (_10656_, _10655_, _02669_);
  nor (_10657_, _10587_, _09034_);
  not (_10658_, _10657_);
  nor (_10659_, _10589_, _05332_);
  and (_10660_, _10659_, _10658_);
  nor (_10661_, _10660_, _10656_);
  nor (_10662_, _10661_, _03243_);
  or (_10663_, _10657_, _03244_);
  nor (_10664_, _10663_, _10604_);
  or (_10665_, _10664_, _02654_);
  nor (_10666_, _10665_, _10662_);
  nor (_10667_, _08981_, _07143_);
  nor (_10668_, _10667_, _10587_);
  and (_10669_, _10668_, _02654_);
  nor (_10670_, _10669_, _10666_);
  and (_10671_, _10670_, _05883_);
  nor (_10672_, _08828_, _07143_);
  nor (_10673_, _10672_, _10587_);
  nor (_10674_, _10673_, _05883_);
  or (_10675_, _10674_, _10671_);
  and (_10676_, _10675_, _03124_);
  nor (_10677_, _10601_, _03124_);
  or (_10678_, _10677_, _02650_);
  or (_10679_, _10678_, _10676_);
  nand (_10680_, _10620_, _02650_);
  and (_10681_, _10680_, _10679_);
  nor (_10682_, _10681_, _03121_);
  and (_10683_, _09037_, _04629_);
  nor (_10684_, _10683_, _10587_);
  and (_10685_, _10684_, _03121_);
  nor (_10686_, _10685_, _10682_);
  or (_10687_, _10686_, _27789_);
  or (_10688_, _27788_, \oc8051_golden_model_1.IE [4]);
  and (_10689_, _10688_, _27053_);
  and (_28805_, _10689_, _10687_);
  not (_10690_, \oc8051_golden_model_1.IE [5]);
  nor (_10691_, _04629_, _10690_);
  and (_10692_, _04629_, _06036_);
  nor (_10693_, _10692_, _10691_);
  and (_10694_, _10693_, _02575_);
  nor (_10695_, _07143_, _04480_);
  nor (_10696_, _10695_, _10691_);
  and (_10697_, _10696_, _05949_);
  and (_10698_, _04629_, \oc8051_golden_model_1.ACC [5]);
  nor (_10699_, _10698_, _10691_);
  and (_10700_, _10699_, _03168_);
  nor (_10701_, _09087_, _07143_);
  nor (_10702_, _10701_, _10691_);
  and (_10703_, _10702_, _02661_);
  nor (_10704_, _10699_, _05903_);
  nor (_10705_, _04505_, _10690_);
  or (_10706_, _10705_, _02661_);
  nor (_10707_, _10706_, _10704_);
  or (_10708_, _10707_, _06504_);
  nor (_10709_, _10708_, _10703_);
  nor (_10710_, _10696_, _03365_);
  nor (_10711_, _10710_, _10709_);
  nor (_10712_, _05433_, _10690_);
  and (_10713_, _09072_, _05433_);
  nor (_10714_, _10713_, _10712_);
  nor (_10715_, _10714_, _03390_);
  nor (_10716_, _10715_, _03168_);
  and (_10717_, _10716_, _10711_);
  nor (_10718_, _10717_, _10700_);
  and (_10719_, _10718_, _03177_);
  and (_10720_, _09099_, _05433_);
  nor (_10721_, _10720_, _10712_);
  nor (_10722_, _10721_, _03177_);
  or (_10723_, _10722_, _10719_);
  and (_10724_, _10723_, _05168_);
  and (_10725_, _09108_, _05433_);
  nor (_10726_, _10725_, _10712_);
  nor (_10727_, _10726_, _05168_);
  nor (_10728_, _10727_, _10724_);
  nor (_10729_, _10728_, _03140_);
  nor (_10730_, _09059_, _07180_);
  nor (_10731_, _10730_, _10712_);
  nor (_10732_, _10731_, _03141_);
  nor (_10733_, _10732_, _05949_);
  not (_10734_, _10733_);
  nor (_10735_, _10734_, _10729_);
  nor (_10736_, _10735_, _10697_);
  nor (_10737_, _10736_, _05959_);
  and (_10738_, _04629_, _03904_);
  nor (_10739_, _10691_, _05963_);
  not (_10740_, _10739_);
  nor (_10741_, _10740_, _10738_);
  or (_10742_, _10741_, _02024_);
  nor (_10743_, _10742_, _10737_);
  nor (_10744_, _09180_, _07143_);
  nor (_10745_, _10744_, _10691_);
  nor (_10746_, _10745_, _03139_);
  or (_10747_, _10746_, _02575_);
  nor (_10748_, _10747_, _10743_);
  nor (_10749_, _10748_, _10694_);
  or (_10750_, _10749_, _02656_);
  and (_10751_, _09195_, _04629_);
  or (_10752_, _10751_, _10691_);
  or (_10753_, _10752_, _05305_);
  and (_10754_, _10753_, _03252_);
  and (_10755_, _10754_, _10750_);
  and (_10756_, _09055_, _04629_);
  nor (_10757_, _10756_, _10691_);
  nor (_10758_, _10757_, _03252_);
  nor (_10759_, _10758_, _10755_);
  nor (_10760_, _10759_, _02669_);
  not (_10761_, _10691_);
  and (_10762_, _10761_, _04787_);
  not (_10763_, _10762_);
  nor (_10764_, _10693_, _05332_);
  and (_10765_, _10764_, _10763_);
  nor (_10766_, _10765_, _10760_);
  nor (_10767_, _10766_, _03243_);
  or (_10768_, _10762_, _03244_);
  nor (_10769_, _10768_, _10699_);
  or (_10770_, _10769_, _02654_);
  nor (_10771_, _10770_, _10767_);
  nor (_10772_, _09194_, _07143_);
  nor (_10773_, _10772_, _10691_);
  and (_10774_, _10773_, _02654_);
  nor (_10775_, _10774_, _10771_);
  and (_10776_, _10775_, _05883_);
  nor (_10777_, _09054_, _07143_);
  nor (_10778_, _10777_, _10691_);
  nor (_10779_, _10778_, _05883_);
  or (_10780_, _10779_, _10776_);
  and (_10781_, _10780_, _03124_);
  nor (_10782_, _10702_, _03124_);
  or (_10783_, _10782_, _02650_);
  or (_10784_, _10783_, _10781_);
  nand (_10785_, _10721_, _02650_);
  and (_10786_, _10785_, _10784_);
  nor (_10787_, _10786_, _03121_);
  and (_10788_, _09248_, _04629_);
  nor (_10789_, _10788_, _10691_);
  and (_10790_, _10789_, _03121_);
  nor (_10791_, _10790_, _10787_);
  or (_10792_, _10791_, _27789_);
  or (_10793_, _27788_, \oc8051_golden_model_1.IE [5]);
  and (_10794_, _10793_, _27053_);
  and (_28808_, _10794_, _10792_);
  not (_10795_, \oc8051_golden_model_1.IE [6]);
  nor (_10796_, _04629_, _10795_);
  and (_10797_, _04629_, _03960_);
  or (_10798_, _10797_, _10796_);
  and (_10799_, _10798_, _05959_);
  nor (_10800_, _05433_, _10795_);
  not (_10801_, _10800_);
  and (_10802_, _10801_, _09320_);
  and (_10803_, _09305_, _05433_);
  nor (_10804_, _10803_, _10800_);
  or (_10805_, _10804_, _05168_);
  nor (_10806_, _10805_, _10802_);
  nor (_10807_, _09301_, _07143_);
  nor (_10808_, _10807_, _10796_);
  and (_10809_, _10808_, _02661_);
  and (_10810_, _04629_, \oc8051_golden_model_1.ACC [6]);
  nor (_10811_, _10810_, _10796_);
  nor (_10812_, _10811_, _05903_);
  nor (_10813_, _04505_, _10795_);
  or (_10814_, _10813_, _02661_);
  nor (_10815_, _10814_, _10812_);
  or (_10816_, _10815_, _06504_);
  nor (_10817_, _10816_, _10809_);
  nor (_10818_, _07143_, _04373_);
  nor (_10819_, _10818_, _10796_);
  nor (_10820_, _10819_, _03365_);
  nor (_10821_, _10804_, _03390_);
  nor (_10822_, _10821_, _10820_);
  nand (_10823_, _10822_, _03179_);
  or (_10824_, _10823_, _10817_);
  nand (_10825_, _10811_, _03168_);
  and (_10826_, _10825_, _10824_);
  and (_10827_, _10826_, _03177_);
  and (_10828_, _09286_, _05433_);
  nor (_10829_, _10828_, _10800_);
  nor (_10830_, _10829_, _03177_);
  or (_10831_, _10830_, _10827_);
  and (_10832_, _10831_, _05168_);
  nor (_10833_, _10832_, _10806_);
  nor (_10834_, _10833_, _03140_);
  nor (_10835_, _09272_, _07180_);
  nor (_10836_, _10835_, _10800_);
  nor (_10837_, _10836_, _03141_);
  nor (_10838_, _10837_, _05949_);
  not (_10839_, _10838_);
  nor (_10840_, _10839_, _10834_);
  and (_10841_, _10819_, _05949_);
  or (_10842_, _10841_, _05959_);
  nor (_10843_, _10842_, _10840_);
  or (_10844_, _10843_, _10799_);
  and (_10845_, _10844_, _03139_);
  and (_10846_, _09388_, _04629_);
  nor (_10847_, _10846_, _10796_);
  nor (_10848_, _10847_, _03139_);
  or (_10849_, _10848_, _06549_);
  or (_10850_, _10849_, _10845_);
  and (_10851_, _09404_, _04629_);
  or (_10852_, _10796_, _05305_);
  or (_10853_, _10852_, _10851_);
  and (_10854_, _04629_, _09395_);
  nor (_10855_, _10854_, _10796_);
  and (_10856_, _10855_, _02575_);
  nor (_10857_, _10856_, _03251_);
  and (_10858_, _10857_, _10853_);
  and (_10859_, _10858_, _10850_);
  and (_10860_, _09268_, _04629_);
  nor (_10861_, _10860_, _10796_);
  nor (_10862_, _10861_, _03252_);
  nor (_10863_, _10862_, _10859_);
  nor (_10864_, _10863_, _02669_);
  nor (_10865_, _10796_, _06119_);
  not (_10866_, _10865_);
  nor (_10867_, _10855_, _05332_);
  and (_10868_, _10867_, _10866_);
  nor (_10869_, _10868_, _10864_);
  nor (_10870_, _10869_, _03243_);
  or (_10871_, _10865_, _03244_);
  nor (_10872_, _10871_, _10811_);
  or (_10873_, _10872_, _02654_);
  nor (_10874_, _10873_, _10870_);
  nor (_10875_, _09403_, _07143_);
  nor (_10876_, _10875_, _10796_);
  and (_10877_, _10876_, _02654_);
  nor (_10878_, _10877_, _10874_);
  and (_10879_, _10878_, _05883_);
  nor (_10880_, _09267_, _07143_);
  nor (_10881_, _10880_, _10796_);
  nor (_10882_, _10881_, _05883_);
  or (_10883_, _10882_, _10879_);
  and (_10884_, _10883_, _03124_);
  nor (_10885_, _10808_, _03124_);
  or (_10886_, _10885_, _02650_);
  or (_10887_, _10886_, _10884_);
  nand (_10888_, _10829_, _02650_);
  and (_10889_, _10888_, _10887_);
  nor (_10890_, _10889_, _03121_);
  and (_10891_, _09456_, _04629_);
  nor (_10892_, _10891_, _10796_);
  and (_10893_, _10892_, _03121_);
  nor (_10894_, _10893_, _10890_);
  or (_10895_, _10894_, _27789_);
  or (_10896_, _27788_, \oc8051_golden_model_1.IE [6]);
  and (_10897_, _10896_, _27053_);
  and (_28809_, _10897_, _10895_);
  not (_10898_, \oc8051_golden_model_1.IP [0]);
  nor (_10899_, _04581_, _10898_);
  nor (_10900_, _04888_, _07034_);
  nor (_10901_, _10900_, _10899_);
  nor (_10902_, _10901_, _03513_);
  and (_10903_, _04581_, _05996_);
  nor (_10904_, _10903_, _10899_);
  nor (_10905_, _10904_, _05332_);
  not (_10906_, _10905_);
  nor (_10907_, _10906_, _10900_);
  and (_10908_, _04581_, _04268_);
  nor (_10909_, _10899_, _05963_);
  not (_10910_, _10909_);
  nor (_10911_, _10910_, _10908_);
  nor (_10912_, _05425_, _10898_);
  and (_10913_, _07997_, _05425_);
  nor (_10914_, _10913_, _10912_);
  nor (_10915_, _10914_, _03390_);
  and (_10916_, _10901_, _02661_);
  and (_10917_, _04581_, \oc8051_golden_model_1.ACC [0]);
  nor (_10918_, _10917_, _10899_);
  nor (_10919_, _10918_, _05903_);
  nor (_10920_, _04505_, _10898_);
  or (_10921_, _10920_, _02661_);
  nor (_10922_, _10921_, _10919_);
  or (_10923_, _10922_, _06504_);
  nor (_10924_, _10923_, _10916_);
  and (_10925_, _04581_, _03716_);
  nor (_10926_, _10925_, _10899_);
  nor (_10927_, _10926_, _03365_);
  or (_10928_, _10927_, _03168_);
  or (_10929_, _10928_, _10924_);
  nor (_10930_, _10929_, _10915_);
  and (_10931_, _10918_, _03168_);
  nor (_10932_, _10931_, _03176_);
  not (_10933_, _10932_);
  nor (_10934_, _10933_, _10930_);
  and (_10935_, _10899_, _03176_);
  or (_10936_, _10935_, _10934_);
  and (_10937_, _10936_, _05168_);
  nor (_10938_, _10901_, _05168_);
  or (_10939_, _10938_, _10937_);
  nor (_10940_, _10939_, _03140_);
  nor (_10941_, _08035_, _07071_);
  or (_10942_, _10912_, _03141_);
  nor (_10943_, _10942_, _10941_);
  or (_10944_, _10943_, _05949_);
  or (_10945_, _10944_, _10940_);
  or (_10946_, _10926_, _06673_);
  and (_10947_, _10946_, _05963_);
  and (_10948_, _10947_, _10945_);
  nor (_10949_, _10948_, _10911_);
  nor (_10950_, _10949_, _02024_);
  nor (_10951_, _08093_, _07034_);
  or (_10952_, _10899_, _03139_);
  nor (_10953_, _10952_, _10951_);
  or (_10954_, _10953_, _02575_);
  nor (_10955_, _10954_, _10950_);
  nand (_10956_, _10904_, _05305_);
  and (_10957_, _10956_, _06549_);
  nor (_10958_, _10957_, _10955_);
  and (_10959_, _07968_, _04581_);
  nor (_10960_, _10959_, _10899_);
  and (_10961_, _10960_, _02656_);
  nor (_10962_, _10961_, _10958_);
  and (_10963_, _10962_, _03252_);
  and (_10964_, _08110_, _04581_);
  nor (_10965_, _10964_, _10899_);
  nor (_10966_, _10965_, _03252_);
  or (_10967_, _10966_, _10963_);
  and (_10968_, _10967_, _05332_);
  nor (_10969_, _10968_, _10907_);
  nor (_10970_, _10969_, _03243_);
  nor (_10971_, _10899_, _04888_);
  or (_10972_, _10971_, _03244_);
  nor (_10973_, _10972_, _10918_);
  or (_10974_, _10973_, _02654_);
  nor (_10975_, _10974_, _10970_);
  nor (_10976_, _07967_, _07034_);
  nor (_10977_, _10976_, _10899_);
  and (_10978_, _10977_, _02654_);
  nor (_10979_, _10978_, _10975_);
  and (_10980_, _10979_, _05883_);
  nor (_10981_, _08109_, _07034_);
  nor (_10982_, _10981_, _10899_);
  nor (_10983_, _10982_, _05883_);
  or (_10984_, _10983_, _10980_);
  and (_10985_, _10984_, _03124_);
  nor (_10986_, _10901_, _03124_);
  nor (_10987_, _10986_, _02650_);
  not (_10988_, _10987_);
  nor (_10989_, _10988_, _10985_);
  nor (_10990_, _10899_, _03122_);
  nor (_10991_, _10990_, _10989_);
  and (_10992_, _10991_, _03513_);
  nor (_10993_, _10992_, _10902_);
  nand (_10994_, _10993_, _27788_);
  or (_10995_, _27788_, \oc8051_golden_model_1.IP [0]);
  and (_10996_, _10995_, _27053_);
  and (_28810_, _10996_, _10994_);
  nor (_10997_, _04581_, \oc8051_golden_model_1.IP [1]);
  not (_10998_, _10997_);
  nor (_10999_, _08325_, _07034_);
  nor (_11000_, _10999_, _03252_);
  and (_11001_, _11000_, _10998_);
  not (_11002_, \oc8051_golden_model_1.IP [1]);
  nor (_11003_, _04581_, _11002_);
  and (_11004_, _04581_, _04218_);
  or (_11005_, _11004_, _11003_);
  and (_11006_, _11005_, _05959_);
  nor (_11007_, _08246_, _07071_);
  nor (_11008_, _05425_, _11002_);
  or (_11009_, _11008_, _03141_);
  or (_11010_, _11009_, _11007_);
  and (_11011_, _08209_, _04581_);
  nor (_11012_, _11011_, _10997_);
  nor (_11013_, _11012_, _02662_);
  and (_11014_, _04581_, _08322_);
  nor (_11015_, _11014_, _10997_);
  and (_11016_, _11015_, _04505_);
  nor (_11017_, _04505_, _11002_);
  or (_11018_, _11017_, _02661_);
  nor (_11019_, _11018_, _11016_);
  or (_11020_, _11019_, _06504_);
  nor (_11021_, _11020_, _11013_);
  nor (_11022_, _07034_, _03777_);
  nor (_11023_, _11022_, _11003_);
  nor (_11024_, _11023_, _03365_);
  and (_11025_, _08213_, _05425_);
  nor (_11026_, _11025_, _11008_);
  nor (_11027_, _11026_, _03390_);
  nor (_11028_, _11027_, _11024_);
  nand (_11029_, _11028_, _03179_);
  or (_11030_, _11029_, _11021_);
  or (_11031_, _11015_, _03179_);
  and (_11032_, _11031_, _11030_);
  and (_11033_, _11032_, _03177_);
  and (_11034_, _08200_, _05425_);
  nor (_11035_, _11034_, _11008_);
  nor (_11036_, _11035_, _03177_);
  or (_11037_, _11036_, _11033_);
  and (_11038_, _11037_, _05168_);
  nor (_11039_, _11008_, _08228_);
  or (_11040_, _11039_, _05168_);
  nor (_11041_, _11040_, _11026_);
  or (_11042_, _11041_, _03140_);
  or (_11043_, _11042_, _11038_);
  and (_11044_, _11043_, _11010_);
  nor (_11045_, _11044_, _05949_);
  and (_11046_, _11023_, _05949_);
  or (_11047_, _11046_, _05959_);
  nor (_11048_, _11047_, _11045_);
  or (_11049_, _11048_, _11006_);
  and (_11050_, _11049_, _03139_);
  nor (_11051_, _08307_, _07034_);
  nor (_11052_, _11051_, _11003_);
  nor (_11053_, _11052_, _03139_);
  nor (_11054_, _11053_, _11050_);
  nor (_11055_, _11054_, _06549_);
  nor (_11056_, _08185_, _07034_);
  nor (_11057_, _11056_, _05305_);
  and (_11058_, _04581_, _03016_);
  nor (_11059_, _11058_, _05245_);
  nor (_11060_, _11059_, _11057_);
  nor (_11061_, _11060_, _10997_);
  nor (_11062_, _11061_, _11055_);
  nor (_11063_, _11062_, _03251_);
  nor (_11064_, _11063_, _11001_);
  nor (_11065_, _11064_, _02669_);
  nor (_11066_, _08184_, _07034_);
  nor (_11067_, _11066_, _05332_);
  and (_11068_, _11067_, _10998_);
  nor (_11069_, _11068_, _11065_);
  nor (_11070_, _11069_, _03243_);
  nor (_11071_, _11003_, _06122_);
  nor (_11072_, _11071_, _03244_);
  and (_11073_, _11072_, _11015_);
  nor (_11074_, _11073_, _11070_);
  nor (_11075_, _11074_, _03241_);
  and (_11076_, _11058_, _04835_);
  nor (_11077_, _11076_, _05357_);
  nand (_11078_, _11014_, _04835_);
  and (_11079_, _11078_, _03239_);
  or (_11080_, _11079_, _11077_);
  and (_11081_, _11080_, _10998_);
  or (_11082_, _11081_, _03123_);
  nor (_11083_, _11082_, _11075_);
  nor (_11084_, _11012_, _03124_);
  or (_11085_, _11084_, _02650_);
  nor (_11086_, _11085_, _11083_);
  nor (_11087_, _11035_, _03122_);
  or (_11088_, _11087_, _03121_);
  nor (_11089_, _11088_, _11086_);
  nor (_11090_, _11011_, _11003_);
  and (_11091_, _11090_, _03121_);
  nor (_11092_, _11091_, _11089_);
  or (_11093_, _11092_, _27789_);
  or (_11094_, _27788_, \oc8051_golden_model_1.IP [1]);
  and (_11095_, _11094_, _27053_);
  and (_28813_, _11095_, _11093_);
  not (_11096_, \oc8051_golden_model_1.IP [2]);
  nor (_11097_, _04581_, _11096_);
  and (_11098_, _04581_, _06009_);
  nor (_11099_, _11098_, _11097_);
  and (_11100_, _11099_, _02575_);
  nor (_11101_, _07034_, _03644_);
  nor (_11102_, _11101_, _11097_);
  and (_11103_, _11102_, _05949_);
  nor (_11104_, _08420_, _07034_);
  nor (_11105_, _11104_, _11097_);
  and (_11106_, _11105_, _02661_);
  and (_11107_, _04581_, \oc8051_golden_model_1.ACC [2]);
  nor (_11108_, _11107_, _11097_);
  nor (_11109_, _11108_, _05903_);
  nor (_11110_, _04505_, _11096_);
  or (_11111_, _11110_, _02661_);
  nor (_11112_, _11111_, _11109_);
  or (_11113_, _11112_, _06504_);
  nor (_11114_, _11113_, _11106_);
  nor (_11115_, _11102_, _03365_);
  nor (_11116_, _05425_, _11096_);
  and (_11117_, _08406_, _05425_);
  nor (_11118_, _11117_, _11116_);
  nor (_11119_, _11118_, _03390_);
  nor (_11120_, _11119_, _11115_);
  nand (_11121_, _11120_, _03179_);
  or (_11122_, _11121_, _11114_);
  nand (_11123_, _11108_, _03168_);
  and (_11124_, _11123_, _11122_);
  nor (_11125_, _11124_, _03176_);
  and (_11126_, _08404_, _05425_);
  nor (_11127_, _11126_, _11116_);
  and (_11128_, _11127_, _03176_);
  or (_11129_, _11128_, _03144_);
  nor (_11130_, _11129_, _11125_);
  nor (_11131_, _11116_, _08446_);
  or (_11132_, _11131_, _05168_);
  nor (_11133_, _11132_, _11118_);
  or (_11134_, _11133_, _11130_);
  and (_11135_, _11134_, _03141_);
  nor (_11136_, _08465_, _07071_);
  nor (_11137_, _11116_, _11136_);
  nor (_11138_, _11137_, _03141_);
  or (_11139_, _11138_, _05949_);
  nor (_11140_, _11139_, _11135_);
  nor (_11141_, _11140_, _11103_);
  nor (_11142_, _11141_, _05959_);
  and (_11143_, _04581_, _04170_);
  nor (_11144_, _11097_, _05963_);
  not (_11145_, _11144_);
  nor (_11146_, _11145_, _11143_);
  or (_11147_, _11146_, _02024_);
  nor (_11148_, _11147_, _11142_);
  nor (_11149_, _08522_, _07034_);
  nor (_11150_, _11149_, _11097_);
  nor (_11151_, _11150_, _03139_);
  or (_11152_, _11151_, _02575_);
  nor (_11153_, _11152_, _11148_);
  nor (_11154_, _11153_, _11100_);
  or (_11155_, _11154_, _02656_);
  and (_11156_, _08537_, _04581_);
  or (_11157_, _11156_, _11097_);
  or (_11158_, _11157_, _05305_);
  and (_11159_, _11158_, _03252_);
  and (_11160_, _11159_, _11155_);
  and (_11161_, _08387_, _04581_);
  nor (_11162_, _11161_, _11097_);
  nor (_11163_, _11162_, _03252_);
  nor (_11164_, _11163_, _11160_);
  nor (_11165_, _11164_, _02669_);
  nor (_11166_, _11097_, _06121_);
  not (_11167_, _11166_);
  nor (_11168_, _11099_, _05332_);
  and (_11169_, _11168_, _11167_);
  nor (_11170_, _11169_, _11165_);
  nor (_11171_, _11170_, _03243_);
  or (_11172_, _11166_, _03244_);
  nor (_11173_, _11172_, _11108_);
  or (_11174_, _11173_, _02654_);
  nor (_11175_, _11174_, _11171_);
  nor (_11176_, _08536_, _07034_);
  nor (_11177_, _11176_, _11097_);
  and (_11178_, _11177_, _02654_);
  nor (_11179_, _11178_, _11175_);
  and (_11180_, _11179_, _05883_);
  nor (_11181_, _08386_, _07034_);
  nor (_11182_, _11181_, _11097_);
  nor (_11183_, _11182_, _05883_);
  or (_11184_, _11183_, _11180_);
  and (_11185_, _11184_, _03124_);
  nor (_11186_, _11105_, _03124_);
  or (_11187_, _11186_, _02650_);
  or (_11188_, _11187_, _11185_);
  nand (_11189_, _11127_, _02650_);
  and (_11190_, _11189_, _11188_);
  nor (_11191_, _11190_, _03121_);
  and (_11192_, _08596_, _04581_);
  nor (_11193_, _11192_, _11097_);
  and (_11194_, _11193_, _03121_);
  nor (_11195_, _11194_, _11191_);
  or (_11196_, _11195_, _27789_);
  or (_11197_, _27788_, \oc8051_golden_model_1.IP [2]);
  and (_11198_, _11197_, _27053_);
  and (_28814_, _11198_, _11196_);
  not (_11199_, \oc8051_golden_model_1.IP [3]);
  nor (_11200_, _04581_, _11199_);
  and (_11201_, _04581_, _05986_);
  nor (_11202_, _11201_, _11200_);
  and (_11203_, _11202_, _02575_);
  nor (_11204_, _07034_, _03859_);
  nor (_11205_, _11204_, _11200_);
  and (_11206_, _11205_, _05949_);
  nor (_11207_, _08627_, _07071_);
  nor (_11208_, _05425_, _11199_);
  or (_11209_, _11208_, _03141_);
  or (_11210_, _11209_, _11207_);
  nor (_11211_, _08646_, _07034_);
  nor (_11212_, _11211_, _11200_);
  and (_11213_, _11212_, _02661_);
  and (_11214_, _04581_, \oc8051_golden_model_1.ACC [3]);
  nor (_11215_, _11214_, _11200_);
  nor (_11216_, _11215_, _05903_);
  nor (_11217_, _04505_, _11199_);
  or (_11218_, _11217_, _02661_);
  nor (_11219_, _11218_, _11216_);
  or (_11220_, _11219_, _06504_);
  nor (_11221_, _11220_, _11213_);
  nor (_11222_, _11205_, _03365_);
  and (_11223_, _08642_, _05425_);
  nor (_11224_, _11223_, _11208_);
  nor (_11225_, _11224_, _03390_);
  nor (_11226_, _11225_, _11222_);
  nand (_11227_, _11226_, _03179_);
  or (_11228_, _11227_, _11221_);
  nand (_11229_, _11215_, _03168_);
  and (_11230_, _11229_, _11228_);
  and (_11231_, _11230_, _03177_);
  and (_11232_, _08640_, _05425_);
  nor (_11233_, _11232_, _11208_);
  nor (_11234_, _11233_, _03177_);
  or (_11235_, _11234_, _11231_);
  and (_11236_, _11235_, _05168_);
  nor (_11237_, _11208_, _08671_);
  or (_11238_, _11224_, _05168_);
  nor (_11239_, _11238_, _11237_);
  or (_11240_, _11239_, _03140_);
  or (_11241_, _11240_, _11236_);
  and (_11242_, _11241_, _11210_);
  nor (_11243_, _11242_, _05949_);
  nor (_11244_, _11243_, _11206_);
  nor (_11245_, _11244_, _05959_);
  and (_11246_, _04581_, _04120_);
  nor (_11247_, _11200_, _05963_);
  not (_11248_, _11247_);
  nor (_11249_, _11248_, _11246_);
  or (_11250_, _11249_, _02024_);
  nor (_11251_, _11250_, _11245_);
  nor (_11252_, _08744_, _07034_);
  nor (_11253_, _11252_, _11200_);
  nor (_11254_, _11253_, _03139_);
  or (_11255_, _11254_, _02575_);
  nor (_11256_, _11255_, _11251_);
  nor (_11257_, _11256_, _11203_);
  or (_11258_, _11257_, _02656_);
  and (_11259_, _08622_, _04581_);
  or (_11260_, _11259_, _11200_);
  or (_11261_, _11260_, _05305_);
  and (_11262_, _11261_, _03252_);
  and (_11263_, _11262_, _11258_);
  and (_11264_, _08618_, _04581_);
  nor (_11265_, _11264_, _11200_);
  nor (_11266_, _11265_, _03252_);
  nor (_11267_, _11266_, _11263_);
  nor (_11268_, _11267_, _02669_);
  nor (_11269_, _11200_, _06120_);
  not (_11270_, _11269_);
  nor (_11271_, _11202_, _05332_);
  and (_11272_, _11271_, _11270_);
  nor (_11273_, _11272_, _11268_);
  nor (_11274_, _11273_, _03243_);
  or (_11275_, _11269_, _03244_);
  nor (_11276_, _11275_, _11215_);
  or (_11277_, _11276_, _02654_);
  nor (_11278_, _11277_, _11274_);
  nor (_11279_, _08621_, _07034_);
  nor (_11280_, _11279_, _11200_);
  and (_11281_, _11280_, _02654_);
  nor (_11282_, _11281_, _11278_);
  and (_11283_, _11282_, _05883_);
  nor (_11284_, _08617_, _07034_);
  nor (_11285_, _11284_, _11200_);
  nor (_11286_, _11285_, _05883_);
  or (_11287_, _11286_, _11283_);
  and (_11288_, _11287_, _03124_);
  nor (_11289_, _11212_, _03124_);
  or (_11290_, _11289_, _02650_);
  or (_11291_, _11290_, _11288_);
  nand (_11292_, _11233_, _02650_);
  and (_11293_, _11292_, _11291_);
  nor (_11294_, _11293_, _03121_);
  and (_11295_, _08807_, _04581_);
  nor (_11296_, _11295_, _11200_);
  and (_11297_, _11296_, _03121_);
  nor (_11298_, _11297_, _11294_);
  or (_11299_, _11298_, _27789_);
  or (_11300_, _27788_, \oc8051_golden_model_1.IP [3]);
  and (_11301_, _11300_, _27053_);
  and (_28815_, _11301_, _11299_);
  not (_11302_, \oc8051_golden_model_1.IP [4]);
  nor (_11303_, _04581_, _11302_);
  and (_11304_, _04581_, _05974_);
  nor (_11305_, _11304_, _11303_);
  and (_11306_, _11305_, _02575_);
  nor (_11307_, _07034_, _04325_);
  nor (_11308_, _11307_, _11303_);
  and (_11309_, _11308_, _05949_);
  nor (_11310_, _08838_, _07034_);
  nor (_11311_, _11310_, _11303_);
  and (_11312_, _11311_, _02661_);
  and (_11313_, _04581_, \oc8051_golden_model_1.ACC [4]);
  nor (_11314_, _11313_, _11303_);
  nor (_11315_, _11314_, _05903_);
  nor (_11316_, _04505_, _11302_);
  or (_11317_, _11316_, _02661_);
  nor (_11318_, _11317_, _11315_);
  or (_11319_, _11318_, _06504_);
  nor (_11320_, _11319_, _11312_);
  nor (_11321_, _11308_, _03365_);
  nor (_11322_, _05425_, _11302_);
  and (_11323_, _08869_, _05425_);
  nor (_11324_, _11323_, _11322_);
  nor (_11325_, _11324_, _03390_);
  nor (_11326_, _11325_, _11321_);
  nand (_11327_, _11326_, _03179_);
  or (_11328_, _11327_, _11320_);
  nand (_11329_, _11314_, _03168_);
  and (_11330_, _11329_, _11328_);
  and (_11331_, _11330_, _03177_);
  and (_11332_, _08880_, _05425_);
  nor (_11333_, _11332_, _11322_);
  nor (_11334_, _11333_, _03177_);
  or (_11335_, _11334_, _11331_);
  and (_11336_, _11335_, _05168_);
  and (_11337_, _08890_, _05425_);
  nor (_11338_, _11337_, _11322_);
  nor (_11339_, _11338_, _05168_);
  nor (_11340_, _11339_, _11336_);
  nor (_11341_, _11340_, _03140_);
  nor (_11342_, _08908_, _07071_);
  nor (_11343_, _11342_, _11322_);
  nor (_11344_, _11343_, _03141_);
  nor (_11345_, _11344_, _05949_);
  not (_11346_, _11345_);
  nor (_11347_, _11346_, _11341_);
  nor (_11348_, _11347_, _11309_);
  nor (_11349_, _11348_, _05959_);
  and (_11350_, _04581_, _04012_);
  nor (_11351_, _11303_, _05963_);
  not (_11352_, _11351_);
  nor (_11353_, _11352_, _11350_);
  or (_11354_, _11353_, _02024_);
  nor (_11355_, _11354_, _11349_);
  nor (_11356_, _08967_, _07034_);
  nor (_11357_, _11356_, _11303_);
  nor (_11358_, _11357_, _03139_);
  or (_11359_, _11358_, _02575_);
  nor (_11360_, _11359_, _11355_);
  nor (_11361_, _11360_, _11306_);
  or (_11362_, _11361_, _02656_);
  and (_11363_, _08982_, _04581_);
  or (_11364_, _11363_, _11303_);
  or (_11365_, _11364_, _05305_);
  and (_11366_, _11365_, _03252_);
  and (_11367_, _11366_, _11362_);
  and (_11368_, _08830_, _04581_);
  nor (_11369_, _11368_, _11303_);
  nor (_11370_, _11369_, _03252_);
  nor (_11371_, _11370_, _11367_);
  nor (_11372_, _11371_, _02669_);
  nor (_11373_, _11303_, _09034_);
  not (_11374_, _11373_);
  nor (_11375_, _11305_, _05332_);
  and (_11376_, _11375_, _11374_);
  nor (_11377_, _11376_, _11372_);
  nor (_11378_, _11377_, _03243_);
  or (_11379_, _11373_, _03244_);
  nor (_11380_, _11379_, _11314_);
  or (_11381_, _11380_, _02654_);
  nor (_11382_, _11381_, _11378_);
  nor (_11383_, _08981_, _07034_);
  nor (_11384_, _11383_, _11303_);
  and (_11385_, _11384_, _02654_);
  nor (_11386_, _11385_, _11382_);
  and (_11387_, _11386_, _05883_);
  nor (_11388_, _08828_, _07034_);
  nor (_11389_, _11388_, _11303_);
  nor (_11390_, _11389_, _05883_);
  or (_11391_, _11390_, _11387_);
  and (_11392_, _11391_, _03124_);
  nor (_11393_, _11311_, _03124_);
  or (_11394_, _11393_, _02650_);
  or (_11395_, _11394_, _11392_);
  nand (_11396_, _11333_, _02650_);
  and (_11397_, _11396_, _11395_);
  nor (_11398_, _11397_, _03121_);
  and (_11399_, _09037_, _04581_);
  nor (_11400_, _11399_, _11303_);
  and (_11401_, _11400_, _03121_);
  nor (_11402_, _11401_, _11398_);
  or (_11403_, _11402_, _27789_);
  or (_11404_, _27788_, \oc8051_golden_model_1.IP [4]);
  and (_11405_, _11404_, _27053_);
  and (_28816_, _11405_, _11403_);
  not (_11406_, \oc8051_golden_model_1.IP [5]);
  nor (_11407_, _04581_, _11406_);
  and (_11408_, _04581_, _06036_);
  nor (_11409_, _11408_, _11407_);
  and (_11410_, _11409_, _02575_);
  nor (_11411_, _07034_, _04480_);
  nor (_11412_, _11411_, _11407_);
  and (_11413_, _11412_, _05949_);
  nor (_11414_, _05425_, _11406_);
  nor (_11415_, _11414_, _09107_);
  and (_11416_, _09072_, _05425_);
  nor (_11417_, _11416_, _11414_);
  or (_11418_, _11417_, _05168_);
  nor (_11419_, _11418_, _11415_);
  nor (_11420_, _09087_, _07034_);
  nor (_11421_, _11420_, _11407_);
  and (_11422_, _11421_, _02661_);
  and (_11423_, _04581_, \oc8051_golden_model_1.ACC [5]);
  nor (_11424_, _11423_, _11407_);
  nor (_11425_, _11424_, _05903_);
  nor (_11426_, _04505_, _11406_);
  or (_11427_, _11426_, _02661_);
  nor (_11428_, _11427_, _11425_);
  or (_11429_, _11428_, _06504_);
  nor (_11430_, _11429_, _11422_);
  nor (_11431_, _11412_, _03365_);
  nor (_11432_, _11417_, _03390_);
  nor (_11433_, _11432_, _11431_);
  nand (_11434_, _11433_, _03179_);
  or (_11435_, _11434_, _11430_);
  nand (_11436_, _11424_, _03168_);
  and (_11437_, _11436_, _11435_);
  and (_11438_, _11437_, _03177_);
  and (_11439_, _09099_, _05425_);
  nor (_11440_, _11439_, _11414_);
  nor (_11441_, _11440_, _03177_);
  or (_11442_, _11441_, _11438_);
  and (_11443_, _11442_, _05168_);
  nor (_11444_, _11443_, _11419_);
  nor (_11445_, _11444_, _03140_);
  nor (_11446_, _09059_, _07071_);
  nor (_11447_, _11446_, _11414_);
  nor (_11448_, _11447_, _03141_);
  nor (_11449_, _11448_, _05949_);
  not (_11450_, _11449_);
  nor (_11451_, _11450_, _11445_);
  nor (_11452_, _11451_, _11413_);
  nor (_11453_, _11452_, _05959_);
  and (_11454_, _04581_, _03904_);
  nor (_11455_, _11407_, _05963_);
  not (_11456_, _11455_);
  nor (_11457_, _11456_, _11454_);
  or (_11458_, _11457_, _02024_);
  nor (_11459_, _11458_, _11453_);
  nor (_11460_, _09180_, _07034_);
  nor (_11461_, _11460_, _11407_);
  nor (_11462_, _11461_, _03139_);
  or (_11463_, _11462_, _02575_);
  nor (_11464_, _11463_, _11459_);
  nor (_11465_, _11464_, _11410_);
  or (_11466_, _11465_, _02656_);
  and (_11467_, _09195_, _04581_);
  or (_11468_, _11467_, _11407_);
  or (_11469_, _11468_, _05305_);
  and (_11470_, _11469_, _03252_);
  and (_11471_, _11470_, _11466_);
  and (_11472_, _09055_, _04581_);
  nor (_11473_, _11472_, _11407_);
  nor (_11474_, _11473_, _03252_);
  nor (_11475_, _11474_, _11471_);
  nor (_11476_, _11475_, _02669_);
  not (_11477_, _11407_);
  and (_11478_, _11477_, _04787_);
  not (_11479_, _11478_);
  nor (_11480_, _11409_, _05332_);
  and (_11481_, _11480_, _11479_);
  nor (_11482_, _11481_, _11476_);
  nor (_11483_, _11482_, _03243_);
  or (_11484_, _11478_, _03244_);
  nor (_11485_, _11484_, _11424_);
  or (_11486_, _11485_, _02654_);
  nor (_11487_, _11486_, _11483_);
  nor (_11488_, _09194_, _07034_);
  nor (_11489_, _11488_, _11407_);
  and (_11490_, _11489_, _02654_);
  nor (_11491_, _11490_, _11487_);
  and (_11492_, _11491_, _05883_);
  nor (_11493_, _09054_, _07034_);
  nor (_11494_, _11493_, _11407_);
  nor (_11495_, _11494_, _05883_);
  or (_11496_, _11495_, _11492_);
  and (_11497_, _11496_, _03124_);
  nor (_11498_, _11421_, _03124_);
  or (_11499_, _11498_, _02650_);
  or (_11500_, _11499_, _11497_);
  nand (_11501_, _11440_, _02650_);
  and (_11502_, _11501_, _11500_);
  nor (_11503_, _11502_, _03121_);
  and (_11504_, _09248_, _04581_);
  nor (_11505_, _11504_, _11407_);
  and (_11506_, _11505_, _03121_);
  nor (_11507_, _11506_, _11503_);
  or (_11508_, _11507_, _27789_);
  or (_11509_, _27788_, \oc8051_golden_model_1.IP [5]);
  and (_11510_, _11509_, _27053_);
  and (_28817_, _11510_, _11508_);
  not (_11511_, \oc8051_golden_model_1.IP [6]);
  nor (_11512_, _04581_, _11511_);
  and (_11513_, _04581_, _03960_);
  or (_11514_, _11513_, _11512_);
  and (_11515_, _11514_, _05959_);
  nor (_11516_, _05425_, _11511_);
  not (_11517_, _11516_);
  and (_11518_, _11517_, _09320_);
  and (_11519_, _09305_, _05425_);
  nor (_11520_, _11519_, _11516_);
  or (_11521_, _11520_, _05168_);
  nor (_11522_, _11521_, _11518_);
  nor (_11523_, _09301_, _07034_);
  nor (_11524_, _11523_, _11512_);
  and (_11525_, _11524_, _02661_);
  and (_11526_, _04581_, \oc8051_golden_model_1.ACC [6]);
  nor (_11527_, _11526_, _11512_);
  nor (_11528_, _11527_, _05903_);
  nor (_11529_, _04505_, _11511_);
  or (_11530_, _11529_, _02661_);
  nor (_11531_, _11530_, _11528_);
  or (_11532_, _11531_, _06504_);
  nor (_11533_, _11532_, _11525_);
  nor (_11534_, _07034_, _04373_);
  nor (_11535_, _11534_, _11512_);
  nor (_11536_, _11535_, _03365_);
  nor (_11537_, _11520_, _03390_);
  nor (_11538_, _11537_, _11536_);
  nand (_11539_, _11538_, _03179_);
  or (_11540_, _11539_, _11533_);
  nand (_11541_, _11527_, _03168_);
  and (_11542_, _11541_, _11540_);
  and (_11543_, _11542_, _03177_);
  and (_11544_, _09286_, _05425_);
  nor (_11545_, _11544_, _11516_);
  nor (_11546_, _11545_, _03177_);
  or (_11547_, _11546_, _11543_);
  and (_11548_, _11547_, _05168_);
  nor (_11549_, _11548_, _11522_);
  nor (_11550_, _11549_, _03140_);
  nor (_11551_, _09272_, _07071_);
  nor (_11552_, _11551_, _11516_);
  nor (_11553_, _11552_, _03141_);
  nor (_11554_, _11553_, _05949_);
  not (_11555_, _11554_);
  nor (_11556_, _11555_, _11550_);
  and (_11557_, _11535_, _05949_);
  or (_11558_, _11557_, _05959_);
  nor (_11559_, _11558_, _11556_);
  or (_11560_, _11559_, _11515_);
  and (_11561_, _11560_, _03139_);
  and (_11562_, _09388_, _04581_);
  nor (_11563_, _11562_, _11512_);
  nor (_11564_, _11563_, _03139_);
  or (_11565_, _11564_, _06549_);
  or (_11566_, _11565_, _11561_);
  and (_11567_, _09404_, _04581_);
  or (_11568_, _11512_, _05305_);
  or (_11569_, _11568_, _11567_);
  and (_11570_, _04581_, _09395_);
  nor (_11571_, _11570_, _11512_);
  and (_11572_, _11571_, _02575_);
  nor (_11573_, _11572_, _03251_);
  and (_11574_, _11573_, _11569_);
  and (_11575_, _11574_, _11566_);
  and (_11576_, _09268_, _04581_);
  nor (_11577_, _11576_, _11512_);
  nor (_11578_, _11577_, _03252_);
  nor (_11579_, _11578_, _11575_);
  nor (_11580_, _11579_, _02669_);
  nor (_11581_, _11512_, _06119_);
  not (_11582_, _11581_);
  nor (_11583_, _11571_, _05332_);
  and (_11584_, _11583_, _11582_);
  nor (_11585_, _11584_, _11580_);
  nor (_11586_, _11585_, _03243_);
  or (_11587_, _11581_, _03244_);
  nor (_11588_, _11587_, _11527_);
  or (_11589_, _11588_, _02654_);
  nor (_11590_, _11589_, _11586_);
  nor (_11591_, _09403_, _07034_);
  nor (_11592_, _11591_, _11512_);
  and (_11593_, _11592_, _02654_);
  nor (_11594_, _11593_, _11590_);
  and (_11595_, _11594_, _05883_);
  nor (_11596_, _09267_, _07034_);
  nor (_11597_, _11596_, _11512_);
  nor (_11598_, _11597_, _05883_);
  or (_11599_, _11598_, _11595_);
  and (_11600_, _11599_, _03124_);
  nor (_11601_, _11524_, _03124_);
  or (_11602_, _11601_, _02650_);
  or (_11603_, _11602_, _11600_);
  nand (_11604_, _11545_, _02650_);
  and (_11605_, _11604_, _11603_);
  nor (_11606_, _11605_, _03121_);
  and (_11607_, _09456_, _04581_);
  nor (_11608_, _11607_, _11512_);
  and (_11609_, _11608_, _03121_);
  nor (_11610_, _11609_, _11606_);
  or (_11611_, _11610_, _27789_);
  or (_11612_, _27788_, \oc8051_golden_model_1.IP [6]);
  and (_11613_, _11612_, _27053_);
  and (_28818_, _11613_, _11611_);
  not (_11614_, \oc8051_golden_model_1.P0 [0]);
  nor (_11615_, _27788_, _11614_);
  or (_28821_, _11615_, rst);
  nor (_11616_, \oc8051_golden_model_1.P0 [1], rst);
  nor (_28822_, _11616_, _00001_);
  not (_11617_, \oc8051_golden_model_1.P0 [2]);
  nor (_11618_, _27788_, _11617_);
  or (_28823_, _11618_, rst);
  nor (_11619_, \oc8051_golden_model_1.P0 [3], rst);
  nor (_28824_, _11619_, _00001_);
  not (_11620_, \oc8051_golden_model_1.P0 [4]);
  nor (_11621_, _27788_, _11620_);
  or (_28825_, _11621_, rst);
  nor (_11622_, \oc8051_golden_model_1.P0 [5], rst);
  nor (_28826_, _11622_, _00001_);
  not (_11623_, \oc8051_golden_model_1.P0 [6]);
  nor (_11624_, _27788_, _11623_);
  or (_28827_, _11624_, rst);
  not (_11625_, \oc8051_golden_model_1.P1 [0]);
  nor (_11626_, _27788_, _11625_);
  or (_28830_, _11626_, rst);
  nor (_11627_, \oc8051_golden_model_1.P1 [1], rst);
  nor (_28831_, _11627_, _00001_);
  not (_11628_, \oc8051_golden_model_1.P1 [2]);
  nor (_11629_, _27788_, _11628_);
  or (_28832_, _11629_, rst);
  nor (_11630_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_28833_, _11630_, _00001_);
  not (_11631_, \oc8051_golden_model_1.P1 [4]);
  nor (_11632_, _27788_, _11631_);
  or (_28834_, _11632_, rst);
  nor (_11633_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_28835_, _11633_, _00001_);
  not (_11634_, \oc8051_golden_model_1.P1 [6]);
  nor (_11635_, _27788_, _11634_);
  or (_28836_, _11635_, rst);
  not (_11636_, \oc8051_golden_model_1.P2 [0]);
  nor (_11637_, _27788_, _11636_);
  or (_28841_, _11637_, rst);
  nor (_11638_, \oc8051_golden_model_1.P2 [1], rst);
  nor (_28842_, _11638_, _00001_);
  not (_11639_, \oc8051_golden_model_1.P2 [2]);
  nor (_11640_, _27788_, _11639_);
  or (_28843_, _11640_, rst);
  nor (_11641_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_28844_, _11641_, _00001_);
  not (_11642_, \oc8051_golden_model_1.P2 [4]);
  nor (_11643_, _27788_, _11642_);
  or (_28845_, _11643_, rst);
  nor (_11644_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_28846_, _11644_, _00001_);
  not (_11645_, \oc8051_golden_model_1.P2 [6]);
  nor (_11646_, _27788_, _11645_);
  or (_28847_, _11646_, rst);
  not (_11647_, \oc8051_golden_model_1.P3 [0]);
  nor (_11648_, _27788_, _11647_);
  or (_28850_, _11648_, rst);
  nor (_11649_, \oc8051_golden_model_1.P3 [1], rst);
  nor (_28851_, _11649_, _00001_);
  not (_11650_, \oc8051_golden_model_1.P3 [2]);
  nor (_11651_, _27788_, _11650_);
  or (_28852_, _11651_, rst);
  nor (_11652_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_28853_, _11652_, _00001_);
  not (_11653_, \oc8051_golden_model_1.P3 [4]);
  nor (_11654_, _27788_, _11653_);
  or (_28854_, _11654_, rst);
  nor (_11655_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_28855_, _11655_, _00001_);
  not (_11656_, \oc8051_golden_model_1.P3 [6]);
  nor (_11657_, _27788_, _11656_);
  or (_28856_, _11657_, rst);
  nand (_11658_, \oc8051_golden_model_1.PSW [0], _27053_);
  nor (_28859_, _11658_, _27788_);
  not (_11659_, \oc8051_golden_model_1.PSW [1]);
  or (_11660_, _11659_, rst);
  nor (_28860_, _11660_, _27788_);
  nand (_11661_, \oc8051_golden_model_1.PSW [2], _27053_);
  nor (_28861_, _11661_, _27788_);
  or (_11662_, _03159_, rst);
  nor (_28862_, _11662_, _27788_);
  not (_11663_, \oc8051_golden_model_1.PSW [4]);
  or (_11664_, _11663_, rst);
  nor (_28863_, _11664_, _27788_);
  not (_11665_, \oc8051_golden_model_1.PSW [5]);
  or (_11666_, _11665_, rst);
  nor (_28864_, _11666_, _27788_);
  nand (_11667_, \oc8051_golden_model_1.PSW [6], _27053_);
  nor (_28867_, _11667_, _27788_);
  not (_11668_, \oc8051_golden_model_1.PCON [0]);
  nor (_11669_, _04623_, _11668_);
  nor (_11670_, _04888_, _06956_);
  nor (_11671_, _11670_, _11669_);
  and (_11672_, _07527_, _02023_);
  and (_11673_, _11672_, _11671_);
  and (_11674_, _04623_, _05996_);
  nor (_11675_, _11674_, _11669_);
  nor (_11676_, _11675_, _05332_);
  not (_11677_, _11676_);
  nor (_11678_, _11677_, _11670_);
  nor (_11679_, _06956_, _04485_);
  nor (_11680_, _11679_, _11669_);
  and (_11681_, _11680_, _05949_);
  and (_11682_, _04623_, \oc8051_golden_model_1.ACC [0]);
  nor (_11683_, _11682_, _11669_);
  nor (_11684_, _11683_, _05903_);
  nor (_11685_, _04505_, _11668_);
  or (_11686_, _11685_, _11684_);
  and (_11687_, _11686_, _02662_);
  nor (_11688_, _11671_, _02662_);
  or (_11689_, _11688_, _11687_);
  and (_11690_, _11689_, _03365_);
  nor (_11691_, _11680_, _03365_);
  nor (_11692_, _11691_, _11690_);
  nor (_11693_, _11692_, _03168_);
  nor (_11694_, _11683_, _03179_);
  nor (_11695_, _11694_, _05949_);
  not (_11696_, _11695_);
  nor (_11697_, _11696_, _11693_);
  nor (_11698_, _11697_, _11681_);
  nor (_11699_, _11698_, _05959_);
  and (_11700_, _04623_, _04268_);
  nor (_11701_, _11669_, _05963_);
  not (_11702_, _11701_);
  nor (_11703_, _11702_, _11700_);
  nor (_11704_, _11703_, _11699_);
  nor (_11705_, _11704_, _02024_);
  nor (_11706_, _08093_, _06956_);
  or (_11707_, _11669_, _03139_);
  nor (_11708_, _11707_, _11706_);
  or (_11709_, _11708_, _02575_);
  nor (_11710_, _11709_, _11705_);
  nand (_11711_, _11675_, _05305_);
  and (_11712_, _11711_, _06549_);
  nor (_11713_, _11712_, _11710_);
  and (_11714_, _07968_, _04623_);
  nor (_11715_, _11714_, _11669_);
  and (_11716_, _11715_, _02656_);
  nor (_11717_, _11716_, _11713_);
  and (_11718_, _11717_, _03252_);
  and (_11719_, _08110_, _04623_);
  nor (_11720_, _11719_, _11669_);
  nor (_11721_, _11720_, _03252_);
  or (_11722_, _11721_, _11718_);
  and (_11723_, _11722_, _05332_);
  nor (_11724_, _11723_, _11678_);
  nor (_11725_, _11724_, _03243_);
  and (_11726_, _08108_, _04623_);
  or (_11727_, _11726_, _11669_);
  and (_11728_, _11727_, _03243_);
  or (_11729_, _11728_, _11725_);
  and (_11730_, _11729_, _05357_);
  nor (_11731_, _07967_, _06956_);
  nor (_11732_, _11731_, _11669_);
  nor (_11733_, _11732_, _05357_);
  or (_11734_, _11733_, _11730_);
  and (_11735_, _11734_, _05883_);
  nor (_11736_, _08109_, _06956_);
  nor (_11737_, _11736_, _11669_);
  nor (_11738_, _11737_, _05883_);
  nor (_11739_, _11738_, _11672_);
  not (_11740_, _11739_);
  nor (_11741_, _11740_, _11735_);
  nor (_11742_, _11741_, _11673_);
  or (_11743_, _11742_, _27789_);
  or (_11744_, _27788_, \oc8051_golden_model_1.PCON [0]);
  and (_11745_, _11744_, _27053_);
  and (_28868_, _11745_, _11743_);
  nor (_11746_, _04623_, \oc8051_golden_model_1.PCON [1]);
  and (_11747_, _08209_, _04623_);
  nor (_11748_, _11747_, _11746_);
  nor (_11749_, _11748_, _03124_);
  not (_11750_, _11746_);
  nor (_11751_, _08184_, _06956_);
  nor (_11752_, _11751_, _05332_);
  and (_11753_, _11752_, _11750_);
  nor (_11754_, _08325_, _06956_);
  nor (_11755_, _11754_, _03252_);
  and (_11756_, _11755_, _11750_);
  and (_11757_, _04623_, _04218_);
  not (_11758_, \oc8051_golden_model_1.PCON [1]);
  nor (_11759_, _04623_, _11758_);
  nor (_11760_, _11759_, _05963_);
  not (_11761_, _11760_);
  nor (_11762_, _11761_, _11757_);
  not (_11763_, _11762_);
  and (_11764_, _04623_, _08322_);
  nor (_11765_, _11764_, _11746_);
  and (_11766_, _11765_, _03168_);
  and (_11767_, _11765_, _04505_);
  nor (_11768_, _04505_, _11758_);
  or (_11769_, _11768_, _11767_);
  and (_11770_, _11769_, _02662_);
  and (_11771_, _11748_, _02661_);
  or (_11772_, _11771_, _11770_);
  and (_11773_, _11772_, _03365_);
  nor (_11774_, _06956_, _03777_);
  nor (_11775_, _11774_, _11759_);
  nor (_11776_, _11775_, _03365_);
  nor (_11777_, _11776_, _11773_);
  nor (_11778_, _11777_, _03168_);
  or (_11779_, _11778_, _05949_);
  nor (_11780_, _11779_, _11766_);
  and (_11781_, _11775_, _05949_);
  nor (_11782_, _11781_, _11780_);
  nor (_11783_, _11782_, _05959_);
  nor (_11784_, _11783_, _02024_);
  and (_11785_, _11784_, _11763_);
  and (_11786_, _08307_, _04623_);
  nor (_11787_, _11786_, _03139_);
  and (_11788_, _11787_, _11750_);
  nor (_11789_, _11788_, _11785_);
  nor (_11790_, _11789_, _06549_);
  nor (_11791_, _08185_, _06956_);
  nor (_11792_, _11791_, _05305_);
  and (_11793_, _04623_, _03016_);
  nor (_11794_, _11793_, _05245_);
  or (_11795_, _11794_, _11792_);
  and (_11796_, _11795_, _11750_);
  nor (_11797_, _11796_, _11790_);
  nor (_11798_, _11797_, _03251_);
  nor (_11799_, _11798_, _11756_);
  nor (_11800_, _11799_, _02669_);
  nor (_11801_, _11800_, _11753_);
  nor (_11802_, _11801_, _03243_);
  nor (_11803_, _11759_, _06122_);
  nor (_11804_, _11803_, _03244_);
  and (_11805_, _11804_, _11765_);
  nor (_11806_, _11805_, _11802_);
  nor (_11807_, _11806_, _03241_);
  and (_11808_, _11793_, _04835_);
  nor (_11809_, _11808_, _05357_);
  nand (_11810_, _11764_, _04835_);
  and (_11811_, _11810_, _03239_);
  or (_11812_, _11811_, _11809_);
  and (_11813_, _11812_, _11750_);
  or (_11814_, _11813_, _03123_);
  nor (_11815_, _11814_, _11807_);
  nor (_11816_, _11815_, _11749_);
  nor (_11817_, _11816_, _03121_);
  nor (_11818_, _11759_, _11747_);
  and (_11819_, _11818_, _03121_);
  nor (_11820_, _11819_, _11817_);
  or (_11821_, _11820_, _27789_);
  or (_11822_, _27788_, \oc8051_golden_model_1.PCON [1]);
  and (_11823_, _11822_, _27053_);
  and (_28869_, _11823_, _11821_);
  not (_11824_, \oc8051_golden_model_1.PCON [2]);
  nor (_11825_, _04623_, _11824_);
  nor (_11826_, _11825_, _06121_);
  not (_11827_, _11826_);
  and (_11828_, _04623_, _06009_);
  nor (_11829_, _11828_, _11825_);
  nor (_11830_, _11829_, _05332_);
  and (_11831_, _11830_, _11827_);
  and (_11832_, _04623_, _04170_);
  nor (_11833_, _11832_, _11825_);
  or (_11834_, _11833_, _05963_);
  and (_11835_, _04623_, \oc8051_golden_model_1.ACC [2]);
  nor (_11836_, _11835_, _11825_);
  nor (_11837_, _11836_, _05903_);
  nor (_11838_, _04505_, _11824_);
  or (_11839_, _11838_, _11837_);
  and (_11840_, _11839_, _02662_);
  nor (_11841_, _08420_, _06956_);
  nor (_11842_, _11841_, _11825_);
  nor (_11843_, _11842_, _02662_);
  or (_11844_, _11843_, _11840_);
  and (_11845_, _11844_, _03365_);
  nor (_11846_, _06956_, _03644_);
  nor (_11847_, _11846_, _11825_);
  nor (_11848_, _11847_, _03365_);
  nor (_11849_, _11848_, _11845_);
  nor (_11850_, _11849_, _03168_);
  nor (_11851_, _11836_, _03179_);
  nor (_11852_, _11851_, _05949_);
  not (_11853_, _11852_);
  nor (_11854_, _11853_, _11850_);
  and (_11855_, _11847_, _05949_);
  or (_11856_, _11855_, _05959_);
  or (_11857_, _11856_, _11854_);
  and (_11858_, _11857_, _03139_);
  and (_11859_, _11858_, _11834_);
  nor (_11860_, _08522_, _06956_);
  or (_11861_, _11825_, _03139_);
  nor (_11862_, _11861_, _11860_);
  or (_11863_, _11862_, _02575_);
  nor (_11864_, _11863_, _11859_);
  nand (_11865_, _11829_, _05305_);
  and (_11866_, _11865_, _06549_);
  nor (_11867_, _11866_, _11864_);
  and (_11868_, _08537_, _04623_);
  nor (_11869_, _11868_, _11825_);
  and (_11870_, _11869_, _02656_);
  nor (_11871_, _11870_, _11867_);
  and (_11872_, _11871_, _03252_);
  and (_11873_, _08387_, _04623_);
  nor (_11874_, _11873_, _11825_);
  nor (_11875_, _11874_, _03252_);
  or (_11876_, _11875_, _11872_);
  and (_11877_, _11876_, _05332_);
  nor (_11878_, _11877_, _11831_);
  nor (_11879_, _11878_, _03243_);
  or (_11880_, _11826_, _03244_);
  nor (_11881_, _11880_, _11836_);
  or (_11882_, _11881_, _02654_);
  nor (_11883_, _11882_, _11879_);
  nor (_11884_, _08536_, _06956_);
  nor (_11885_, _11884_, _11825_);
  and (_11886_, _11885_, _02654_);
  nor (_11887_, _11886_, _11883_);
  and (_11888_, _11887_, _05883_);
  nor (_11889_, _08386_, _06956_);
  nor (_11890_, _11889_, _11825_);
  nor (_11891_, _11890_, _05883_);
  or (_11892_, _11891_, _11888_);
  and (_11893_, _11892_, _03124_);
  nor (_11894_, _11842_, _03124_);
  or (_11895_, _11894_, _11893_);
  and (_11896_, _11895_, _03513_);
  and (_11897_, _08596_, _04623_);
  nor (_11898_, _11897_, _11825_);
  nor (_11899_, _11898_, _03513_);
  or (_11900_, _11899_, _11896_);
  or (_11901_, _11900_, _27789_);
  or (_11902_, _27788_, \oc8051_golden_model_1.PCON [2]);
  and (_11903_, _11902_, _27053_);
  and (_28872_, _11903_, _11901_);
  not (_11904_, \oc8051_golden_model_1.PCON [3]);
  nor (_11905_, _04623_, _11904_);
  nor (_11906_, _11905_, _06120_);
  not (_11907_, _11906_);
  and (_11908_, _04623_, _05986_);
  nor (_11909_, _11908_, _11905_);
  nor (_11910_, _11909_, _05332_);
  and (_11911_, _11910_, _11907_);
  and (_11912_, _04623_, \oc8051_golden_model_1.ACC [3]);
  nor (_11913_, _11912_, _11905_);
  nor (_11914_, _11913_, _05903_);
  nor (_11915_, _04505_, _11904_);
  or (_11916_, _11915_, _11914_);
  and (_11917_, _11916_, _02662_);
  nor (_11918_, _08646_, _06956_);
  nor (_11919_, _11918_, _11905_);
  nor (_11920_, _11919_, _02662_);
  or (_11921_, _11920_, _11917_);
  and (_11922_, _11921_, _03365_);
  nor (_11923_, _06956_, _03859_);
  nor (_11924_, _11923_, _11905_);
  nor (_11925_, _11924_, _03365_);
  nor (_11926_, _11925_, _11922_);
  nor (_11927_, _11926_, _03168_);
  nor (_11928_, _11913_, _03179_);
  nor (_11929_, _11928_, _05949_);
  not (_11930_, _11929_);
  nor (_11931_, _11930_, _11927_);
  and (_11932_, _11924_, _05949_);
  or (_11933_, _11932_, _05959_);
  or (_11934_, _11933_, _11931_);
  and (_11935_, _04623_, _04120_);
  nor (_11936_, _11935_, _11905_);
  or (_11937_, _11936_, _05963_);
  and (_11938_, _11937_, _03139_);
  and (_11939_, _11938_, _11934_);
  nor (_11940_, _08744_, _06956_);
  or (_11941_, _11905_, _03139_);
  nor (_11942_, _11941_, _11940_);
  or (_11943_, _11942_, _02575_);
  nor (_11944_, _11943_, _11939_);
  nand (_11945_, _11909_, _05305_);
  and (_11946_, _11945_, _06549_);
  nor (_11947_, _11946_, _11944_);
  and (_11948_, _08622_, _04623_);
  nor (_11949_, _11948_, _11905_);
  and (_11950_, _11949_, _02656_);
  nor (_11951_, _11950_, _11947_);
  and (_11952_, _11951_, _03252_);
  and (_11953_, _08618_, _04623_);
  nor (_11954_, _11953_, _11905_);
  nor (_11955_, _11954_, _03252_);
  or (_11956_, _11955_, _11952_);
  and (_11957_, _11956_, _05332_);
  nor (_11958_, _11957_, _11911_);
  nor (_11959_, _11958_, _03243_);
  or (_11960_, _11906_, _03244_);
  nor (_11961_, _11960_, _11913_);
  or (_11962_, _11961_, _02654_);
  nor (_11963_, _11962_, _11959_);
  nor (_11964_, _08621_, _06956_);
  nor (_11965_, _11964_, _11905_);
  and (_11966_, _11965_, _02654_);
  nor (_11967_, _11966_, _11963_);
  and (_11968_, _11967_, _05883_);
  nor (_11969_, _08617_, _06956_);
  nor (_11970_, _11969_, _11905_);
  nor (_11971_, _11970_, _05883_);
  or (_11972_, _11971_, _11968_);
  and (_11973_, _11972_, _03124_);
  nor (_11974_, _11919_, _03124_);
  or (_11975_, _11974_, _11973_);
  and (_11976_, _11975_, _03513_);
  and (_11977_, _08807_, _04623_);
  nor (_11978_, _11977_, _11905_);
  nor (_11979_, _11978_, _03513_);
  or (_11980_, _11979_, _11976_);
  or (_11981_, _11980_, _27789_);
  or (_11982_, _27788_, \oc8051_golden_model_1.PCON [3]);
  and (_11983_, _11982_, _27053_);
  and (_28873_, _11983_, _11981_);
  not (_11984_, \oc8051_golden_model_1.PCON [4]);
  nor (_11985_, _04623_, _11984_);
  and (_11986_, _08830_, _04623_);
  nor (_11987_, _11986_, _11985_);
  nor (_11988_, _11987_, _03252_);
  and (_11989_, _04623_, _05974_);
  nor (_11990_, _11989_, _11985_);
  and (_11991_, _11990_, _02575_);
  and (_11992_, _04623_, \oc8051_golden_model_1.ACC [4]);
  nor (_11993_, _11992_, _11985_);
  nor (_11994_, _11993_, _03179_);
  nor (_11995_, _11993_, _05903_);
  nor (_11996_, _04505_, _11984_);
  or (_11997_, _11996_, _11995_);
  and (_11998_, _11997_, _02662_);
  nor (_11999_, _08838_, _06956_);
  nor (_12000_, _11999_, _11985_);
  nor (_12001_, _12000_, _02662_);
  or (_12002_, _12001_, _11998_);
  and (_12003_, _12002_, _03365_);
  nor (_12004_, _06956_, _04325_);
  nor (_12005_, _12004_, _11985_);
  nor (_12006_, _12005_, _03365_);
  nor (_12007_, _12006_, _12003_);
  nor (_12008_, _12007_, _03168_);
  or (_12009_, _12008_, _05949_);
  nor (_12010_, _12009_, _11994_);
  and (_12011_, _12005_, _05949_);
  nor (_12012_, _12011_, _12010_);
  nor (_12013_, _12012_, _05959_);
  and (_12014_, _04623_, _04012_);
  nor (_12015_, _11985_, _05963_);
  not (_12016_, _12015_);
  nor (_12017_, _12016_, _12014_);
  or (_12018_, _12017_, _02024_);
  nor (_12019_, _12018_, _12013_);
  nor (_12020_, _08967_, _06956_);
  nor (_12021_, _12020_, _11985_);
  nor (_12022_, _12021_, _03139_);
  or (_12023_, _12022_, _02575_);
  nor (_12024_, _12023_, _12019_);
  nor (_12025_, _12024_, _11991_);
  or (_12026_, _12025_, _02656_);
  and (_12027_, _08982_, _04623_);
  or (_12028_, _12027_, _11985_);
  or (_12029_, _12028_, _05305_);
  and (_12030_, _12029_, _03252_);
  and (_12031_, _12030_, _12026_);
  nor (_12032_, _12031_, _11988_);
  nor (_12033_, _12032_, _02669_);
  nor (_12034_, _11985_, _09034_);
  not (_12035_, _12034_);
  nor (_12036_, _11990_, _05332_);
  and (_12037_, _12036_, _12035_);
  nor (_12038_, _12037_, _12033_);
  nor (_12039_, _12038_, _03243_);
  or (_12040_, _12034_, _03244_);
  nor (_12041_, _12040_, _11993_);
  or (_12042_, _12041_, _02654_);
  nor (_12043_, _12042_, _12039_);
  nor (_12044_, _08981_, _06956_);
  nor (_12045_, _12044_, _11985_);
  and (_12046_, _12045_, _02654_);
  nor (_12047_, _12046_, _12043_);
  and (_12048_, _12047_, _05883_);
  nor (_12049_, _08828_, _06956_);
  nor (_12050_, _12049_, _11985_);
  nor (_12051_, _12050_, _05883_);
  or (_12052_, _12051_, _12048_);
  and (_12053_, _12052_, _03124_);
  nor (_12054_, _12000_, _03124_);
  nor (_12055_, _12054_, _03121_);
  not (_12056_, _12055_);
  nor (_12057_, _12056_, _12053_);
  and (_12058_, _09037_, _04623_);
  nor (_12059_, _12058_, _11985_);
  and (_12060_, _12059_, _03121_);
  nor (_12061_, _12060_, _12057_);
  or (_12062_, _12061_, _27789_);
  or (_12063_, _27788_, \oc8051_golden_model_1.PCON [4]);
  and (_12064_, _12063_, _27053_);
  and (_28874_, _12064_, _12062_);
  not (_12065_, \oc8051_golden_model_1.PCON [5]);
  nor (_12066_, _04623_, _12065_);
  and (_12067_, _09055_, _04623_);
  nor (_12068_, _12067_, _12066_);
  nor (_12069_, _12068_, _03252_);
  and (_12070_, _04623_, _06036_);
  nor (_12071_, _12070_, _12066_);
  and (_12072_, _12071_, _02575_);
  nor (_12073_, _06956_, _04480_);
  nor (_12074_, _12073_, _12066_);
  and (_12075_, _12074_, _05949_);
  and (_12076_, _04623_, \oc8051_golden_model_1.ACC [5]);
  nor (_12077_, _12076_, _12066_);
  nor (_12078_, _12077_, _05903_);
  nor (_12079_, _04505_, _12065_);
  or (_12080_, _12079_, _12078_);
  and (_12081_, _12080_, _02662_);
  nor (_12082_, _09087_, _06956_);
  nor (_12083_, _12082_, _12066_);
  nor (_12084_, _12083_, _02662_);
  or (_12085_, _12084_, _12081_);
  and (_12086_, _12085_, _03365_);
  nor (_12087_, _12074_, _03365_);
  nor (_12088_, _12087_, _12086_);
  nor (_12089_, _12088_, _03168_);
  nor (_12090_, _12077_, _03179_);
  nor (_12091_, _12090_, _05949_);
  not (_12092_, _12091_);
  nor (_12093_, _12092_, _12089_);
  nor (_12094_, _12093_, _12075_);
  nor (_12095_, _12094_, _05959_);
  and (_12096_, _04623_, _03904_);
  nor (_12097_, _12066_, _05963_);
  not (_12098_, _12097_);
  nor (_12099_, _12098_, _12096_);
  or (_12100_, _12099_, _02024_);
  nor (_12101_, _12100_, _12095_);
  nor (_12102_, _09180_, _06956_);
  nor (_12103_, _12102_, _12066_);
  nor (_12104_, _12103_, _03139_);
  or (_12106_, _12104_, _02575_);
  nor (_12107_, _12106_, _12101_);
  nor (_12109_, _12107_, _12072_);
  or (_12110_, _12109_, _02656_);
  and (_12112_, _09195_, _04623_);
  or (_12113_, _12112_, _12066_);
  or (_12115_, _12113_, _05305_);
  and (_12116_, _12115_, _03252_);
  and (_12118_, _12116_, _12110_);
  nor (_12119_, _12118_, _12069_);
  nor (_12121_, _12119_, _02669_);
  not (_12122_, _12066_);
  and (_12124_, _12122_, _04787_);
  not (_12125_, _12124_);
  nor (_12127_, _12071_, _05332_);
  and (_12128_, _12127_, _12125_);
  nor (_12130_, _12128_, _12121_);
  nor (_12131_, _12130_, _03243_);
  or (_12133_, _12124_, _03244_);
  nor (_12134_, _12133_, _12077_);
  or (_12136_, _12134_, _02654_);
  nor (_12137_, _12136_, _12131_);
  nor (_12139_, _09194_, _06956_);
  nor (_12140_, _12139_, _12066_);
  and (_12142_, _12140_, _02654_);
  nor (_12143_, _12142_, _12137_);
  and (_12144_, _12143_, _05883_);
  nor (_12145_, _09054_, _06956_);
  nor (_12146_, _12145_, _12066_);
  nor (_12147_, _12146_, _05883_);
  or (_12148_, _12147_, _12144_);
  and (_12149_, _12148_, _03124_);
  nor (_12150_, _12083_, _03124_);
  or (_12151_, _12150_, _12149_);
  and (_12152_, _12151_, _03513_);
  and (_12153_, _09248_, _04623_);
  nor (_12154_, _12153_, _12066_);
  nor (_12155_, _12154_, _03513_);
  or (_12156_, _12155_, _12152_);
  or (_12157_, _12156_, _27789_);
  or (_12158_, _27788_, \oc8051_golden_model_1.PCON [5]);
  and (_12159_, _12158_, _27053_);
  and (_28875_, _12159_, _12157_);
  not (_12160_, \oc8051_golden_model_1.PCON [6]);
  nor (_12161_, _04623_, _12160_);
  and (_12162_, _09268_, _04623_);
  nor (_12163_, _12162_, _12161_);
  nor (_12164_, _12163_, _03252_);
  and (_12165_, _04623_, _03960_);
  or (_12166_, _12165_, _12161_);
  and (_12167_, _12166_, _05959_);
  and (_12168_, _04623_, \oc8051_golden_model_1.ACC [6]);
  nor (_12169_, _12168_, _12161_);
  nor (_12170_, _12169_, _05903_);
  nor (_12171_, _04505_, _12160_);
  or (_12172_, _12171_, _12170_);
  and (_12173_, _12172_, _02662_);
  nor (_12174_, _09301_, _06956_);
  nor (_12175_, _12174_, _12161_);
  nor (_12176_, _12175_, _02662_);
  or (_12177_, _12176_, _12173_);
  and (_12178_, _12177_, _03365_);
  nor (_12179_, _06956_, _04373_);
  nor (_12180_, _12179_, _12161_);
  nor (_12181_, _12180_, _03365_);
  nor (_12182_, _12181_, _12178_);
  nor (_12183_, _12182_, _03168_);
  nor (_12184_, _12169_, _03179_);
  nor (_12185_, _12184_, _05949_);
  not (_12186_, _12185_);
  nor (_12187_, _12186_, _12183_);
  and (_12188_, _12180_, _05949_);
  or (_12190_, _12188_, _05959_);
  nor (_12192_, _12190_, _12187_);
  or (_12193_, _12192_, _12167_);
  and (_12195_, _12193_, _03139_);
  and (_12196_, _09388_, _04623_);
  nor (_12198_, _12196_, _12161_);
  nor (_12199_, _12198_, _03139_);
  or (_12201_, _12199_, _06549_);
  or (_12202_, _12201_, _12195_);
  and (_12204_, _09404_, _04623_);
  or (_12205_, _12161_, _05305_);
  or (_12207_, _12205_, _12204_);
  and (_12208_, _04623_, _09395_);
  nor (_12210_, _12208_, _12161_);
  and (_12211_, _12210_, _02575_);
  nor (_12213_, _12211_, _03251_);
  and (_12214_, _12213_, _12207_);
  and (_12216_, _12214_, _12202_);
  nor (_12217_, _12216_, _12164_);
  nor (_12219_, _12217_, _02669_);
  nor (_12220_, _12161_, _06119_);
  not (_12222_, _12220_);
  nor (_12223_, _12210_, _05332_);
  and (_12224_, _12223_, _12222_);
  nor (_12225_, _12224_, _12219_);
  nor (_12226_, _12225_, _03243_);
  or (_12227_, _12220_, _03244_);
  nor (_12228_, _12227_, _12169_);
  or (_12229_, _12228_, _02654_);
  nor (_12230_, _12229_, _12226_);
  nor (_12231_, _09403_, _06956_);
  nor (_12232_, _12231_, _12161_);
  and (_12233_, _12232_, _02654_);
  nor (_12234_, _12233_, _12230_);
  and (_12235_, _12234_, _05883_);
  nor (_12236_, _09267_, _06956_);
  nor (_12237_, _12236_, _12161_);
  nor (_12238_, _12237_, _05883_);
  or (_12239_, _12238_, _12235_);
  and (_12240_, _12239_, _03124_);
  nor (_12241_, _12175_, _03124_);
  or (_12242_, _12241_, _12240_);
  and (_12243_, _12242_, _03513_);
  and (_12244_, _09456_, _04623_);
  nor (_12245_, _12244_, _12161_);
  nor (_12246_, _12245_, _03513_);
  or (_12247_, _12246_, _12243_);
  or (_12248_, _12247_, _27789_);
  or (_12249_, _27788_, \oc8051_golden_model_1.PCON [6]);
  and (_12250_, _12249_, _27053_);
  and (_28876_, _12250_, _12248_);
  not (_12251_, \oc8051_golden_model_1.SBUF [0]);
  nor (_12252_, _04626_, _12251_);
  nor (_12253_, _04888_, _06866_);
  nor (_12254_, _12253_, _12252_);
  and (_12255_, _12254_, _11672_);
  and (_12256_, _04626_, \oc8051_golden_model_1.ACC [0]);
  nor (_12257_, _12256_, _12252_);
  nor (_12258_, _12257_, _03179_);
  nor (_12259_, _12258_, _05949_);
  nor (_12260_, _12254_, _02662_);
  nor (_12261_, _04505_, _12251_);
  nor (_12262_, _12257_, _05903_);
  nor (_12263_, _12262_, _12261_);
  nor (_12264_, _12263_, _02661_);
  or (_12265_, _12264_, _03162_);
  nor (_12266_, _12265_, _12260_);
  or (_12267_, _12266_, _03168_);
  and (_12268_, _12267_, _12259_);
  and (_12269_, _04626_, _03716_);
  nor (_12270_, _05949_, _03162_);
  or (_12271_, _12270_, _12252_);
  nor (_12272_, _12271_, _12269_);
  nor (_12273_, _12272_, _12268_);
  nor (_12274_, _12273_, _05959_);
  and (_12275_, _04626_, _04268_);
  nor (_12276_, _12252_, _05963_);
  not (_12277_, _12276_);
  nor (_12278_, _12277_, _12275_);
  nor (_12279_, _12278_, _12274_);
  nor (_12280_, _12279_, _02024_);
  nor (_12281_, _08093_, _06866_);
  or (_12282_, _12252_, _03139_);
  nor (_12283_, _12282_, _12281_);
  or (_12284_, _12283_, _02575_);
  nor (_12285_, _12284_, _12280_);
  and (_12286_, _04626_, _05996_);
  nor (_12287_, _12286_, _12252_);
  nand (_12288_, _12287_, _05305_);
  and (_12289_, _12288_, _06549_);
  nor (_12290_, _12289_, _12285_);
  and (_12291_, _07968_, _04626_);
  nor (_12292_, _12291_, _12252_);
  and (_12293_, _12292_, _02656_);
  nor (_12294_, _12293_, _12290_);
  and (_12295_, _12294_, _03252_);
  and (_12296_, _08110_, _04626_);
  nor (_12297_, _12296_, _12252_);
  nor (_12298_, _12297_, _03252_);
  or (_12299_, _12298_, _12295_);
  and (_12300_, _12299_, _05332_);
  or (_12301_, _12287_, _05332_);
  nor (_12302_, _12301_, _12253_);
  nor (_12303_, _12302_, _12300_);
  nor (_12304_, _12303_, _03243_);
  and (_12305_, _08108_, _04626_);
  or (_12306_, _12305_, _12252_);
  and (_12307_, _12306_, _03243_);
  or (_12308_, _12307_, _12304_);
  and (_12309_, _12308_, _05357_);
  nor (_12310_, _07967_, _06866_);
  nor (_12311_, _12310_, _12252_);
  nor (_12312_, _12311_, _05357_);
  or (_12313_, _12312_, _12309_);
  and (_12314_, _12313_, _05883_);
  nor (_12315_, _08109_, _06866_);
  nor (_12316_, _12315_, _12252_);
  nor (_12317_, _12316_, _05883_);
  nor (_12318_, _12317_, _11672_);
  not (_12319_, _12318_);
  nor (_12320_, _12319_, _12314_);
  nor (_12321_, _12320_, _12255_);
  or (_12322_, _12321_, _27789_);
  or (_12323_, _27788_, \oc8051_golden_model_1.SBUF [0]);
  and (_12324_, _12323_, _27053_);
  and (_28877_, _12324_, _12322_);
  nor (_12325_, _04626_, \oc8051_golden_model_1.SBUF [1]);
  and (_12326_, _08209_, _04626_);
  nor (_12327_, _12326_, _12325_);
  nor (_12328_, _12327_, _03124_);
  not (_12329_, _12325_);
  nor (_12330_, _08325_, _06866_);
  nor (_12331_, _12330_, _03252_);
  and (_12332_, _12331_, _12329_);
  and (_12333_, _04626_, _04218_);
  not (_12334_, \oc8051_golden_model_1.SBUF [1]);
  nor (_12335_, _04626_, _12334_);
  nor (_12336_, _12335_, _05963_);
  not (_12337_, _12336_);
  nor (_12338_, _12337_, _12333_);
  not (_12339_, _12338_);
  and (_12340_, _04626_, _08322_);
  nor (_12341_, _12340_, _12325_);
  and (_12342_, _12341_, _03168_);
  and (_12343_, _12341_, _04505_);
  nor (_12344_, _04505_, _12334_);
  or (_12345_, _12344_, _12343_);
  and (_12346_, _12345_, _02662_);
  and (_12347_, _12327_, _02661_);
  or (_12348_, _12347_, _12346_);
  and (_12349_, _12348_, _03365_);
  nor (_12350_, _06866_, _03777_);
  nor (_12351_, _12350_, _12335_);
  nor (_12352_, _12351_, _03365_);
  nor (_12353_, _12352_, _12349_);
  nor (_12354_, _12353_, _03168_);
  or (_12355_, _12354_, _05949_);
  nor (_12356_, _12355_, _12342_);
  and (_12357_, _12351_, _05949_);
  nor (_12358_, _12357_, _12356_);
  nor (_12359_, _12358_, _05959_);
  nor (_12360_, _12359_, _02024_);
  and (_12361_, _12360_, _12339_);
  and (_12362_, _08307_, _04626_);
  nor (_12363_, _12362_, _03139_);
  and (_12364_, _12363_, _12329_);
  nor (_12365_, _12364_, _12361_);
  nor (_12366_, _12365_, _06549_);
  nor (_12367_, _08185_, _06866_);
  nor (_12368_, _12367_, _05305_);
  and (_12369_, _04626_, _03016_);
  nor (_12370_, _12369_, _05245_);
  or (_12371_, _12370_, _12368_);
  and (_12372_, _12371_, _12329_);
  nor (_12373_, _12372_, _12366_);
  nor (_12374_, _12373_, _03251_);
  nor (_12375_, _12374_, _12332_);
  nor (_12376_, _12375_, _02669_);
  nor (_12377_, _08184_, _06866_);
  nor (_12378_, _12377_, _05332_);
  and (_12379_, _12378_, _12329_);
  nor (_12380_, _12379_, _12376_);
  nor (_12381_, _12380_, _03243_);
  nor (_12382_, _12335_, _06122_);
  nor (_12383_, _12382_, _03244_);
  and (_12384_, _12383_, _12341_);
  nor (_12385_, _12384_, _12381_);
  nor (_12386_, _12385_, _03241_);
  and (_12387_, _12369_, _04835_);
  nor (_12388_, _12387_, _05357_);
  and (_12389_, _12340_, _04835_);
  nor (_12390_, _12389_, _05883_);
  or (_12391_, _12390_, _12388_);
  and (_12392_, _12391_, _12329_);
  or (_12393_, _12392_, _03123_);
  nor (_12394_, _12393_, _12386_);
  nor (_12395_, _12394_, _12328_);
  nor (_12396_, _12395_, _03121_);
  nor (_12397_, _12335_, _12326_);
  and (_12398_, _12397_, _03121_);
  nor (_12399_, _12398_, _12396_);
  or (_12400_, _12399_, _27789_);
  or (_12401_, _27788_, \oc8051_golden_model_1.SBUF [1]);
  and (_12402_, _12401_, _27053_);
  and (_28878_, _12402_, _12400_);
  not (_12403_, \oc8051_golden_model_1.SBUF [2]);
  nor (_12404_, _04626_, _12403_);
  and (_12405_, _04626_, _04170_);
  nor (_12406_, _12405_, _12404_);
  or (_12407_, _12406_, _05963_);
  and (_12408_, _04626_, \oc8051_golden_model_1.ACC [2]);
  nor (_12409_, _12408_, _12404_);
  nor (_12410_, _12409_, _03179_);
  nor (_12411_, _12409_, _05903_);
  nor (_12412_, _04505_, _12403_);
  or (_12413_, _12412_, _12411_);
  and (_12414_, _12413_, _02662_);
  nor (_12415_, _08420_, _06866_);
  nor (_12416_, _12415_, _12404_);
  nor (_12417_, _12416_, _02662_);
  or (_12418_, _12417_, _12414_);
  and (_12419_, _12418_, _03365_);
  nor (_12420_, _06866_, _03644_);
  nor (_12421_, _12420_, _12404_);
  nor (_12422_, _12421_, _03365_);
  nor (_12423_, _12422_, _12419_);
  nor (_12424_, _12423_, _03168_);
  or (_12425_, _12424_, _05949_);
  nor (_12426_, _12425_, _12410_);
  and (_12427_, _12421_, _05949_);
  or (_12428_, _12427_, _05959_);
  or (_12429_, _12428_, _12426_);
  and (_12430_, _12429_, _03139_);
  and (_12431_, _12430_, _12407_);
  nor (_12432_, _08522_, _06866_);
  or (_12433_, _12404_, _03139_);
  nor (_12434_, _12433_, _12432_);
  or (_12435_, _12434_, _02575_);
  nor (_12436_, _12435_, _12431_);
  and (_12437_, _04626_, _06009_);
  nor (_12438_, _12437_, _12404_);
  nand (_12439_, _12438_, _05305_);
  and (_12440_, _12439_, _06549_);
  nor (_12441_, _12440_, _12436_);
  and (_12442_, _08537_, _04626_);
  nor (_12443_, _12442_, _12404_);
  and (_12444_, _12443_, _02656_);
  nor (_12445_, _12444_, _12441_);
  and (_12446_, _12445_, _03252_);
  and (_12447_, _08387_, _04626_);
  nor (_12448_, _12447_, _12404_);
  nor (_12449_, _12448_, _03252_);
  or (_12450_, _12449_, _12446_);
  and (_12451_, _12450_, _05332_);
  nor (_12452_, _12404_, _06121_);
  not (_12453_, _12452_);
  nor (_12454_, _12438_, _05332_);
  and (_12455_, _12454_, _12453_);
  nor (_12456_, _12455_, _12451_);
  nor (_12457_, _12456_, _03243_);
  or (_12458_, _12452_, _03244_);
  nor (_12459_, _12458_, _12409_);
  or (_12460_, _12459_, _02654_);
  nor (_12461_, _12460_, _12457_);
  nor (_12462_, _08536_, _06866_);
  nor (_12463_, _12462_, _12404_);
  and (_12464_, _12463_, _02654_);
  nor (_12465_, _12464_, _12461_);
  and (_12466_, _12465_, _05883_);
  nor (_12467_, _08386_, _06866_);
  nor (_12468_, _12467_, _12404_);
  nor (_12469_, _12468_, _05883_);
  or (_12470_, _12469_, _12466_);
  and (_12471_, _12470_, _03124_);
  nor (_12472_, _12416_, _03124_);
  or (_12473_, _12472_, _12471_);
  and (_12474_, _12473_, _03513_);
  and (_12475_, _08596_, _04626_);
  nor (_12476_, _12475_, _12404_);
  nor (_12477_, _12476_, _03513_);
  or (_12478_, _12477_, _12474_);
  or (_12479_, _12478_, _27789_);
  or (_12480_, _27788_, \oc8051_golden_model_1.SBUF [2]);
  and (_12481_, _12480_, _27053_);
  and (_28879_, _12481_, _12479_);
  not (_12482_, \oc8051_golden_model_1.SBUF [3]);
  nor (_12483_, _04626_, _12482_);
  nor (_12484_, _12483_, _06120_);
  not (_12485_, _12484_);
  and (_12486_, _04626_, _05986_);
  nor (_12487_, _12486_, _12483_);
  nor (_12488_, _12487_, _05332_);
  and (_12489_, _12488_, _12485_);
  and (_12490_, _04626_, \oc8051_golden_model_1.ACC [3]);
  nor (_12491_, _12490_, _12483_);
  nor (_12492_, _12491_, _05903_);
  nor (_12493_, _04505_, _12482_);
  or (_12494_, _12493_, _12492_);
  and (_12495_, _12494_, _02662_);
  nor (_12496_, _08646_, _06866_);
  nor (_12497_, _12496_, _12483_);
  nor (_12498_, _12497_, _02662_);
  or (_12499_, _12498_, _12495_);
  and (_12500_, _12499_, _03365_);
  nor (_12501_, _06866_, _03859_);
  nor (_12502_, _12501_, _12483_);
  nor (_12503_, _12502_, _03365_);
  nor (_12504_, _12503_, _12500_);
  nor (_12505_, _12504_, _03168_);
  nor (_12506_, _12491_, _03179_);
  nor (_12507_, _12506_, _05949_);
  not (_12508_, _12507_);
  nor (_12509_, _12508_, _12505_);
  and (_12510_, _12502_, _05949_);
  or (_12511_, _12510_, _05959_);
  or (_12512_, _12511_, _12509_);
  and (_12513_, _04626_, _04120_);
  nor (_12514_, _12513_, _12483_);
  or (_12515_, _12514_, _05963_);
  and (_12516_, _12515_, _03139_);
  and (_12517_, _12516_, _12512_);
  nor (_12518_, _08744_, _06866_);
  or (_12519_, _12483_, _03139_);
  nor (_12520_, _12519_, _12518_);
  or (_12521_, _12520_, _02575_);
  nor (_12522_, _12521_, _12517_);
  nand (_12523_, _12487_, _05305_);
  and (_12524_, _12523_, _06549_);
  nor (_12525_, _12524_, _12522_);
  and (_12526_, _08622_, _04626_);
  nor (_12527_, _12526_, _12483_);
  and (_12528_, _12527_, _02656_);
  nor (_12529_, _12528_, _12525_);
  and (_12530_, _12529_, _03252_);
  and (_12531_, _08618_, _04626_);
  nor (_12532_, _12531_, _12483_);
  nor (_12533_, _12532_, _03252_);
  or (_12534_, _12533_, _12530_);
  and (_12535_, _12534_, _05332_);
  nor (_12536_, _12535_, _12489_);
  nor (_12537_, _12536_, _03243_);
  or (_12538_, _12484_, _03244_);
  nor (_12539_, _12538_, _12491_);
  or (_12540_, _12539_, _02654_);
  nor (_12541_, _12540_, _12537_);
  nor (_12542_, _08621_, _06866_);
  nor (_12543_, _12542_, _12483_);
  and (_12544_, _12543_, _02654_);
  nor (_12545_, _12544_, _12541_);
  and (_12546_, _12545_, _05883_);
  nor (_12547_, _08617_, _06866_);
  nor (_12548_, _12547_, _12483_);
  nor (_12549_, _12548_, _05883_);
  or (_12550_, _12549_, _12546_);
  and (_12551_, _12550_, _03124_);
  nor (_12552_, _12497_, _03124_);
  or (_12553_, _12552_, _12551_);
  and (_12554_, _12553_, _03513_);
  and (_12555_, _08807_, _04626_);
  nor (_12556_, _12555_, _12483_);
  nor (_12557_, _12556_, _03513_);
  or (_12558_, _12557_, _12554_);
  or (_12559_, _12558_, _27789_);
  or (_12560_, _27788_, \oc8051_golden_model_1.SBUF [3]);
  and (_12561_, _12560_, _27053_);
  and (_28880_, _12561_, _12559_);
  not (_12562_, \oc8051_golden_model_1.SBUF [4]);
  nor (_12563_, _04626_, _12562_);
  and (_12564_, _08830_, _04626_);
  nor (_12565_, _12564_, _12563_);
  nor (_12566_, _12565_, _03252_);
  and (_12567_, _04626_, _05974_);
  nor (_12568_, _12567_, _12563_);
  and (_12569_, _12568_, _02575_);
  and (_12570_, _04626_, \oc8051_golden_model_1.ACC [4]);
  nor (_12571_, _12570_, _12563_);
  nor (_12572_, _12571_, _03179_);
  nor (_12573_, _12571_, _05903_);
  nor (_12574_, _04505_, _12562_);
  or (_12575_, _12574_, _12573_);
  and (_12576_, _12575_, _02662_);
  nor (_12577_, _08838_, _06866_);
  nor (_12578_, _12577_, _12563_);
  nor (_12579_, _12578_, _02662_);
  or (_12580_, _12579_, _12576_);
  and (_12581_, _12580_, _03365_);
  nor (_12582_, _06866_, _04325_);
  nor (_12583_, _12582_, _12563_);
  nor (_12584_, _12583_, _03365_);
  nor (_12585_, _12584_, _12581_);
  nor (_12586_, _12585_, _03168_);
  or (_12587_, _12586_, _05949_);
  nor (_12588_, _12587_, _12572_);
  and (_12589_, _12583_, _05949_);
  nor (_12590_, _12589_, _12588_);
  nor (_12591_, _12590_, _05959_);
  and (_12592_, _04626_, _04012_);
  nor (_12593_, _12563_, _05963_);
  not (_12594_, _12593_);
  nor (_12595_, _12594_, _12592_);
  or (_12596_, _12595_, _02024_);
  nor (_12597_, _12596_, _12591_);
  nor (_12598_, _08967_, _06866_);
  nor (_12599_, _12598_, _12563_);
  nor (_12600_, _12599_, _03139_);
  or (_12601_, _12600_, _02575_);
  nor (_12602_, _12601_, _12597_);
  nor (_12603_, _12602_, _12569_);
  or (_12604_, _12603_, _02656_);
  and (_12605_, _08982_, _04626_);
  or (_12606_, _12605_, _12563_);
  or (_12607_, _12606_, _05305_);
  and (_12608_, _12607_, _03252_);
  and (_12609_, _12608_, _12604_);
  nor (_12610_, _12609_, _12566_);
  nor (_12611_, _12610_, _02669_);
  nor (_12612_, _12563_, _09034_);
  not (_12613_, _12612_);
  nor (_12614_, _12568_, _05332_);
  and (_12615_, _12614_, _12613_);
  nor (_12616_, _12615_, _12611_);
  nor (_12617_, _12616_, _03243_);
  or (_12618_, _12612_, _03244_);
  nor (_12619_, _12618_, _12571_);
  or (_12620_, _12619_, _02654_);
  nor (_12621_, _12620_, _12617_);
  nor (_12622_, _08981_, _06866_);
  nor (_12623_, _12622_, _12563_);
  and (_12624_, _12623_, _02654_);
  nor (_12625_, _12624_, _12621_);
  and (_12626_, _12625_, _05883_);
  nor (_12627_, _08828_, _06866_);
  nor (_12628_, _12627_, _12563_);
  nor (_12629_, _12628_, _05883_);
  or (_12630_, _12629_, _12626_);
  and (_12631_, _12630_, _03124_);
  nor (_12632_, _12578_, _03124_);
  or (_12633_, _12632_, _12631_);
  and (_12634_, _12633_, _03513_);
  and (_12635_, _09037_, _04626_);
  nor (_12636_, _12635_, _12563_);
  nor (_12637_, _12636_, _03513_);
  or (_12638_, _12637_, _12634_);
  or (_12639_, _12638_, _27789_);
  or (_12640_, _27788_, \oc8051_golden_model_1.SBUF [4]);
  and (_12641_, _12640_, _27053_);
  and (_28881_, _12641_, _12639_);
  not (_12642_, \oc8051_golden_model_1.SBUF [5]);
  nor (_12643_, _04626_, _12642_);
  and (_12644_, _09055_, _04626_);
  nor (_12645_, _12644_, _12643_);
  nor (_12646_, _12645_, _03252_);
  and (_12647_, _04626_, _06036_);
  nor (_12648_, _12647_, _12643_);
  and (_12649_, _12648_, _02575_);
  nor (_12650_, _06866_, _04480_);
  nor (_12651_, _12650_, _12643_);
  and (_12652_, _12651_, _05949_);
  and (_12653_, _04626_, \oc8051_golden_model_1.ACC [5]);
  nor (_12654_, _12653_, _12643_);
  nor (_12655_, _12654_, _05903_);
  nor (_12656_, _04505_, _12642_);
  or (_12657_, _12656_, _12655_);
  and (_12658_, _12657_, _02662_);
  nor (_12659_, _09087_, _06866_);
  nor (_12660_, _12659_, _12643_);
  nor (_12661_, _12660_, _02662_);
  or (_12662_, _12661_, _12658_);
  and (_12663_, _12662_, _03365_);
  nor (_12664_, _12651_, _03365_);
  nor (_12665_, _12664_, _12663_);
  nor (_12666_, _12665_, _03168_);
  nor (_12667_, _12654_, _03179_);
  nor (_12668_, _12667_, _05949_);
  not (_12669_, _12668_);
  nor (_12670_, _12669_, _12666_);
  nor (_12671_, _12670_, _12652_);
  nor (_12672_, _12671_, _05959_);
  and (_12673_, _04626_, _03904_);
  nor (_12674_, _12643_, _05963_);
  not (_12675_, _12674_);
  nor (_12676_, _12675_, _12673_);
  or (_12677_, _12676_, _02024_);
  nor (_12678_, _12677_, _12672_);
  nor (_12679_, _09180_, _06866_);
  nor (_12680_, _12679_, _12643_);
  nor (_12681_, _12680_, _03139_);
  or (_12682_, _12681_, _02575_);
  nor (_12683_, _12682_, _12678_);
  nor (_12684_, _12683_, _12649_);
  or (_12685_, _12684_, _02656_);
  and (_12686_, _09195_, _04626_);
  or (_12687_, _12686_, _12643_);
  or (_12688_, _12687_, _05305_);
  and (_12689_, _12688_, _03252_);
  and (_12690_, _12689_, _12685_);
  nor (_12691_, _12690_, _12646_);
  nor (_12692_, _12691_, _02669_);
  not (_12693_, _12643_);
  and (_12694_, _12693_, _04787_);
  not (_12695_, _12694_);
  nor (_12696_, _12648_, _05332_);
  and (_12697_, _12696_, _12695_);
  nor (_12698_, _12697_, _12692_);
  nor (_12699_, _12698_, _03243_);
  or (_12700_, _12694_, _03244_);
  nor (_12701_, _12700_, _12654_);
  or (_12702_, _12701_, _02654_);
  nor (_12703_, _12702_, _12699_);
  nor (_12704_, _09194_, _06866_);
  nor (_12705_, _12704_, _12643_);
  and (_12706_, _12705_, _02654_);
  nor (_12707_, _12706_, _12703_);
  and (_12708_, _12707_, _05883_);
  nor (_12709_, _09054_, _06866_);
  nor (_12710_, _12709_, _12643_);
  nor (_12711_, _12710_, _05883_);
  or (_12712_, _12711_, _12708_);
  and (_12713_, _12712_, _03124_);
  nor (_12714_, _12660_, _03124_);
  or (_12715_, _12714_, _12713_);
  and (_12716_, _12715_, _03513_);
  and (_12717_, _09248_, _04626_);
  nor (_12718_, _12717_, _12643_);
  nor (_12719_, _12718_, _03513_);
  or (_12720_, _12719_, _12716_);
  or (_12721_, _12720_, _27789_);
  or (_12722_, _27788_, \oc8051_golden_model_1.SBUF [5]);
  and (_12723_, _12722_, _27053_);
  and (_28882_, _12723_, _12721_);
  not (_12724_, \oc8051_golden_model_1.SBUF [6]);
  nor (_12725_, _04626_, _12724_);
  and (_12726_, _09268_, _04626_);
  nor (_12727_, _12726_, _12725_);
  nor (_12728_, _12727_, _03252_);
  and (_12729_, _04626_, _03960_);
  or (_12730_, _12729_, _12725_);
  and (_12731_, _12730_, _05959_);
  and (_12732_, _04626_, \oc8051_golden_model_1.ACC [6]);
  nor (_12733_, _12732_, _12725_);
  nor (_12734_, _12733_, _03179_);
  nor (_12735_, _12733_, _05903_);
  nor (_12736_, _04505_, _12724_);
  or (_12737_, _12736_, _12735_);
  and (_12738_, _12737_, _02662_);
  nor (_12739_, _09301_, _06866_);
  nor (_12740_, _12739_, _12725_);
  nor (_12741_, _12740_, _02662_);
  or (_12742_, _12741_, _12738_);
  and (_12743_, _12742_, _03365_);
  nor (_12744_, _06866_, _04373_);
  nor (_12745_, _12744_, _12725_);
  nor (_12746_, _12745_, _03365_);
  nor (_12747_, _12746_, _12743_);
  nor (_12748_, _12747_, _03168_);
  or (_12749_, _12748_, _05949_);
  nor (_12750_, _12749_, _12734_);
  and (_12751_, _12745_, _05949_);
  or (_12752_, _12751_, _05959_);
  nor (_12753_, _12752_, _12750_);
  or (_12754_, _12753_, _12731_);
  and (_12755_, _12754_, _03139_);
  and (_12756_, _09388_, _04626_);
  nor (_12757_, _12756_, _12725_);
  nor (_12758_, _12757_, _03139_);
  or (_12759_, _12758_, _06549_);
  or (_12760_, _12759_, _12755_);
  and (_12761_, _09404_, _04626_);
  or (_12762_, _12725_, _05305_);
  or (_12763_, _12762_, _12761_);
  and (_12764_, _04626_, _09395_);
  nor (_12765_, _12764_, _12725_);
  and (_12766_, _12765_, _02575_);
  nor (_12767_, _12766_, _03251_);
  and (_12768_, _12767_, _12763_);
  and (_12769_, _12768_, _12760_);
  nor (_12770_, _12769_, _12728_);
  nor (_12771_, _12770_, _02669_);
  nor (_12772_, _12725_, _06119_);
  not (_12773_, _12772_);
  nor (_12774_, _12765_, _05332_);
  and (_12775_, _12774_, _12773_);
  nor (_12776_, _12775_, _12771_);
  nor (_12777_, _12776_, _03243_);
  or (_12778_, _12772_, _03244_);
  nor (_12779_, _12778_, _12733_);
  or (_12780_, _12779_, _02654_);
  nor (_12781_, _12780_, _12777_);
  nor (_12782_, _09403_, _06866_);
  nor (_12783_, _12782_, _12725_);
  and (_12784_, _12783_, _02654_);
  nor (_12785_, _12784_, _12781_);
  and (_12786_, _12785_, _05883_);
  nor (_12787_, _09267_, _06866_);
  nor (_12788_, _12787_, _12725_);
  nor (_12789_, _12788_, _05883_);
  or (_12790_, _12789_, _12786_);
  and (_12791_, _12790_, _03124_);
  nor (_12792_, _12740_, _03124_);
  or (_12793_, _12792_, _12791_);
  and (_12794_, _12793_, _03513_);
  and (_12795_, _09456_, _04626_);
  nor (_12796_, _12795_, _12725_);
  nor (_12797_, _12796_, _03513_);
  or (_12798_, _12797_, _12794_);
  or (_12799_, _12798_, _27789_);
  or (_12800_, _27788_, \oc8051_golden_model_1.SBUF [6]);
  and (_12801_, _12800_, _27053_);
  and (_28883_, _12801_, _12799_);
  not (_12802_, \oc8051_golden_model_1.SCON [0]);
  nor (_12803_, _04615_, _12802_);
  nor (_12804_, _04888_, _06755_);
  nor (_12805_, _12804_, _12803_);
  nor (_12806_, _12805_, _03513_);
  and (_12807_, _04615_, _04268_);
  nor (_12808_, _12803_, _05963_);
  not (_12809_, _12808_);
  nor (_12810_, _12809_, _12807_);
  nor (_12811_, _05431_, _12802_);
  and (_12812_, _07997_, _05431_);
  nor (_12813_, _12812_, _12811_);
  nor (_12814_, _12813_, _03390_);
  and (_12815_, _12805_, _02661_);
  and (_12816_, _04615_, \oc8051_golden_model_1.ACC [0]);
  nor (_12817_, _12816_, _12803_);
  nor (_12818_, _12817_, _05903_);
  nor (_12819_, _04505_, _12802_);
  or (_12820_, _12819_, _02661_);
  nor (_12821_, _12820_, _12818_);
  or (_12822_, _12821_, _06504_);
  nor (_12823_, _12822_, _12815_);
  and (_12824_, _04615_, _03716_);
  nor (_12825_, _12824_, _12803_);
  nor (_12826_, _12825_, _03365_);
  or (_12827_, _12826_, _03168_);
  or (_12828_, _12827_, _12823_);
  nor (_12829_, _12828_, _12814_);
  and (_12830_, _12817_, _03168_);
  nor (_12831_, _12830_, _03176_);
  not (_12832_, _12831_);
  nor (_12833_, _12832_, _12829_);
  and (_12834_, _12803_, _03176_);
  or (_12835_, _12834_, _12833_);
  and (_12836_, _12835_, _05168_);
  nor (_12837_, _12805_, _05168_);
  or (_12838_, _12837_, _12836_);
  nor (_12839_, _12838_, _03140_);
  nor (_12840_, _08035_, _06792_);
  or (_12841_, _12811_, _03141_);
  nor (_12842_, _12841_, _12840_);
  or (_12843_, _12842_, _05949_);
  or (_12844_, _12843_, _12839_);
  or (_12845_, _12825_, _06673_);
  and (_12846_, _12845_, _05963_);
  and (_12847_, _12846_, _12844_);
  nor (_12848_, _12847_, _12810_);
  nor (_12849_, _12848_, _02024_);
  nor (_12850_, _08093_, _06755_);
  or (_12851_, _12803_, _03139_);
  nor (_12852_, _12851_, _12850_);
  or (_12853_, _12852_, _02575_);
  nor (_12854_, _12853_, _12849_);
  and (_12855_, _04615_, _05996_);
  nor (_12856_, _12855_, _12803_);
  nand (_12857_, _12856_, _05305_);
  and (_12858_, _12857_, _06549_);
  nor (_12859_, _12858_, _12854_);
  and (_12860_, _07968_, _04615_);
  nor (_12861_, _12860_, _12803_);
  and (_12862_, _12861_, _02656_);
  nor (_12863_, _12862_, _12859_);
  and (_12864_, _12863_, _03252_);
  and (_12865_, _08110_, _04615_);
  nor (_12866_, _12865_, _12803_);
  nor (_12867_, _12866_, _03252_);
  or (_12868_, _12867_, _12864_);
  and (_12869_, _12868_, _05332_);
  or (_12870_, _12856_, _05332_);
  nor (_12871_, _12870_, _12804_);
  nor (_12872_, _12871_, _12869_);
  nor (_12873_, _12872_, _03243_);
  nor (_12874_, _12803_, _04888_);
  or (_12875_, _12874_, _03244_);
  nor (_12876_, _12875_, _12817_);
  or (_12877_, _12876_, _02654_);
  nor (_12878_, _12877_, _12873_);
  nor (_12879_, _07967_, _06755_);
  nor (_12880_, _12879_, _12803_);
  and (_12881_, _12880_, _02654_);
  nor (_12882_, _12881_, _12878_);
  and (_12883_, _12882_, _05883_);
  nor (_12884_, _08109_, _06755_);
  nor (_12885_, _12884_, _12803_);
  nor (_12886_, _12885_, _05883_);
  or (_12887_, _12886_, _12883_);
  and (_12888_, _12887_, _03124_);
  nor (_12889_, _12805_, _03124_);
  nor (_12890_, _12889_, _02650_);
  not (_12891_, _12890_);
  nor (_12892_, _12891_, _12888_);
  nor (_12893_, _12803_, _03122_);
  nor (_12894_, _12893_, _12892_);
  and (_12895_, _12894_, _03513_);
  nor (_12896_, _12895_, _12806_);
  nand (_12897_, _12896_, _27788_);
  or (_12898_, _27788_, \oc8051_golden_model_1.SCON [0]);
  and (_12899_, _12898_, _27053_);
  and (_28886_, _12899_, _12897_);
  nor (_12900_, _04615_, \oc8051_golden_model_1.SCON [1]);
  not (_12901_, _12900_);
  nor (_12902_, _08325_, _06755_);
  nor (_12903_, _12902_, _03252_);
  and (_12904_, _12903_, _12901_);
  not (_12905_, \oc8051_golden_model_1.SCON [1]);
  nor (_12906_, _04615_, _12905_);
  and (_12907_, _04615_, _04218_);
  or (_12908_, _12907_, _12906_);
  and (_12909_, _12908_, _05959_);
  nor (_12910_, _08246_, _06792_);
  nor (_12911_, _05431_, _12905_);
  or (_12912_, _12911_, _03141_);
  or (_12913_, _12912_, _12910_);
  and (_12914_, _08209_, _04615_);
  nor (_12915_, _12914_, _12900_);
  nor (_12916_, _12915_, _02662_);
  and (_12917_, _04615_, _08322_);
  nor (_12918_, _12917_, _12900_);
  and (_12919_, _12918_, _04505_);
  nor (_12920_, _04505_, _12905_);
  or (_12921_, _12920_, _02661_);
  nor (_12922_, _12921_, _12919_);
  or (_12923_, _12922_, _06504_);
  nor (_12924_, _12923_, _12916_);
  nor (_12925_, _06755_, _03777_);
  nor (_12926_, _12925_, _12906_);
  nor (_12927_, _12926_, _03365_);
  and (_12928_, _08213_, _05431_);
  nor (_12929_, _12928_, _12911_);
  nor (_12930_, _12929_, _03390_);
  nor (_12931_, _12930_, _12927_);
  nand (_12932_, _12931_, _03179_);
  or (_12933_, _12932_, _12924_);
  or (_12934_, _12918_, _03179_);
  and (_12935_, _12934_, _12933_);
  and (_12936_, _12935_, _03177_);
  and (_12937_, _08200_, _05431_);
  nor (_12938_, _12937_, _12911_);
  nor (_12939_, _12938_, _03177_);
  or (_12940_, _12939_, _12936_);
  and (_12941_, _12940_, _05168_);
  nor (_12942_, _12911_, _08228_);
  or (_12943_, _12942_, _05168_);
  nor (_12944_, _12943_, _12929_);
  or (_12945_, _12944_, _03140_);
  or (_12946_, _12945_, _12941_);
  and (_12947_, _12946_, _12913_);
  nor (_12948_, _12947_, _05949_);
  and (_12949_, _12926_, _05949_);
  or (_12950_, _12949_, _05959_);
  nor (_12951_, _12950_, _12948_);
  or (_12952_, _12951_, _12909_);
  and (_12953_, _12952_, _03139_);
  nor (_12954_, _08307_, _06755_);
  nor (_12955_, _12954_, _12906_);
  nor (_12956_, _12955_, _03139_);
  nor (_12957_, _12956_, _12953_);
  nor (_12958_, _12957_, _06549_);
  nor (_12959_, _08185_, _06755_);
  nor (_12960_, _12959_, _05305_);
  and (_12961_, _04615_, _03016_);
  nor (_12962_, _12961_, _05245_);
  or (_12963_, _12962_, _12960_);
  and (_12964_, _12963_, _12901_);
  nor (_12965_, _12964_, _12958_);
  nor (_12966_, _12965_, _03251_);
  nor (_12967_, _12966_, _12904_);
  nor (_12968_, _12967_, _02669_);
  nor (_12969_, _08184_, _06755_);
  nor (_12970_, _12969_, _05332_);
  and (_12971_, _12970_, _12901_);
  nor (_12972_, _12971_, _12968_);
  nor (_12973_, _12972_, _03243_);
  nor (_12974_, _12906_, _06122_);
  nor (_12975_, _12974_, _03244_);
  and (_12976_, _12975_, _12918_);
  nor (_12977_, _12976_, _12973_);
  nor (_12978_, _12977_, _03241_);
  and (_12979_, _12961_, _04835_);
  nor (_12980_, _12979_, _05357_);
  nand (_12981_, _12917_, _04835_);
  and (_12982_, _12981_, _03239_);
  or (_12983_, _12982_, _12980_);
  and (_12984_, _12983_, _12901_);
  or (_12985_, _12984_, _03123_);
  nor (_12986_, _12985_, _12978_);
  nor (_12987_, _12915_, _03124_);
  or (_12988_, _12987_, _02650_);
  nor (_12989_, _12988_, _12986_);
  nor (_12990_, _12938_, _03122_);
  or (_12991_, _12990_, _03121_);
  nor (_12992_, _12991_, _12989_);
  nor (_12993_, _12914_, _12906_);
  and (_12994_, _12993_, _03121_);
  nor (_12995_, _12994_, _12992_);
  or (_12996_, _12995_, _27789_);
  or (_12997_, _27788_, \oc8051_golden_model_1.SCON [1]);
  and (_12998_, _12997_, _27053_);
  and (_28887_, _12998_, _12996_);
  not (_12999_, \oc8051_golden_model_1.SCON [2]);
  nor (_13000_, _04615_, _12999_);
  and (_13001_, _04615_, _06009_);
  nor (_13002_, _13001_, _13000_);
  and (_13003_, _13002_, _02575_);
  nor (_13004_, _06755_, _03644_);
  nor (_13005_, _13004_, _13000_);
  and (_13006_, _13005_, _05949_);
  nor (_13007_, _08420_, _06755_);
  nor (_13008_, _13007_, _13000_);
  and (_13009_, _13008_, _02661_);
  and (_13010_, _04615_, \oc8051_golden_model_1.ACC [2]);
  nor (_13011_, _13010_, _13000_);
  nor (_13012_, _13011_, _05903_);
  nor (_13013_, _04505_, _12999_);
  or (_13014_, _13013_, _02661_);
  nor (_13015_, _13014_, _13012_);
  or (_13016_, _13015_, _06504_);
  nor (_13017_, _13016_, _13009_);
  nor (_13018_, _13005_, _03365_);
  nor (_13019_, _05431_, _12999_);
  and (_13020_, _08406_, _05431_);
  nor (_13021_, _13020_, _13019_);
  nor (_13022_, _13021_, _03390_);
  nor (_13023_, _13022_, _13018_);
  nand (_13024_, _13023_, _03179_);
  or (_13025_, _13024_, _13017_);
  nand (_13026_, _13011_, _03168_);
  and (_13027_, _13026_, _13025_);
  nor (_13028_, _13027_, _03176_);
  and (_13029_, _08404_, _05431_);
  nor (_13030_, _13029_, _13019_);
  and (_13031_, _13030_, _03176_);
  or (_13032_, _13031_, _03144_);
  nor (_13033_, _13032_, _13028_);
  nor (_13034_, _13019_, _08446_);
  or (_13035_, _13034_, _05168_);
  nor (_13036_, _13035_, _13021_);
  or (_13037_, _13036_, _13033_);
  and (_13038_, _13037_, _03141_);
  nor (_13039_, _08465_, _06792_);
  nor (_13040_, _13019_, _13039_);
  nor (_13041_, _13040_, _03141_);
  or (_13042_, _13041_, _05949_);
  nor (_13043_, _13042_, _13038_);
  nor (_13044_, _13043_, _13006_);
  nor (_13045_, _13044_, _05959_);
  and (_13046_, _04615_, _04170_);
  nor (_13047_, _13000_, _05963_);
  not (_13048_, _13047_);
  nor (_13049_, _13048_, _13046_);
  or (_13050_, _13049_, _02024_);
  nor (_13051_, _13050_, _13045_);
  nor (_13052_, _08522_, _06755_);
  nor (_13053_, _13052_, _13000_);
  nor (_13054_, _13053_, _03139_);
  or (_13055_, _13054_, _02575_);
  nor (_13056_, _13055_, _13051_);
  nor (_13057_, _13056_, _13003_);
  or (_13058_, _13057_, _02656_);
  and (_13059_, _08537_, _04615_);
  or (_13060_, _13059_, _13000_);
  or (_13061_, _13060_, _05305_);
  and (_13062_, _13061_, _03252_);
  and (_13063_, _13062_, _13058_);
  and (_13064_, _08387_, _04615_);
  nor (_13065_, _13064_, _13000_);
  nor (_13066_, _13065_, _03252_);
  nor (_13067_, _13066_, _13063_);
  nor (_13068_, _13067_, _02669_);
  nor (_13069_, _13000_, _06121_);
  not (_13070_, _13069_);
  nor (_13071_, _13002_, _05332_);
  and (_13072_, _13071_, _13070_);
  nor (_13073_, _13072_, _13068_);
  nor (_13074_, _13073_, _03243_);
  or (_13075_, _13069_, _03244_);
  nor (_13076_, _13075_, _13011_);
  or (_13077_, _13076_, _02654_);
  nor (_13078_, _13077_, _13074_);
  nor (_13079_, _08536_, _06755_);
  nor (_13080_, _13079_, _13000_);
  and (_13081_, _13080_, _02654_);
  nor (_13082_, _13081_, _13078_);
  and (_13083_, _13082_, _05883_);
  nor (_13084_, _08386_, _06755_);
  nor (_13085_, _13084_, _13000_);
  nor (_13086_, _13085_, _05883_);
  or (_13087_, _13086_, _13083_);
  and (_13088_, _13087_, _03124_);
  nor (_13089_, _13008_, _03124_);
  or (_13090_, _13089_, _02650_);
  or (_13091_, _13090_, _13088_);
  nand (_13092_, _13030_, _02650_);
  and (_13093_, _13092_, _13091_);
  nor (_13094_, _13093_, _03121_);
  and (_13095_, _08596_, _04615_);
  nor (_13096_, _13095_, _13000_);
  and (_13097_, _13096_, _03121_);
  nor (_13098_, _13097_, _13094_);
  or (_13099_, _13098_, _27789_);
  or (_13100_, _27788_, \oc8051_golden_model_1.SCON [2]);
  and (_13101_, _13100_, _27053_);
  and (_28888_, _13101_, _13099_);
  not (_13102_, \oc8051_golden_model_1.SCON [3]);
  nor (_13103_, _04615_, _13102_);
  and (_13104_, _04615_, _05986_);
  nor (_13105_, _13104_, _13103_);
  and (_13106_, _13105_, _02575_);
  nor (_13107_, _06755_, _03859_);
  nor (_13108_, _13107_, _13103_);
  and (_13109_, _13108_, _05949_);
  nor (_13110_, _08627_, _06792_);
  nor (_13111_, _05431_, _13102_);
  or (_13112_, _13111_, _03141_);
  or (_13113_, _13112_, _13110_);
  nor (_13114_, _08646_, _06755_);
  nor (_13115_, _13114_, _13103_);
  and (_13116_, _13115_, _02661_);
  and (_13117_, _04615_, \oc8051_golden_model_1.ACC [3]);
  nor (_13118_, _13117_, _13103_);
  nor (_13119_, _13118_, _05903_);
  nor (_13120_, _04505_, _13102_);
  or (_13121_, _13120_, _02661_);
  nor (_13122_, _13121_, _13119_);
  or (_13123_, _13122_, _06504_);
  nor (_13124_, _13123_, _13116_);
  nor (_13125_, _13108_, _03365_);
  and (_13126_, _08642_, _05431_);
  nor (_13127_, _13126_, _13111_);
  nor (_13128_, _13127_, _03390_);
  nor (_13129_, _13128_, _13125_);
  nand (_13130_, _13129_, _03179_);
  or (_13131_, _13130_, _13124_);
  nand (_13132_, _13118_, _03168_);
  and (_13133_, _13132_, _13131_);
  and (_13134_, _13133_, _03177_);
  and (_13135_, _08640_, _05431_);
  nor (_13136_, _13135_, _13111_);
  nor (_13137_, _13136_, _03177_);
  or (_13138_, _13137_, _13134_);
  and (_13139_, _13138_, _05168_);
  nor (_13140_, _13111_, _08671_);
  or (_13141_, _13127_, _05168_);
  nor (_13142_, _13141_, _13140_);
  or (_13143_, _13142_, _03140_);
  or (_13144_, _13143_, _13139_);
  and (_13145_, _13144_, _13113_);
  nor (_13146_, _13145_, _05949_);
  nor (_13147_, _13146_, _13109_);
  nor (_13148_, _13147_, _05959_);
  and (_13149_, _04615_, _04120_);
  nor (_13150_, _13103_, _05963_);
  not (_13151_, _13150_);
  nor (_13152_, _13151_, _13149_);
  or (_13153_, _13152_, _02024_);
  nor (_13154_, _13153_, _13148_);
  nor (_13155_, _08744_, _06755_);
  nor (_13156_, _13155_, _13103_);
  nor (_13157_, _13156_, _03139_);
  or (_13158_, _13157_, _02575_);
  nor (_13159_, _13158_, _13154_);
  nor (_13160_, _13159_, _13106_);
  or (_13161_, _13160_, _02656_);
  and (_13162_, _08622_, _04615_);
  or (_13163_, _13162_, _13103_);
  or (_13164_, _13163_, _05305_);
  and (_13165_, _13164_, _03252_);
  and (_13166_, _13165_, _13161_);
  and (_13167_, _08618_, _04615_);
  nor (_13168_, _13167_, _13103_);
  nor (_13169_, _13168_, _03252_);
  nor (_13170_, _13169_, _13166_);
  nor (_13171_, _13170_, _02669_);
  nor (_13172_, _13103_, _06120_);
  not (_13173_, _13172_);
  nor (_13174_, _13105_, _05332_);
  and (_13175_, _13174_, _13173_);
  nor (_13176_, _13175_, _13171_);
  nor (_13177_, _13176_, _03243_);
  or (_13178_, _13172_, _03244_);
  nor (_13179_, _13178_, _13118_);
  or (_13180_, _13179_, _02654_);
  nor (_13181_, _13180_, _13177_);
  nor (_13182_, _08621_, _06755_);
  nor (_13183_, _13182_, _13103_);
  and (_13184_, _13183_, _02654_);
  nor (_13185_, _13184_, _13181_);
  and (_13186_, _13185_, _05883_);
  nor (_13187_, _08617_, _06755_);
  nor (_13188_, _13187_, _13103_);
  nor (_13189_, _13188_, _05883_);
  or (_13190_, _13189_, _13186_);
  and (_13191_, _13190_, _03124_);
  nor (_13192_, _13115_, _03124_);
  or (_13193_, _13192_, _02650_);
  or (_13194_, _13193_, _13191_);
  nand (_13195_, _13136_, _02650_);
  and (_13196_, _13195_, _13194_);
  nor (_13197_, _13196_, _03121_);
  and (_13198_, _08807_, _04615_);
  nor (_13199_, _13198_, _13103_);
  and (_13200_, _13199_, _03121_);
  nor (_13201_, _13200_, _13197_);
  or (_13202_, _13201_, _27789_);
  or (_13203_, _27788_, \oc8051_golden_model_1.SCON [3]);
  and (_13204_, _13203_, _27053_);
  and (_28889_, _13204_, _13202_);
  not (_13205_, \oc8051_golden_model_1.SCON [4]);
  nor (_13206_, _04615_, _13205_);
  and (_13207_, _04615_, _05974_);
  nor (_13208_, _13207_, _13206_);
  and (_13209_, _13208_, _02575_);
  nor (_13210_, _06755_, _04325_);
  nor (_13211_, _13210_, _13206_);
  and (_13212_, _13211_, _05949_);
  nor (_13213_, _05431_, _13205_);
  nor (_13214_, _13213_, _08889_);
  and (_13215_, _08869_, _05431_);
  nor (_13216_, _13215_, _13213_);
  or (_13217_, _13216_, _05168_);
  nor (_13218_, _13217_, _13214_);
  nor (_13219_, _08838_, _06755_);
  nor (_13220_, _13219_, _13206_);
  and (_13221_, _13220_, _02661_);
  and (_13222_, _04615_, \oc8051_golden_model_1.ACC [4]);
  nor (_13223_, _13222_, _13206_);
  nor (_13224_, _13223_, _05903_);
  nor (_13225_, _04505_, _13205_);
  or (_13226_, _13225_, _02661_);
  nor (_13227_, _13226_, _13224_);
  or (_13228_, _13227_, _06504_);
  nor (_13229_, _13228_, _13221_);
  nor (_13230_, _13211_, _03365_);
  nor (_13231_, _13216_, _03390_);
  nor (_13232_, _13231_, _13230_);
  nand (_13233_, _13232_, _03179_);
  or (_13234_, _13233_, _13229_);
  nand (_13235_, _13223_, _03168_);
  and (_13236_, _13235_, _13234_);
  and (_13237_, _13236_, _03177_);
  and (_13238_, _08880_, _05431_);
  nor (_13239_, _13238_, _13213_);
  nor (_13240_, _13239_, _03177_);
  or (_13241_, _13240_, _13237_);
  and (_13242_, _13241_, _05168_);
  nor (_13243_, _13242_, _13218_);
  nor (_13244_, _13243_, _03140_);
  nor (_13245_, _08908_, _06792_);
  nor (_13246_, _13245_, _13213_);
  nor (_13247_, _13246_, _03141_);
  nor (_13248_, _13247_, _05949_);
  not (_13249_, _13248_);
  nor (_13250_, _13249_, _13244_);
  nor (_13251_, _13250_, _13212_);
  nor (_13252_, _13251_, _05959_);
  and (_13253_, _04615_, _04012_);
  nor (_13254_, _13206_, _05963_);
  not (_13255_, _13254_);
  nor (_13256_, _13255_, _13253_);
  or (_13257_, _13256_, _02024_);
  nor (_13258_, _13257_, _13252_);
  nor (_13259_, _08967_, _06755_);
  nor (_13260_, _13259_, _13206_);
  nor (_13261_, _13260_, _03139_);
  or (_13262_, _13261_, _02575_);
  nor (_13263_, _13262_, _13258_);
  nor (_13264_, _13263_, _13209_);
  or (_13265_, _13264_, _02656_);
  and (_13266_, _08982_, _04615_);
  or (_13267_, _13266_, _13206_);
  or (_13268_, _13267_, _05305_);
  and (_13269_, _13268_, _03252_);
  and (_13270_, _13269_, _13265_);
  and (_13271_, _08830_, _04615_);
  nor (_13272_, _13271_, _13206_);
  nor (_13273_, _13272_, _03252_);
  nor (_13274_, _13273_, _13270_);
  nor (_13275_, _13274_, _02669_);
  nor (_13276_, _13206_, _09034_);
  not (_13277_, _13276_);
  nor (_13278_, _13208_, _05332_);
  and (_13279_, _13278_, _13277_);
  nor (_13280_, _13279_, _13275_);
  nor (_13281_, _13280_, _03243_);
  or (_13282_, _13276_, _03244_);
  nor (_13283_, _13282_, _13223_);
  or (_13284_, _13283_, _02654_);
  nor (_13285_, _13284_, _13281_);
  nor (_13286_, _08981_, _06755_);
  nor (_13287_, _13286_, _13206_);
  and (_13288_, _13287_, _02654_);
  nor (_13289_, _13288_, _13285_);
  and (_13290_, _13289_, _05883_);
  nor (_13291_, _08828_, _06755_);
  nor (_13292_, _13291_, _13206_);
  nor (_13293_, _13292_, _05883_);
  or (_13294_, _13293_, _13290_);
  and (_13295_, _13294_, _03124_);
  nor (_13296_, _13220_, _03124_);
  or (_13297_, _13296_, _02650_);
  or (_13298_, _13297_, _13295_);
  nand (_13299_, _13239_, _02650_);
  and (_13300_, _13299_, _13298_);
  nor (_13301_, _13300_, _03121_);
  and (_13302_, _09037_, _04615_);
  nor (_13303_, _13302_, _13206_);
  and (_13304_, _13303_, _03121_);
  nor (_13305_, _13304_, _13301_);
  or (_13306_, _13305_, _27789_);
  or (_13307_, _27788_, \oc8051_golden_model_1.SCON [4]);
  and (_13308_, _13307_, _27053_);
  and (_28892_, _13308_, _13306_);
  not (_13309_, \oc8051_golden_model_1.SCON [5]);
  nor (_13310_, _04615_, _13309_);
  and (_13311_, _04615_, _06036_);
  nor (_13312_, _13311_, _13310_);
  and (_13313_, _13312_, _02575_);
  nor (_13314_, _06755_, _04480_);
  nor (_13315_, _13314_, _13310_);
  and (_13316_, _13315_, _05949_);
  nor (_13317_, _05431_, _13309_);
  nor (_13318_, _13317_, _09107_);
  and (_13319_, _09072_, _05431_);
  nor (_13320_, _13319_, _13317_);
  or (_13321_, _13320_, _05168_);
  nor (_13322_, _13321_, _13318_);
  nor (_13323_, _09087_, _06755_);
  nor (_13324_, _13323_, _13310_);
  and (_13325_, _13324_, _02661_);
  and (_13326_, _04615_, \oc8051_golden_model_1.ACC [5]);
  nor (_13327_, _13326_, _13310_);
  nor (_13328_, _13327_, _05903_);
  nor (_13329_, _04505_, _13309_);
  or (_13330_, _13329_, _02661_);
  nor (_13331_, _13330_, _13328_);
  or (_13332_, _13331_, _06504_);
  nor (_13333_, _13332_, _13325_);
  nor (_13334_, _13315_, _03365_);
  nor (_13335_, _13320_, _03390_);
  nor (_13336_, _13335_, _13334_);
  nand (_13337_, _13336_, _03179_);
  or (_13338_, _13337_, _13333_);
  nand (_13339_, _13327_, _03168_);
  and (_13340_, _13339_, _13338_);
  and (_13341_, _13340_, _03177_);
  and (_13342_, _09099_, _05431_);
  nor (_13343_, _13342_, _13317_);
  nor (_13344_, _13343_, _03177_);
  or (_13345_, _13344_, _13341_);
  and (_13346_, _13345_, _05168_);
  nor (_13347_, _13346_, _13322_);
  nor (_13348_, _13347_, _03140_);
  nor (_13349_, _09059_, _06792_);
  nor (_13350_, _13349_, _13317_);
  nor (_13351_, _13350_, _03141_);
  nor (_13352_, _13351_, _05949_);
  not (_13353_, _13352_);
  nor (_13354_, _13353_, _13348_);
  nor (_13355_, _13354_, _13316_);
  nor (_13356_, _13355_, _05959_);
  and (_13357_, _04615_, _03904_);
  nor (_13358_, _13310_, _05963_);
  not (_13359_, _13358_);
  nor (_13360_, _13359_, _13357_);
  or (_13361_, _13360_, _02024_);
  nor (_13362_, _13361_, _13356_);
  nor (_13363_, _09180_, _06755_);
  nor (_13364_, _13363_, _13310_);
  nor (_13365_, _13364_, _03139_);
  or (_13366_, _13365_, _02575_);
  nor (_13367_, _13366_, _13362_);
  nor (_13368_, _13367_, _13313_);
  or (_13369_, _13368_, _02656_);
  and (_13370_, _09195_, _04615_);
  or (_13371_, _13370_, _13310_);
  or (_13372_, _13371_, _05305_);
  and (_13373_, _13372_, _03252_);
  and (_13374_, _13373_, _13369_);
  and (_13375_, _09055_, _04615_);
  nor (_13376_, _13375_, _13310_);
  nor (_13377_, _13376_, _03252_);
  nor (_13378_, _13377_, _13374_);
  nor (_13379_, _13378_, _02669_);
  not (_13380_, _13310_);
  and (_13381_, _13380_, _04787_);
  not (_13382_, _13381_);
  nor (_13383_, _13312_, _05332_);
  and (_13384_, _13383_, _13382_);
  nor (_13385_, _13384_, _13379_);
  nor (_13386_, _13385_, _03243_);
  or (_13387_, _13381_, _03244_);
  nor (_13388_, _13387_, _13327_);
  or (_13389_, _13388_, _02654_);
  nor (_13390_, _13389_, _13386_);
  nor (_13391_, _09194_, _06755_);
  nor (_13392_, _13391_, _13310_);
  and (_13393_, _13392_, _02654_);
  nor (_13394_, _13393_, _13390_);
  and (_13395_, _13394_, _05883_);
  nor (_13396_, _09054_, _06755_);
  nor (_13397_, _13396_, _13310_);
  nor (_13398_, _13397_, _05883_);
  or (_13399_, _13398_, _13395_);
  and (_13400_, _13399_, _03124_);
  nor (_13401_, _13324_, _03124_);
  or (_13402_, _13401_, _02650_);
  or (_13403_, _13402_, _13400_);
  nand (_13404_, _13343_, _02650_);
  and (_13405_, _13404_, _13403_);
  nor (_13406_, _13405_, _03121_);
  and (_13407_, _09248_, _04615_);
  nor (_13408_, _13407_, _13310_);
  and (_13409_, _13408_, _03121_);
  nor (_13410_, _13409_, _13406_);
  or (_13411_, _13410_, _27789_);
  or (_13412_, _27788_, \oc8051_golden_model_1.SCON [5]);
  and (_13413_, _13412_, _27053_);
  and (_28893_, _13413_, _13411_);
  not (_13414_, \oc8051_golden_model_1.SCON [6]);
  nor (_13415_, _04615_, _13414_);
  and (_13416_, _04615_, _03960_);
  or (_13417_, _13416_, _13415_);
  and (_13418_, _13417_, _05959_);
  nor (_13419_, _05431_, _13414_);
  not (_13420_, _13419_);
  and (_13421_, _13420_, _09320_);
  and (_13422_, _09305_, _05431_);
  nor (_13423_, _13422_, _13419_);
  or (_13424_, _13423_, _05168_);
  nor (_13425_, _13424_, _13421_);
  nor (_13426_, _09301_, _06755_);
  nor (_13427_, _13426_, _13415_);
  and (_13428_, _13427_, _02661_);
  and (_13429_, _04615_, \oc8051_golden_model_1.ACC [6]);
  nor (_13430_, _13429_, _13415_);
  nor (_13431_, _13430_, _05903_);
  nor (_13432_, _04505_, _13414_);
  or (_13433_, _13432_, _02661_);
  nor (_13434_, _13433_, _13431_);
  or (_13435_, _13434_, _06504_);
  nor (_13436_, _13435_, _13428_);
  nor (_13437_, _06755_, _04373_);
  nor (_13438_, _13437_, _13415_);
  nor (_13439_, _13438_, _03365_);
  nor (_13440_, _13423_, _03390_);
  nor (_13441_, _13440_, _13439_);
  nand (_13442_, _13441_, _03179_);
  or (_13443_, _13442_, _13436_);
  nand (_13444_, _13430_, _03168_);
  and (_13445_, _13444_, _13443_);
  and (_13446_, _13445_, _03177_);
  and (_13447_, _09286_, _05431_);
  nor (_13448_, _13447_, _13419_);
  nor (_13449_, _13448_, _03177_);
  or (_13450_, _13449_, _13446_);
  and (_13451_, _13450_, _05168_);
  nor (_13452_, _13451_, _13425_);
  nor (_13453_, _13452_, _03140_);
  nor (_13454_, _09272_, _06792_);
  nor (_13455_, _13454_, _13419_);
  nor (_13456_, _13455_, _03141_);
  nor (_13457_, _13456_, _05949_);
  not (_13458_, _13457_);
  nor (_13459_, _13458_, _13453_);
  and (_13460_, _13438_, _05949_);
  or (_13461_, _13460_, _05959_);
  nor (_13462_, _13461_, _13459_);
  or (_13463_, _13462_, _13418_);
  and (_13464_, _13463_, _03139_);
  and (_13465_, _09388_, _04615_);
  nor (_13466_, _13465_, _13415_);
  nor (_13467_, _13466_, _03139_);
  or (_13468_, _13467_, _06549_);
  or (_13469_, _13468_, _13464_);
  and (_13470_, _09404_, _04615_);
  or (_13471_, _13415_, _05305_);
  or (_13472_, _13471_, _13470_);
  and (_13473_, _04615_, _09395_);
  nor (_13474_, _13473_, _13415_);
  and (_13475_, _13474_, _02575_);
  nor (_13476_, _13475_, _03251_);
  and (_13477_, _13476_, _13472_);
  and (_13478_, _13477_, _13469_);
  and (_13479_, _09268_, _04615_);
  nor (_13480_, _13479_, _13415_);
  nor (_13481_, _13480_, _03252_);
  nor (_13482_, _13481_, _13478_);
  nor (_13483_, _13482_, _02669_);
  nor (_13484_, _13415_, _06119_);
  not (_13485_, _13484_);
  nor (_13486_, _13474_, _05332_);
  and (_13487_, _13486_, _13485_);
  nor (_13488_, _13487_, _13483_);
  nor (_13489_, _13488_, _03243_);
  or (_13490_, _13484_, _03244_);
  nor (_13491_, _13490_, _13430_);
  or (_13492_, _13491_, _02654_);
  nor (_13493_, _13492_, _13489_);
  nor (_13494_, _09403_, _06755_);
  nor (_13495_, _13494_, _13415_);
  and (_13496_, _13495_, _02654_);
  nor (_13497_, _13496_, _13493_);
  and (_13498_, _13497_, _05883_);
  nor (_13499_, _09267_, _06755_);
  nor (_13500_, _13499_, _13415_);
  nor (_13501_, _13500_, _05883_);
  or (_13502_, _13501_, _13498_);
  and (_13503_, _13502_, _03124_);
  nor (_13504_, _13427_, _03124_);
  or (_13505_, _13504_, _02650_);
  or (_13506_, _13505_, _13503_);
  nand (_13507_, _13448_, _02650_);
  and (_13508_, _13507_, _13506_);
  nor (_13509_, _13508_, _03121_);
  and (_13510_, _09456_, _04615_);
  nor (_13511_, _13510_, _13415_);
  and (_13512_, _13511_, _03121_);
  nor (_13513_, _13512_, _13509_);
  or (_13514_, _13513_, _27789_);
  or (_13515_, _27788_, \oc8051_golden_model_1.SCON [6]);
  and (_13516_, _13515_, _27053_);
  and (_28894_, _13516_, _13514_);
  nor (_13517_, _04879_, _03417_);
  nor (_13518_, _08109_, _06608_);
  nor (_13519_, _13518_, _13517_);
  nor (_13520_, _13519_, _05883_);
  and (_13521_, _04879_, \oc8051_golden_model_1.ACC [0]);
  nor (_13522_, _13521_, _13517_);
  nor (_13523_, _13522_, _05903_);
  nor (_13524_, _04505_, _03417_);
  or (_13525_, _13524_, _13523_);
  and (_13526_, _13525_, _02662_);
  nor (_13527_, _04888_, _06608_);
  nor (_13528_, _13527_, _13517_);
  nor (_13529_, _13528_, _02662_);
  or (_13530_, _13529_, _13526_);
  and (_13531_, _13530_, _03365_);
  or (_13532_, _13531_, _03418_);
  and (_13533_, _13532_, _03179_);
  nor (_13534_, _13522_, _03179_);
  or (_13535_, _13534_, _13533_);
  and (_13536_, _13535_, _03430_);
  nor (_13537_, _07263_, _05949_);
  not (_13538_, _13537_);
  nor (_13539_, _13538_, _13536_);
  or (_13540_, _06608_, _04485_);
  nor (_13541_, _13517_, _06673_);
  and (_13542_, _13541_, _13540_);
  nor (_13543_, _13542_, _13539_);
  nor (_13544_, _13543_, _05959_);
  nor (_13545_, _13517_, _05963_);
  or (_13546_, _06608_, _04270_);
  and (_13547_, _13546_, _13545_);
  nor (_13548_, _13547_, _13544_);
  nor (_13549_, _13548_, _02024_);
  or (_13550_, _08093_, _06608_);
  nor (_13551_, _13517_, _03139_);
  and (_13552_, _13551_, _13550_);
  or (_13553_, _13552_, _02575_);
  nor (_13554_, _13553_, _13549_);
  and (_13555_, _04879_, _05996_);
  nor (_13556_, _13555_, _13517_);
  nand (_13557_, _13556_, _05305_);
  and (_13558_, _13557_, _06549_);
  nor (_13559_, _13558_, _13554_);
  and (_13560_, _07968_, _04879_);
  nor (_13561_, _13560_, _13517_);
  and (_13562_, _13561_, _02656_);
  nor (_13563_, _13562_, _13559_);
  and (_13564_, _13563_, _03252_);
  and (_13565_, _08110_, _04879_);
  nor (_13566_, _13565_, _13517_);
  nor (_13567_, _13566_, _03252_);
  or (_13568_, _13567_, _13564_);
  and (_13569_, _13568_, _05332_);
  nor (_13570_, _13556_, _05332_);
  not (_13571_, _13570_);
  nor (_13572_, _13571_, _13527_);
  nor (_13573_, _13572_, _13569_);
  nor (_13574_, _13573_, _03243_);
  and (_13575_, _08108_, _04879_);
  or (_13576_, _13575_, _13517_);
  and (_13577_, _13576_, _03243_);
  or (_13578_, _13577_, _13574_);
  and (_13579_, _13578_, _05357_);
  nor (_13580_, _07967_, _06718_);
  nor (_13581_, _13580_, _13517_);
  nor (_13582_, _13581_, _05357_);
  or (_13583_, _13582_, _13579_);
  and (_13584_, _13583_, _05883_);
  or (_13585_, _13584_, _11672_);
  nor (_13586_, _13585_, _13520_);
  and (_13587_, _13528_, _11672_);
  nor (_13588_, _13587_, _13586_);
  and (_13589_, _13588_, _27788_);
  nor (_13590_, _27788_, _03417_);
  or (_13591_, _13590_, rst);
  or (_28896_, _13591_, _13589_);
  nor (_13592_, _04879_, _03565_);
  and (_13593_, _08209_, _04564_);
  nor (_13594_, _13593_, _13592_);
  nor (_13595_, _13594_, _03513_);
  and (_13596_, _03109_, \oc8051_golden_model_1.SP [1]);
  nor (_13597_, _04879_, \oc8051_golden_model_1.SP [1]);
  not (_13598_, _13597_);
  or (_13599_, _08325_, _06718_);
  and (_13600_, _13599_, _03251_);
  and (_13601_, _13600_, _13598_);
  and (_13602_, _01967_, _03565_);
  not (_13603_, _01967_);
  and (_13604_, _04879_, \oc8051_golden_model_1.ACC [1]);
  or (_13605_, _13604_, _13592_);
  and (_13606_, _13605_, _04505_);
  nor (_13607_, _04505_, _03565_);
  or (_13608_, _13607_, _13606_);
  and (_13609_, _13608_, _01988_);
  nor (_13610_, _01988_, \oc8051_golden_model_1.SP [1]);
  or (_13611_, _13610_, _13609_);
  and (_13612_, _13611_, _02662_);
  nor (_13613_, _13597_, _13593_);
  and (_13614_, _13613_, _02661_);
  or (_13615_, _13614_, _13612_);
  and (_13616_, _13615_, _01995_);
  nor (_13617_, _01995_, \oc8051_golden_model_1.SP [1]);
  or (_13618_, _13617_, _03162_);
  or (_13619_, _13618_, _13616_);
  nand (_13620_, _03783_, _03162_);
  and (_13621_, _13620_, _13619_);
  and (_13622_, _13621_, _03179_);
  and (_13623_, _13605_, _03168_);
  or (_13624_, _13623_, _13622_);
  and (_13625_, _13624_, _03430_);
  or (_13626_, _13625_, _06666_);
  nor (_13627_, _13626_, _07409_);
  nor (_13628_, _06665_, _03565_);
  or (_13629_, _13628_, _05949_);
  nor (_13630_, _13629_, _13627_);
  nand (_13631_, _04564_, _03777_);
  nor (_13632_, _13597_, _06673_);
  and (_13633_, _13632_, _13631_);
  nor (_13634_, _13633_, _05959_);
  not (_13635_, _13634_);
  nor (_13636_, _13635_, _13630_);
  nor (_13637_, _13592_, _05963_);
  or (_13638_, _06608_, _04221_);
  and (_13639_, _13638_, _13637_);
  nor (_13640_, _13639_, _02024_);
  not (_13641_, _13640_);
  nor (_13642_, _13641_, _13636_);
  nor (_13643_, _13597_, _03139_);
  nand (_13644_, _08307_, _04879_);
  and (_13645_, _13644_, _13643_);
  nor (_13646_, _13645_, _13642_);
  nor (_13647_, _13646_, _02575_);
  and (_13648_, _04879_, _05984_);
  or (_13649_, _13648_, _13592_);
  and (_13650_, _13649_, _02575_);
  or (_13651_, _13650_, _13647_);
  and (_13652_, _13651_, _13603_);
  or (_13653_, _13652_, _13602_);
  and (_13654_, _13653_, _05305_);
  or (_13655_, _08185_, _06718_);
  and (_13656_, _13655_, _02656_);
  and (_13657_, _13656_, _13598_);
  nor (_13658_, _13657_, _13654_);
  nor (_13659_, _13658_, _03251_);
  nor (_13660_, _13659_, _13601_);
  nor (_13661_, _13660_, _02669_);
  or (_13662_, _08184_, _06718_);
  and (_13663_, _13662_, _02669_);
  and (_13664_, _13663_, _13598_);
  nor (_13665_, _13664_, _13661_);
  nor (_13666_, _13665_, _05339_);
  and (_13667_, _01965_, _03565_);
  nor (_13668_, _13592_, _06122_);
  nor (_13669_, _13668_, _03244_);
  and (_13670_, _13669_, _13605_);
  or (_13671_, _13670_, _13667_);
  nor (_13672_, _13671_, _13666_);
  nor (_13673_, _13672_, _03241_);
  and (_13674_, _08324_, _04879_);
  nor (_13675_, _13674_, _05883_);
  and (_13676_, _04564_, _03016_);
  nand (_13677_, _13676_, _04835_);
  and (_13678_, _13677_, _02654_);
  nor (_13679_, _13678_, _13675_);
  or (_13680_, _13679_, _13597_);
  and (_13681_, _13680_, _06612_);
  not (_13682_, _13681_);
  nor (_13683_, _13682_, _13673_);
  nor (_13684_, _13683_, _13596_);
  nor (_13685_, _03108_, _01936_);
  not (_13686_, _13685_);
  nor (_13687_, _13686_, _13684_);
  nor (_13688_, _13685_, _03565_);
  nor (_13689_, _13688_, _03123_);
  not (_13690_, _13689_);
  nor (_13691_, _13690_, _13687_);
  and (_13692_, _13613_, _03123_);
  nor (_13693_, _13692_, _06742_);
  not (_13694_, _13693_);
  nor (_13695_, _13694_, _13691_);
  nor (_13696_, _06741_, _03565_);
  nor (_13697_, _13696_, _03121_);
  not (_13698_, _13697_);
  nor (_13699_, _13698_, _13695_);
  nor (_13700_, _13699_, _13595_);
  nor (_13701_, _13700_, _27789_);
  nor (_13702_, _27788_, _03565_);
  or (_13703_, _13702_, rst);
  or (_28897_, _13703_, _13701_);
  and (_13704_, _07762_, _01936_);
  nor (_13705_, _04879_, _03111_);
  and (_13706_, _08387_, _04564_);
  nor (_13707_, _13706_, _13705_);
  nor (_13708_, _13707_, _03252_);
  and (_13709_, _09800_, _01967_);
  or (_13710_, _06608_, _03644_);
  nor (_13711_, _13705_, _06673_);
  and (_13712_, _13711_, _13710_);
  nor (_13713_, _09800_, _02000_);
  nor (_13714_, _04505_, _03111_);
  and (_13715_, _04879_, \oc8051_golden_model_1.ACC [2]);
  nor (_13716_, _13715_, _13705_);
  nor (_13717_, _13716_, _05903_);
  or (_13718_, _13717_, _13714_);
  and (_13719_, _13718_, _01988_);
  nor (_13720_, _09800_, _01988_);
  nor (_13721_, _13720_, _13719_);
  nor (_13722_, _13721_, _02661_);
  nor (_13723_, _08420_, _06608_);
  nor (_13724_, _13723_, _13705_);
  nor (_13725_, _13724_, _02662_);
  or (_13726_, _13725_, _13722_);
  and (_13727_, _13726_, _01995_);
  nor (_13728_, _09800_, _01995_);
  or (_13729_, _13728_, _03162_);
  or (_13730_, _13729_, _13727_);
  nand (_13731_, _03162_, _03115_);
  and (_13732_, _13731_, _13730_);
  and (_13733_, _13732_, _03179_);
  nor (_13734_, _13716_, _03179_);
  or (_13735_, _13734_, _13733_);
  and (_13736_, _13735_, _03430_);
  or (_13737_, _13736_, _07698_);
  and (_13738_, _13737_, _02000_);
  or (_13739_, _13738_, _13713_);
  and (_13740_, _13739_, _07791_);
  and (_13741_, _07762_, _02025_);
  nor (_13742_, _13741_, _05949_);
  not (_13743_, _13742_);
  nor (_13744_, _13743_, _13740_);
  nor (_13745_, _13744_, _13712_);
  nor (_13746_, _13745_, _05959_);
  nor (_13747_, _13705_, _05963_);
  or (_13748_, _06608_, _04168_);
  and (_13749_, _13748_, _13747_);
  or (_13750_, _13749_, _02024_);
  nor (_13751_, _13750_, _13746_);
  nor (_13752_, _08522_, _06718_);
  nor (_13753_, _13752_, _13705_);
  nor (_13754_, _13753_, _03139_);
  or (_13755_, _13754_, _02575_);
  or (_13756_, _13755_, _13751_);
  and (_13757_, _04879_, _06009_);
  nor (_13758_, _13757_, _13705_);
  nand (_13759_, _13758_, _02575_);
  and (_13760_, _13759_, _13756_);
  nor (_13761_, _13760_, _01967_);
  nor (_13762_, _13761_, _13709_);
  and (_13763_, _13762_, _05305_);
  and (_13764_, _08537_, _04879_);
  nor (_13765_, _13764_, _13705_);
  nor (_13766_, _13765_, _05305_);
  or (_13767_, _13766_, _13763_);
  and (_13768_, _13767_, _03252_);
  nor (_13769_, _13768_, _13708_);
  nor (_13770_, _13769_, _02669_);
  nor (_13771_, _13705_, _06121_);
  not (_13772_, _13771_);
  nor (_13773_, _13758_, _05332_);
  and (_13774_, _13773_, _13772_);
  nor (_13775_, _13774_, _13770_);
  nor (_13776_, _13775_, _05339_);
  and (_13777_, _07762_, _01965_);
  or (_13778_, _13771_, _03244_);
  nor (_13779_, _13778_, _13716_);
  or (_13780_, _13779_, _13777_);
  or (_13781_, _13780_, _02654_);
  nor (_13782_, _13781_, _13776_);
  nor (_13783_, _08536_, _06718_);
  nor (_13784_, _13783_, _13705_);
  and (_13785_, _13784_, _02654_);
  nor (_13786_, _13785_, _13782_);
  and (_13787_, _13786_, _05883_);
  nor (_13788_, _08386_, _06718_);
  nor (_13789_, _13788_, _13705_);
  nor (_13790_, _13789_, _05883_);
  or (_13791_, _13790_, _13787_);
  and (_13792_, _13791_, _06612_);
  and (_13793_, _09800_, _03109_);
  or (_13794_, _13793_, _13792_);
  and (_13795_, _13794_, _05408_);
  or (_13796_, _13795_, _13704_);
  and (_13797_, _13796_, _03126_);
  and (_13798_, _09800_, _03108_);
  or (_13799_, _13798_, _03123_);
  nor (_13800_, _13799_, _13797_);
  and (_13801_, _13724_, _03123_);
  or (_13802_, _13801_, _06742_);
  nor (_13803_, _13802_, _13800_);
  nor (_13804_, _09800_, _06741_);
  nor (_13805_, _13804_, _03121_);
  not (_13806_, _13805_);
  nor (_13807_, _13806_, _13803_);
  and (_13808_, _08596_, _04879_);
  nor (_13809_, _13808_, _13705_);
  and (_13810_, _13809_, _03121_);
  nor (_13811_, _13810_, _13807_);
  and (_13812_, _13811_, _27788_);
  nor (_13813_, _27788_, _03111_);
  or (_13814_, _13813_, rst);
  or (_28898_, _13814_, _13812_);
  nor (_13815_, _04879_, _03800_);
  and (_13816_, _08807_, _04564_);
  nor (_13817_, _13816_, _13815_);
  nor (_13818_, _13817_, _03513_);
  nor (_13819_, _08646_, _06608_);
  nor (_13820_, _13819_, _13815_);
  nor (_13821_, _13820_, _03124_);
  and (_13822_, _08618_, _04564_);
  nor (_13823_, _13822_, _13815_);
  nor (_13824_, _13823_, _03252_);
  and (_13825_, _09618_, _01967_);
  and (_13826_, _04879_, \oc8051_golden_model_1.ACC [3]);
  nor (_13827_, _13826_, _13815_);
  nor (_13828_, _13827_, _05903_);
  nor (_13829_, _04505_, _03800_);
  or (_13830_, _13829_, _04504_);
  nor (_13831_, _13830_, _13828_);
  nor (_13832_, _07765_, _01988_);
  nor (_13833_, _13832_, _13831_);
  and (_13834_, _13833_, _02662_);
  nor (_13835_, _13820_, _02662_);
  or (_13836_, _13835_, _13834_);
  and (_13837_, _13836_, _01995_);
  nor (_13838_, _09618_, _01995_);
  or (_13839_, _13838_, _03162_);
  or (_13840_, _13839_, _13837_);
  nand (_13841_, _03805_, _03162_);
  and (_13842_, _13841_, _13840_);
  and (_13843_, _13842_, _03179_);
  nor (_13844_, _13827_, _03179_);
  or (_13845_, _13844_, _13843_);
  and (_13846_, _13845_, _03430_);
  or (_13847_, _13846_, _06666_);
  nor (_13848_, _13847_, _07594_);
  nor (_13849_, _07765_, _06665_);
  or (_13850_, _13849_, _05949_);
  nor (_13851_, _13850_, _13848_);
  nor (_13852_, _06608_, _03859_);
  nor (_13853_, _13852_, _13815_);
  nor (_13854_, _13853_, _06673_);
  nor (_13855_, _13854_, _05959_);
  not (_13856_, _13855_);
  nor (_13857_, _13856_, _13851_);
  nor (_13858_, _13815_, _05963_);
  or (_13859_, _06608_, _04118_);
  and (_13860_, _13859_, _13858_);
  or (_13861_, _13860_, _02024_);
  nor (_13862_, _13861_, _13857_);
  nor (_13863_, _08744_, _06718_);
  nor (_13864_, _13863_, _13815_);
  nor (_13865_, _13864_, _03139_);
  or (_13866_, _13865_, _02575_);
  or (_13867_, _13866_, _13862_);
  and (_13868_, _04879_, _05986_);
  nor (_13869_, _13868_, _13815_);
  nand (_13870_, _13869_, _02575_);
  and (_13871_, _13870_, _13867_);
  nor (_13872_, _13871_, _01967_);
  nor (_13873_, _13872_, _13825_);
  and (_13874_, _13873_, _05305_);
  and (_13875_, _08622_, _04879_);
  nor (_13876_, _13875_, _13815_);
  nor (_13877_, _13876_, _05305_);
  or (_13878_, _13877_, _13874_);
  and (_13879_, _13878_, _03252_);
  nor (_13880_, _13879_, _13824_);
  nor (_13881_, _13880_, _02669_);
  not (_13882_, _13815_);
  and (_13883_, _13882_, _04649_);
  or (_13884_, _13883_, _05332_);
  nor (_13885_, _13884_, _13869_);
  nor (_13886_, _13885_, _13881_);
  nor (_13887_, _13886_, _05339_);
  and (_13888_, _07765_, _01965_);
  nor (_13889_, _13888_, _02654_);
  or (_13890_, _13827_, _03244_);
  or (_13891_, _13890_, _13883_);
  nand (_13892_, _13891_, _13889_);
  nor (_13893_, _13892_, _13887_);
  nor (_13894_, _08621_, _06718_);
  nor (_13895_, _13894_, _13815_);
  and (_13896_, _13895_, _02654_);
  nor (_13897_, _13896_, _13893_);
  and (_13898_, _13897_, _05883_);
  nor (_13899_, _08617_, _06718_);
  nor (_13900_, _13899_, _13815_);
  nor (_13901_, _13900_, _05883_);
  or (_13902_, _13901_, _13898_);
  and (_13903_, _13902_, _06612_);
  nor (_13904_, _03802_, _03800_);
  nor (_13905_, _13904_, _03803_);
  nor (_13906_, _13905_, _06612_);
  or (_13907_, _13906_, _01936_);
  or (_13908_, _13907_, _13903_);
  nand (_13909_, _09618_, _01936_);
  and (_13910_, _13909_, _13908_);
  and (_13911_, _13910_, _03126_);
  nor (_13912_, _13905_, _03126_);
  or (_13913_, _13912_, _13911_);
  and (_13914_, _13913_, _03124_);
  or (_13915_, _13914_, _06742_);
  nor (_13916_, _13915_, _13821_);
  nor (_13917_, _07765_, _06741_);
  nor (_13918_, _13917_, _03121_);
  not (_13919_, _13918_);
  nor (_13920_, _13919_, _13916_);
  nor (_13921_, _13920_, _13818_);
  nand (_13922_, _13921_, _27788_);
  or (_13923_, _27788_, \oc8051_golden_model_1.SP [3]);
  and (_13924_, _13923_, _27053_);
  and (_28899_, _13924_, _13922_);
  nor (_13925_, _04879_, _06642_);
  and (_13926_, _09037_, _04564_);
  nor (_13927_, _13926_, _13925_);
  nor (_13928_, _13927_, _03513_);
  nor (_13929_, _08838_, _06608_);
  nor (_13930_, _13929_, _13925_);
  nor (_13931_, _13930_, _03124_);
  and (_13932_, _08830_, _04564_);
  nor (_13933_, _13932_, _13925_);
  nor (_13934_, _13933_, _03252_);
  nor (_13935_, _04505_, _06642_);
  and (_13936_, _04879_, \oc8051_golden_model_1.ACC [4]);
  nor (_13937_, _13936_, _13925_);
  nor (_13938_, _13937_, _05903_);
  or (_13939_, _13938_, _13935_);
  and (_13940_, _13939_, _01988_);
  nor (_13941_, _06623_, \oc8051_golden_model_1.SP [4]);
  nor (_13942_, _13941_, _06624_);
  and (_13943_, _13942_, _04504_);
  nor (_13944_, _13943_, _13940_);
  nor (_13945_, _13944_, _02661_);
  nor (_13946_, _13930_, _02662_);
  or (_13947_, _13946_, _13945_);
  and (_13948_, _13947_, _01995_);
  and (_13949_, _13942_, _07558_);
  or (_13950_, _13949_, _13948_);
  and (_13951_, _13950_, _03365_);
  and (_13952_, _06643_, _03417_);
  nor (_13953_, _03804_, _06642_);
  nor (_13954_, _13953_, _13952_);
  nor (_13955_, _13954_, _03365_);
  or (_13956_, _13955_, _13951_);
  and (_13957_, _13956_, _03179_);
  nor (_13958_, _13937_, _03179_);
  or (_13959_, _13958_, _13957_);
  and (_13960_, _13959_, _03430_);
  and (_13961_, _06656_, _06642_);
  nor (_13962_, _13961_, _06657_);
  and (_13963_, _13962_, _03187_);
  nor (_13964_, _13963_, _06666_);
  not (_13965_, _13964_);
  nor (_13966_, _13965_, _13960_);
  nor (_13967_, _13942_, _06665_);
  or (_13968_, _13967_, _05949_);
  nor (_13969_, _13968_, _13966_);
  nor (_13970_, _06608_, _04325_);
  nor (_13971_, _13970_, _13925_);
  nor (_13972_, _13971_, _06673_);
  nor (_13973_, _13972_, _05959_);
  not (_13974_, _13973_);
  nor (_13975_, _13974_, _13969_);
  nor (_13976_, _13925_, _05963_);
  or (_13977_, _06608_, _04014_);
  and (_13978_, _13977_, _13976_);
  nor (_13979_, _13978_, _02024_);
  not (_13980_, _13979_);
  nor (_13981_, _13980_, _13975_);
  nor (_13982_, _08967_, _06608_);
  nor (_13983_, _13982_, _13925_);
  nor (_13984_, _13983_, _03139_);
  or (_13985_, _13984_, _13981_);
  and (_13986_, _13985_, _05245_);
  and (_13987_, _04879_, _05974_);
  nor (_13988_, _13987_, _13925_);
  nor (_13989_, _13988_, _05245_);
  or (_13990_, _13989_, _13986_);
  and (_13991_, _13990_, _13603_);
  and (_13992_, _13942_, _01967_);
  or (_13993_, _13992_, _13991_);
  and (_13994_, _13993_, _05305_);
  and (_13995_, _08982_, _04879_);
  nor (_13996_, _13995_, _13925_);
  nor (_13997_, _13996_, _05305_);
  or (_13998_, _13997_, _13994_);
  and (_13999_, _13998_, _03252_);
  nor (_14000_, _13999_, _13934_);
  nor (_14001_, _14000_, _02669_);
  nor (_14002_, _13925_, _09034_);
  not (_14003_, _14002_);
  nor (_14004_, _13988_, _05332_);
  and (_14005_, _14004_, _14003_);
  nor (_14006_, _14005_, _14001_);
  nor (_14007_, _14006_, _05339_);
  and (_14008_, _13942_, _01965_);
  or (_14009_, _14002_, _03244_);
  nor (_14010_, _14009_, _13937_);
  or (_14011_, _14010_, _14008_);
  or (_14012_, _14011_, _02654_);
  nor (_14013_, _14012_, _14007_);
  nor (_14014_, _08981_, _06718_);
  nor (_14015_, _14014_, _13925_);
  and (_14016_, _14015_, _02654_);
  nor (_14017_, _14016_, _14013_);
  and (_14018_, _14017_, _05883_);
  nor (_14019_, _08828_, _06718_);
  nor (_14020_, _14019_, _13925_);
  nor (_14021_, _14020_, _05883_);
  or (_14022_, _14021_, _14018_);
  and (_14023_, _14022_, _06612_);
  nor (_14024_, _03803_, _06642_);
  nor (_14025_, _14024_, _06643_);
  nor (_14026_, _14025_, _06612_);
  or (_14027_, _14026_, _01936_);
  or (_14028_, _14027_, _14023_);
  or (_14029_, _13942_, _05408_);
  and (_14030_, _14029_, _14028_);
  and (_14031_, _14030_, _03126_);
  nor (_14032_, _14025_, _03126_);
  or (_14033_, _14032_, _14031_);
  and (_14034_, _14033_, _03124_);
  or (_14035_, _14034_, _06742_);
  nor (_14036_, _14035_, _13931_);
  nor (_14037_, _13942_, _06741_);
  nor (_14038_, _14037_, _03121_);
  not (_14039_, _14038_);
  nor (_14040_, _14039_, _14036_);
  nor (_14041_, _14040_, _13928_);
  nand (_14042_, _14041_, _27788_);
  or (_14043_, _27788_, \oc8051_golden_model_1.SP [4]);
  and (_14044_, _14043_, _27053_);
  and (_28900_, _14044_, _14042_);
  nor (_14045_, _04879_, _06641_);
  and (_14046_, _09248_, _04564_);
  nor (_14047_, _14046_, _14045_);
  nor (_14048_, _14047_, _03513_);
  nor (_14049_, _09087_, _06608_);
  nor (_14050_, _14049_, _14045_);
  nor (_14051_, _14050_, _03124_);
  and (_14052_, _09055_, _04564_);
  nor (_14053_, _14052_, _14045_);
  nor (_14054_, _14053_, _03252_);
  and (_14055_, _14050_, _02661_);
  and (_14056_, _04879_, \oc8051_golden_model_1.ACC [5]);
  nor (_14057_, _14056_, _14045_);
  nor (_14058_, _14057_, _05903_);
  nor (_14059_, _04505_, _06641_);
  or (_14060_, _14059_, _04504_);
  nor (_14061_, _14060_, _14058_);
  nor (_14062_, _06624_, \oc8051_golden_model_1.SP [5]);
  nor (_14063_, _14062_, _06625_);
  nor (_14064_, _14063_, _01988_);
  nor (_14065_, _14064_, _14061_);
  nor (_14066_, _14065_, _02661_);
  or (_14067_, _14066_, _14055_);
  nor (_14068_, _14067_, _07558_);
  not (_14069_, _14063_);
  nor (_14070_, _14069_, _01995_);
  or (_14071_, _14070_, _03162_);
  nor (_14072_, _14071_, _14068_);
  and (_14073_, _06644_, _03417_);
  nor (_14074_, _13952_, _06641_);
  nor (_14075_, _14074_, _14073_);
  and (_14076_, _14075_, _03162_);
  nor (_14077_, _14076_, _14072_);
  and (_14078_, _14077_, _03179_);
  nor (_14079_, _14057_, _03179_);
  or (_14080_, _14079_, _14078_);
  and (_14081_, _14080_, _03430_);
  nor (_14082_, _06657_, \oc8051_golden_model_1.SP [5]);
  nor (_14083_, _14082_, _06658_);
  and (_14084_, _14083_, _03187_);
  nor (_14085_, _14084_, _06666_);
  not (_14086_, _14085_);
  nor (_14087_, _14086_, _14081_);
  nor (_14088_, _14063_, _06665_);
  or (_14089_, _14088_, _05949_);
  nor (_14090_, _14089_, _14087_);
  nor (_14091_, _06608_, _04480_);
  nor (_14092_, _14091_, _14045_);
  nor (_14093_, _14092_, _06673_);
  nor (_14094_, _14093_, _05959_);
  not (_14095_, _14094_);
  nor (_14096_, _14095_, _14090_);
  nor (_14097_, _14045_, _05963_);
  or (_14098_, _06718_, _03906_);
  and (_14099_, _14098_, _14097_);
  or (_14100_, _14099_, _02024_);
  nor (_14101_, _14100_, _14096_);
  nor (_14102_, _09180_, _06718_);
  nor (_14103_, _14102_, _14045_);
  nor (_14104_, _14103_, _03139_);
  or (_14105_, _14104_, _02575_);
  or (_14106_, _14105_, _14101_);
  and (_14107_, _04879_, _06036_);
  nor (_14108_, _14107_, _14045_);
  nand (_14109_, _14108_, _02575_);
  and (_14110_, _14109_, _14106_);
  nor (_14111_, _14110_, _01967_);
  and (_14112_, _14069_, _01967_);
  nor (_14113_, _14112_, _14111_);
  and (_14114_, _14113_, _05305_);
  and (_14115_, _09195_, _04879_);
  nor (_14116_, _14115_, _14045_);
  nor (_14117_, _14116_, _05305_);
  or (_14118_, _14117_, _14114_);
  and (_14119_, _14118_, _03252_);
  nor (_14120_, _14119_, _14054_);
  nor (_14121_, _14120_, _02669_);
  not (_14122_, _14045_);
  and (_14123_, _14122_, _04787_);
  or (_14124_, _14123_, _05332_);
  nor (_14125_, _14124_, _14108_);
  nor (_14126_, _14125_, _14121_);
  nor (_14127_, _14126_, _05339_);
  and (_14128_, _14063_, _01965_);
  nor (_14129_, _14128_, _02654_);
  or (_14130_, _14057_, _03244_);
  or (_14131_, _14130_, _14123_);
  nand (_14132_, _14131_, _14129_);
  nor (_14133_, _14132_, _14127_);
  nor (_14134_, _09194_, _06718_);
  nor (_14135_, _14134_, _14045_);
  and (_14136_, _14135_, _02654_);
  nor (_14137_, _14136_, _14133_);
  and (_14138_, _14137_, _05883_);
  nor (_14139_, _09054_, _06718_);
  nor (_14140_, _14139_, _14045_);
  nor (_14141_, _14140_, _05883_);
  or (_14142_, _14141_, _14138_);
  and (_14143_, _14142_, _06612_);
  nor (_14144_, _06643_, _06641_);
  nor (_14145_, _14144_, _06644_);
  nor (_14146_, _14145_, _06612_);
  or (_14147_, _14146_, _01936_);
  or (_14148_, _14147_, _14143_);
  nand (_14149_, _14069_, _01936_);
  and (_14150_, _14149_, _14148_);
  and (_14151_, _14150_, _03126_);
  nor (_14152_, _14145_, _03126_);
  or (_14153_, _14152_, _14151_);
  and (_14154_, _14153_, _03124_);
  or (_14155_, _14154_, _06742_);
  nor (_14156_, _14155_, _14051_);
  nor (_14157_, _14063_, _06741_);
  nor (_14158_, _14157_, _03121_);
  not (_14159_, _14158_);
  nor (_14160_, _14159_, _14156_);
  nor (_14161_, _14160_, _14048_);
  nand (_14162_, _14161_, _27788_);
  or (_14163_, _27788_, \oc8051_golden_model_1.SP [5]);
  and (_14164_, _14163_, _27053_);
  and (_28901_, _14164_, _14162_);
  nor (_14165_, _04879_, _06640_);
  and (_14166_, _09268_, _04564_);
  nor (_14167_, _14166_, _14165_);
  nor (_14168_, _14167_, _03252_);
  and (_14169_, _04879_, _03960_);
  or (_14170_, _14169_, _14165_);
  and (_14171_, _14170_, _05959_);
  nor (_14172_, _04505_, _06640_);
  and (_14173_, _04879_, \oc8051_golden_model_1.ACC [6]);
  nor (_14174_, _14173_, _14165_);
  nor (_14175_, _14174_, _05903_);
  or (_14176_, _14175_, _14172_);
  and (_14177_, _14176_, _01988_);
  nor (_14178_, _06625_, \oc8051_golden_model_1.SP [6]);
  nor (_14179_, _14178_, _06626_);
  not (_14180_, _14179_);
  nor (_14181_, _14180_, _01988_);
  nor (_14182_, _14181_, _14177_);
  nor (_14183_, _14182_, _02661_);
  nor (_14184_, _09301_, _06608_);
  nor (_14185_, _14184_, _14165_);
  nor (_14186_, _14185_, _02662_);
  or (_14187_, _14186_, _14183_);
  and (_14188_, _14187_, _01995_);
  nor (_14189_, _14180_, _01995_);
  or (_14190_, _14189_, _14188_);
  and (_14191_, _14190_, _03365_);
  nor (_14192_, _14073_, _06640_);
  nor (_14193_, _14192_, _06646_);
  nor (_14194_, _14193_, _03365_);
  or (_14195_, _14194_, _14191_);
  and (_14196_, _14195_, _03179_);
  nor (_14197_, _14174_, _03179_);
  or (_14198_, _14197_, _14196_);
  and (_14199_, _14198_, _03430_);
  nor (_14200_, _06658_, \oc8051_golden_model_1.SP [6]);
  nor (_14201_, _14200_, _06659_);
  and (_14202_, _14201_, _03187_);
  nor (_14203_, _14202_, _14199_);
  nor (_14204_, _14203_, _06666_);
  nor (_14205_, _14180_, _06665_);
  nor (_14206_, _14205_, _05949_);
  not (_14207_, _14206_);
  nor (_14208_, _14207_, _14204_);
  or (_14209_, _06608_, _04373_);
  nor (_14210_, _14165_, _06673_);
  and (_14211_, _14210_, _14209_);
  or (_14212_, _14211_, _05959_);
  nor (_14213_, _14212_, _14208_);
  or (_14214_, _14213_, _14171_);
  and (_14215_, _14214_, _03139_);
  and (_14216_, _09388_, _04564_);
  nor (_14217_, _14216_, _14165_);
  nor (_14218_, _14217_, _03139_);
  or (_14219_, _14218_, _02575_);
  or (_14220_, _14219_, _14215_);
  and (_14221_, _04879_, _09395_);
  nor (_14222_, _14221_, _14165_);
  nand (_14223_, _14222_, _02575_);
  and (_14224_, _14223_, _14220_);
  nor (_14225_, _14224_, _01967_);
  and (_14226_, _14180_, _01967_);
  nor (_14227_, _14226_, _14225_);
  and (_14228_, _14227_, _05305_);
  and (_14229_, _09404_, _04879_);
  nor (_14230_, _14229_, _14165_);
  nor (_14231_, _14230_, _05305_);
  or (_14232_, _14231_, _14228_);
  and (_14233_, _14232_, _03252_);
  nor (_14234_, _14233_, _14168_);
  nor (_14235_, _14234_, _02669_);
  nor (_14236_, _14165_, _06119_);
  not (_14237_, _14236_);
  nor (_14238_, _14222_, _05332_);
  and (_14239_, _14238_, _14237_);
  nor (_14240_, _14239_, _14235_);
  nor (_14241_, _14240_, _05339_);
  and (_14242_, _14179_, _01965_);
  or (_14243_, _14236_, _03244_);
  nor (_14244_, _14243_, _14174_);
  or (_14245_, _14244_, _14242_);
  or (_14246_, _14245_, _02654_);
  nor (_14247_, _14246_, _14241_);
  nor (_14248_, _09403_, _06718_);
  nor (_14249_, _14248_, _14165_);
  and (_14250_, _14249_, _02654_);
  nor (_14251_, _14250_, _14247_);
  and (_14252_, _14251_, _05883_);
  nor (_14253_, _09267_, _06718_);
  nor (_14254_, _14253_, _14165_);
  nor (_14255_, _14254_, _05883_);
  or (_14256_, _14255_, _14252_);
  and (_14257_, _14256_, _06612_);
  nor (_14258_, _06644_, _06640_);
  nor (_14259_, _14258_, _06645_);
  nor (_14260_, _14259_, _06612_);
  or (_14261_, _14260_, _01936_);
  or (_14262_, _14261_, _14257_);
  nand (_14263_, _14180_, _01936_);
  and (_14264_, _14263_, _14262_);
  nor (_14265_, _14264_, _03108_);
  and (_14266_, _14259_, _03108_);
  nor (_14267_, _14266_, _14265_);
  nor (_14268_, _14267_, _03123_);
  and (_14269_, _14185_, _03123_);
  nor (_14270_, _14269_, _06742_);
  not (_14271_, _14270_);
  nor (_14272_, _14271_, _14268_);
  nor (_14273_, _14180_, _06741_);
  nor (_14274_, _14273_, _03121_);
  not (_14275_, _14274_);
  nor (_14276_, _14275_, _14272_);
  and (_14277_, _09456_, _04879_);
  nor (_14278_, _14277_, _14165_);
  and (_14279_, _14278_, _03121_);
  nor (_14280_, _14279_, _14276_);
  or (_14281_, _14280_, _27789_);
  or (_14282_, _27788_, \oc8051_golden_model_1.SP [6]);
  and (_14283_, _14282_, _27053_);
  and (_28902_, _14283_, _14281_);
  not (_14284_, \oc8051_golden_model_1.TCON [0]);
  nor (_14285_, _04597_, _14284_);
  nor (_14286_, _04888_, _06476_);
  nor (_14287_, _14286_, _14285_);
  nor (_14288_, _14287_, _03513_);
  and (_14289_, _04597_, _05996_);
  nor (_14290_, _14289_, _14285_);
  nor (_14291_, _14290_, _05332_);
  not (_14292_, _14291_);
  nor (_14293_, _14292_, _14286_);
  and (_14294_, _04597_, _04268_);
  nor (_14295_, _14285_, _05963_);
  not (_14296_, _14295_);
  nor (_14297_, _14296_, _14294_);
  nor (_14298_, _05440_, _14284_);
  and (_14299_, _07997_, _05440_);
  nor (_14300_, _14299_, _14298_);
  nor (_14301_, _14300_, _03390_);
  and (_14302_, _14287_, _02661_);
  and (_14303_, _04597_, \oc8051_golden_model_1.ACC [0]);
  nor (_14304_, _14303_, _14285_);
  nor (_14305_, _14304_, _05903_);
  nor (_14306_, _04505_, _14284_);
  or (_14307_, _14306_, _02661_);
  nor (_14308_, _14307_, _14305_);
  or (_14309_, _14308_, _06504_);
  nor (_14310_, _14309_, _14302_);
  and (_14311_, _04597_, _03716_);
  nor (_14312_, _14311_, _14285_);
  nor (_14313_, _14312_, _03365_);
  or (_14314_, _14313_, _03168_);
  or (_14315_, _14314_, _14310_);
  nor (_14316_, _14315_, _14301_);
  and (_14317_, _14304_, _03168_);
  nor (_14318_, _14317_, _03176_);
  not (_14319_, _14318_);
  nor (_14320_, _14319_, _14316_);
  and (_14321_, _14285_, _03176_);
  or (_14322_, _14321_, _14320_);
  and (_14323_, _14322_, _05168_);
  nor (_14324_, _14287_, _05168_);
  or (_14325_, _14324_, _14323_);
  nor (_14326_, _14325_, _03140_);
  nor (_14327_, _08035_, _06529_);
  or (_14328_, _14298_, _03141_);
  nor (_14329_, _14328_, _14327_);
  or (_14330_, _14329_, _05949_);
  or (_14331_, _14330_, _14326_);
  or (_14332_, _14312_, _06673_);
  and (_14333_, _14332_, _05963_);
  and (_14334_, _14333_, _14331_);
  nor (_14335_, _14334_, _14297_);
  nor (_14336_, _14335_, _02024_);
  nor (_14337_, _08093_, _06476_);
  or (_14338_, _14285_, _03139_);
  nor (_14339_, _14338_, _14337_);
  or (_14340_, _14339_, _02575_);
  nor (_14341_, _14340_, _14336_);
  nand (_14342_, _14290_, _05305_);
  and (_14343_, _14342_, _06549_);
  nor (_14344_, _14343_, _14341_);
  and (_14345_, _07968_, _04597_);
  nor (_14346_, _14345_, _14285_);
  and (_14347_, _14346_, _02656_);
  nor (_14348_, _14347_, _14344_);
  and (_14349_, _14348_, _03252_);
  and (_14350_, _08110_, _04597_);
  nor (_14351_, _14350_, _14285_);
  nor (_14352_, _14351_, _03252_);
  or (_14353_, _14352_, _14349_);
  and (_14354_, _14353_, _05332_);
  nor (_14355_, _14354_, _14293_);
  nor (_14356_, _14355_, _03243_);
  nor (_14357_, _14285_, _04888_);
  or (_14358_, _14357_, _03244_);
  nor (_14359_, _14358_, _14304_);
  or (_14360_, _14359_, _02654_);
  nor (_14361_, _14360_, _14356_);
  nor (_14362_, _07967_, _06476_);
  nor (_14363_, _14362_, _14285_);
  and (_14364_, _14363_, _02654_);
  nor (_14365_, _14364_, _14361_);
  and (_14366_, _14365_, _05883_);
  nor (_14367_, _08109_, _06476_);
  nor (_14368_, _14367_, _14285_);
  nor (_14369_, _14368_, _05883_);
  or (_14370_, _14369_, _14366_);
  and (_14371_, _14370_, _03124_);
  nor (_14372_, _14287_, _03124_);
  nor (_14373_, _14372_, _02650_);
  not (_14374_, _14373_);
  nor (_14375_, _14374_, _14371_);
  nor (_14376_, _14285_, _03122_);
  nor (_14377_, _14376_, _14375_);
  and (_14378_, _14377_, _03513_);
  nor (_14379_, _14378_, _14288_);
  nand (_14380_, _14379_, _27788_);
  or (_14381_, _27788_, \oc8051_golden_model_1.TCON [0]);
  and (_14382_, _14381_, _27053_);
  and (_28905_, _14382_, _14380_);
  or (_14383_, _08325_, _06476_);
  or (_14384_, _04597_, \oc8051_golden_model_1.TCON [1]);
  and (_14385_, _14384_, _03251_);
  and (_14386_, _14385_, _14383_);
  nor (_14387_, _08246_, _06529_);
  not (_14388_, \oc8051_golden_model_1.TCON [1]);
  nor (_14389_, _05440_, _14388_);
  or (_14390_, _14389_, _03141_);
  or (_14391_, _14390_, _14387_);
  and (_14392_, _08209_, _04597_);
  not (_14393_, _14392_);
  and (_14394_, _14393_, _14384_);
  or (_14395_, _14394_, _02662_);
  nand (_14396_, _04597_, _08322_);
  and (_14397_, _14396_, _14384_);
  and (_14398_, _14397_, _04505_);
  nor (_14399_, _04505_, _14388_);
  or (_14400_, _14399_, _02661_);
  or (_14401_, _14400_, _14398_);
  and (_14402_, _14401_, _03163_);
  and (_14403_, _14402_, _14395_);
  nor (_14404_, _04597_, _14388_);
  nor (_14405_, _06476_, _03777_);
  or (_14406_, _14405_, _14404_);
  and (_14407_, _14406_, _03162_);
  and (_14408_, _08213_, _05440_);
  or (_14409_, _14408_, _14389_);
  and (_14410_, _14409_, _03150_);
  or (_14411_, _14410_, _14407_);
  or (_14412_, _14411_, _03168_);
  or (_14413_, _14412_, _14403_);
  or (_14414_, _14397_, _03179_);
  and (_14415_, _14414_, _14413_);
  or (_14416_, _14415_, _03176_);
  and (_14417_, _08200_, _05440_);
  or (_14418_, _14417_, _14389_);
  or (_14419_, _14418_, _03177_);
  and (_14420_, _14419_, _05168_);
  and (_14421_, _14420_, _14416_);
  and (_14422_, _08229_, _05440_);
  or (_14423_, _14422_, _14389_);
  and (_14424_, _14423_, _03144_);
  or (_14425_, _14424_, _03140_);
  or (_14426_, _14425_, _14421_);
  and (_14427_, _14426_, _14391_);
  or (_14428_, _14427_, _05949_);
  or (_14429_, _14406_, _06673_);
  and (_14430_, _14429_, _14428_);
  or (_14431_, _14430_, _05959_);
  and (_14432_, _04597_, _04218_);
  or (_14433_, _14404_, _05963_);
  or (_14434_, _14433_, _14432_);
  and (_14435_, _14434_, _03139_);
  and (_14436_, _14435_, _14431_);
  nor (_14437_, _08307_, _06476_);
  or (_14438_, _14437_, _14404_);
  and (_14439_, _14438_, _02024_);
  or (_14440_, _14439_, _14436_);
  and (_14441_, _14440_, _02657_);
  or (_14442_, _08185_, _06476_);
  and (_14443_, _14442_, _02656_);
  nand (_14444_, _04597_, _03016_);
  and (_14445_, _14444_, _02575_);
  or (_14446_, _14445_, _14443_);
  and (_14447_, _14446_, _14384_);
  or (_14448_, _14447_, _14441_);
  and (_14449_, _14448_, _03252_);
  or (_14450_, _14449_, _14386_);
  and (_14451_, _14450_, _05332_);
  or (_14452_, _08184_, _06476_);
  and (_14453_, _14384_, _02669_);
  and (_14454_, _14453_, _14452_);
  or (_14455_, _14454_, _14451_);
  and (_14456_, _14455_, _03244_);
  or (_14457_, _14404_, _06122_);
  and (_14458_, _14397_, _03243_);
  and (_14459_, _14458_, _14457_);
  or (_14460_, _14459_, _14456_);
  and (_14461_, _14460_, _03240_);
  or (_14462_, _14444_, _06122_);
  and (_14463_, _14462_, _02654_);
  or (_14464_, _14396_, _06122_);
  and (_14465_, _14464_, _03239_);
  or (_14466_, _14465_, _14463_);
  and (_14467_, _14466_, _14384_);
  or (_14468_, _14467_, _03123_);
  or (_14469_, _14468_, _14461_);
  or (_14470_, _14394_, _03124_);
  and (_14471_, _14470_, _03122_);
  and (_14472_, _14471_, _14469_);
  and (_14473_, _14418_, _02650_);
  or (_14474_, _14473_, _03121_);
  or (_14475_, _14474_, _14472_);
  or (_14476_, _14392_, _14404_);
  or (_14477_, _14476_, _03513_);
  and (_14478_, _14477_, _14475_);
  and (_14479_, _14478_, _27788_);
  nor (_14480_, _27788_, _14388_);
  or (_14481_, _14480_, rst);
  or (_28906_, _14481_, _14479_);
  not (_14482_, \oc8051_golden_model_1.TCON [2]);
  nor (_14483_, _04597_, _14482_);
  and (_14484_, _04597_, _06009_);
  nor (_14485_, _14484_, _14483_);
  and (_14486_, _14485_, _02575_);
  nor (_14487_, _06476_, _03644_);
  nor (_14488_, _14487_, _14483_);
  and (_14489_, _14488_, _05949_);
  nor (_14490_, _08420_, _06476_);
  nor (_14491_, _14490_, _14483_);
  and (_14492_, _14491_, _02661_);
  and (_14493_, _04597_, \oc8051_golden_model_1.ACC [2]);
  nor (_14494_, _14493_, _14483_);
  nor (_14495_, _14494_, _05903_);
  nor (_14496_, _04505_, _14482_);
  or (_14497_, _14496_, _02661_);
  nor (_14498_, _14497_, _14495_);
  or (_14499_, _14498_, _06504_);
  nor (_14500_, _14499_, _14492_);
  nor (_14501_, _14488_, _03365_);
  nor (_14502_, _05440_, _14482_);
  and (_14503_, _08406_, _05440_);
  nor (_14504_, _14503_, _14502_);
  nor (_14505_, _14504_, _03390_);
  nor (_14506_, _14505_, _14501_);
  nand (_14507_, _14506_, _03179_);
  or (_14508_, _14507_, _14500_);
  nand (_14509_, _14494_, _03168_);
  and (_14510_, _14509_, _14508_);
  nor (_14511_, _14510_, _03176_);
  and (_14512_, _08404_, _05440_);
  nor (_14513_, _14512_, _14502_);
  and (_14514_, _14513_, _03176_);
  or (_14515_, _14514_, _03144_);
  nor (_14516_, _14515_, _14511_);
  and (_14517_, _08447_, _05440_);
  nor (_14518_, _14517_, _14502_);
  nor (_14519_, _14518_, _05168_);
  or (_14520_, _14519_, _14516_);
  and (_14521_, _14520_, _03141_);
  nor (_14522_, _08465_, _06529_);
  nor (_14523_, _14502_, _14522_);
  nor (_14524_, _14523_, _03141_);
  or (_14525_, _14524_, _05949_);
  nor (_14526_, _14525_, _14521_);
  nor (_14527_, _14526_, _14489_);
  nor (_14528_, _14527_, _05959_);
  and (_14529_, _04597_, _04170_);
  nor (_14530_, _14483_, _05963_);
  not (_14531_, _14530_);
  nor (_14532_, _14531_, _14529_);
  or (_14533_, _14532_, _02024_);
  nor (_14534_, _14533_, _14528_);
  nor (_14535_, _08522_, _06476_);
  nor (_14536_, _14535_, _14483_);
  nor (_14537_, _14536_, _03139_);
  or (_14538_, _14537_, _02575_);
  nor (_14539_, _14538_, _14534_);
  nor (_14540_, _14539_, _14486_);
  or (_14541_, _14540_, _02656_);
  and (_14542_, _08537_, _04597_);
  or (_14543_, _14542_, _14483_);
  or (_14544_, _14543_, _05305_);
  and (_14545_, _14544_, _03252_);
  and (_14546_, _14545_, _14541_);
  and (_14547_, _08387_, _04597_);
  nor (_14548_, _14547_, _14483_);
  nor (_14549_, _14548_, _03252_);
  nor (_14550_, _14549_, _14546_);
  nor (_14551_, _14550_, _02669_);
  nor (_14552_, _14483_, _06121_);
  not (_14553_, _14552_);
  nor (_14554_, _14485_, _05332_);
  and (_14555_, _14554_, _14553_);
  nor (_14556_, _14555_, _14551_);
  nor (_14557_, _14556_, _03243_);
  or (_14558_, _14552_, _03244_);
  nor (_14559_, _14558_, _14494_);
  or (_14560_, _14559_, _02654_);
  nor (_14561_, _14560_, _14557_);
  nor (_14562_, _08536_, _06476_);
  nor (_14563_, _14562_, _14483_);
  and (_14564_, _14563_, _02654_);
  nor (_14565_, _14564_, _14561_);
  and (_14566_, _14565_, _05883_);
  nor (_14567_, _08386_, _06476_);
  nor (_14568_, _14567_, _14483_);
  nor (_14569_, _14568_, _05883_);
  or (_14570_, _14569_, _14566_);
  and (_14571_, _14570_, _03124_);
  nor (_14572_, _14491_, _03124_);
  or (_14573_, _14572_, _02650_);
  or (_14574_, _14573_, _14571_);
  nand (_14575_, _14513_, _02650_);
  and (_14576_, _14575_, _14574_);
  nor (_14577_, _14576_, _03121_);
  and (_14578_, _08596_, _04597_);
  nor (_14579_, _14578_, _14483_);
  and (_14580_, _14579_, _03121_);
  nor (_14581_, _14580_, _14577_);
  or (_14582_, _14581_, _27789_);
  or (_14583_, _27788_, \oc8051_golden_model_1.TCON [2]);
  and (_14584_, _14583_, _27053_);
  and (_28907_, _14584_, _14582_);
  not (_14585_, \oc8051_golden_model_1.TCON [3]);
  nor (_14586_, _04597_, _14585_);
  and (_14587_, _04597_, _05986_);
  nor (_14588_, _14587_, _14586_);
  and (_14589_, _14588_, _02575_);
  nor (_14590_, _06476_, _03859_);
  nor (_14591_, _14590_, _14586_);
  and (_14592_, _14591_, _05949_);
  nor (_14593_, _08627_, _06529_);
  nor (_14594_, _05440_, _14585_);
  or (_14595_, _14594_, _03141_);
  or (_14596_, _14595_, _14593_);
  nor (_14597_, _08646_, _06476_);
  nor (_14598_, _14597_, _14586_);
  and (_14599_, _14598_, _02661_);
  and (_14600_, _04597_, \oc8051_golden_model_1.ACC [3]);
  nor (_14601_, _14600_, _14586_);
  nor (_14602_, _14601_, _05903_);
  nor (_14603_, _04505_, _14585_);
  or (_14604_, _14603_, _02661_);
  nor (_14605_, _14604_, _14602_);
  or (_14606_, _14605_, _06504_);
  nor (_14607_, _14606_, _14599_);
  nor (_14608_, _14591_, _03365_);
  and (_14609_, _08642_, _05440_);
  nor (_14610_, _14609_, _14594_);
  nor (_14611_, _14610_, _03390_);
  nor (_14612_, _14611_, _14608_);
  nand (_14613_, _14612_, _03179_);
  or (_14614_, _14613_, _14607_);
  nand (_14615_, _14601_, _03168_);
  and (_14616_, _14615_, _14614_);
  and (_14617_, _14616_, _03177_);
  and (_14618_, _08640_, _05440_);
  nor (_14619_, _14618_, _14594_);
  nor (_14620_, _14619_, _03177_);
  or (_14621_, _14620_, _14617_);
  and (_14622_, _14621_, _05168_);
  nor (_14623_, _14594_, _08671_);
  or (_14624_, _14610_, _05168_);
  nor (_14625_, _14624_, _14623_);
  or (_14626_, _14625_, _03140_);
  or (_14627_, _14626_, _14622_);
  and (_14628_, _14627_, _14596_);
  nor (_14629_, _14628_, _05949_);
  nor (_14630_, _14629_, _14592_);
  nor (_14631_, _14630_, _05959_);
  and (_14632_, _04597_, _04120_);
  nor (_14633_, _14586_, _05963_);
  not (_14634_, _14633_);
  nor (_14635_, _14634_, _14632_);
  or (_14636_, _14635_, _02024_);
  nor (_14637_, _14636_, _14631_);
  nor (_14638_, _08744_, _06476_);
  nor (_14639_, _14638_, _14586_);
  nor (_14640_, _14639_, _03139_);
  or (_14641_, _14640_, _02575_);
  nor (_14642_, _14641_, _14637_);
  nor (_14643_, _14642_, _14589_);
  or (_14644_, _14643_, _02656_);
  and (_14645_, _08622_, _04597_);
  or (_14646_, _14645_, _14586_);
  or (_14647_, _14646_, _05305_);
  and (_14648_, _14647_, _03252_);
  and (_14649_, _14648_, _14644_);
  and (_14650_, _08618_, _04597_);
  nor (_14651_, _14650_, _14586_);
  nor (_14652_, _14651_, _03252_);
  nor (_14653_, _14652_, _14649_);
  nor (_14654_, _14653_, _02669_);
  nor (_14655_, _14586_, _06120_);
  not (_14656_, _14655_);
  nor (_14657_, _14588_, _05332_);
  and (_14658_, _14657_, _14656_);
  nor (_14659_, _14658_, _14654_);
  nor (_14660_, _14659_, _03243_);
  or (_14661_, _14655_, _03244_);
  nor (_14662_, _14661_, _14601_);
  or (_14663_, _14662_, _02654_);
  nor (_14664_, _14663_, _14660_);
  nor (_14665_, _08621_, _06476_);
  nor (_14666_, _14665_, _14586_);
  and (_14667_, _14666_, _02654_);
  nor (_14668_, _14667_, _14664_);
  and (_14669_, _14668_, _05883_);
  nor (_14670_, _08617_, _06476_);
  nor (_14671_, _14670_, _14586_);
  nor (_14672_, _14671_, _05883_);
  or (_14673_, _14672_, _14669_);
  and (_14674_, _14673_, _03124_);
  nor (_14675_, _14598_, _03124_);
  or (_14676_, _14675_, _02650_);
  or (_14677_, _14676_, _14674_);
  nand (_14678_, _14619_, _02650_);
  and (_14679_, _14678_, _14677_);
  nor (_14680_, _14679_, _03121_);
  and (_14681_, _08807_, _04597_);
  nor (_14682_, _14681_, _14586_);
  and (_14683_, _14682_, _03121_);
  nor (_14684_, _14683_, _14680_);
  or (_14685_, _14684_, _27789_);
  or (_14686_, _27788_, \oc8051_golden_model_1.TCON [3]);
  and (_14687_, _14686_, _27053_);
  and (_28908_, _14687_, _14685_);
  not (_14688_, \oc8051_golden_model_1.TCON [4]);
  nor (_14689_, _04597_, _14688_);
  and (_14690_, _04597_, _05974_);
  nor (_14691_, _14690_, _14689_);
  and (_14692_, _14691_, _02575_);
  nor (_14693_, _06476_, _04325_);
  nor (_14694_, _14693_, _14689_);
  and (_14695_, _14694_, _05949_);
  nor (_14696_, _05440_, _14688_);
  nor (_14697_, _14696_, _08889_);
  and (_14698_, _08869_, _05440_);
  nor (_14699_, _14698_, _14696_);
  or (_14700_, _14699_, _05168_);
  nor (_14701_, _14700_, _14697_);
  nor (_14702_, _08838_, _06476_);
  nor (_14703_, _14702_, _14689_);
  and (_14704_, _14703_, _02661_);
  and (_14705_, _04597_, \oc8051_golden_model_1.ACC [4]);
  nor (_14706_, _14705_, _14689_);
  nor (_14707_, _14706_, _05903_);
  nor (_14708_, _04505_, _14688_);
  or (_14709_, _14708_, _02661_);
  nor (_14710_, _14709_, _14707_);
  or (_14711_, _14710_, _06504_);
  nor (_14712_, _14711_, _14704_);
  nor (_14713_, _14694_, _03365_);
  nor (_14714_, _14699_, _03390_);
  nor (_14715_, _14714_, _14713_);
  nand (_14716_, _14715_, _03179_);
  or (_14717_, _14716_, _14712_);
  nand (_14718_, _14706_, _03168_);
  and (_14719_, _14718_, _14717_);
  and (_14720_, _14719_, _03177_);
  and (_14721_, _08880_, _05440_);
  nor (_14722_, _14721_, _14696_);
  nor (_14723_, _14722_, _03177_);
  or (_14724_, _14723_, _14720_);
  and (_14725_, _14724_, _05168_);
  nor (_14726_, _14725_, _14701_);
  nor (_14727_, _14726_, _03140_);
  nor (_14728_, _08908_, _06529_);
  nor (_14729_, _14728_, _14696_);
  nor (_14730_, _14729_, _03141_);
  nor (_14731_, _14730_, _05949_);
  not (_14732_, _14731_);
  nor (_14733_, _14732_, _14727_);
  nor (_14734_, _14733_, _14695_);
  nor (_14735_, _14734_, _05959_);
  and (_14736_, _04597_, _04012_);
  nor (_14737_, _14689_, _05963_);
  not (_14738_, _14737_);
  nor (_14739_, _14738_, _14736_);
  or (_14740_, _14739_, _02024_);
  nor (_14741_, _14740_, _14735_);
  nor (_14742_, _08967_, _06476_);
  nor (_14743_, _14742_, _14689_);
  nor (_14744_, _14743_, _03139_);
  or (_14745_, _14744_, _02575_);
  nor (_14746_, _14745_, _14741_);
  nor (_14747_, _14746_, _14692_);
  or (_14748_, _14747_, _02656_);
  and (_14749_, _08982_, _04597_);
  or (_14750_, _14749_, _14689_);
  or (_14751_, _14750_, _05305_);
  and (_14752_, _14751_, _03252_);
  and (_14753_, _14752_, _14748_);
  and (_14754_, _08830_, _04597_);
  nor (_14755_, _14754_, _14689_);
  nor (_14756_, _14755_, _03252_);
  nor (_14757_, _14756_, _14753_);
  nor (_14758_, _14757_, _02669_);
  nor (_14759_, _14689_, _09034_);
  not (_14760_, _14759_);
  nor (_14761_, _14691_, _05332_);
  and (_14762_, _14761_, _14760_);
  nor (_14763_, _14762_, _14758_);
  nor (_14764_, _14763_, _03243_);
  or (_14765_, _14759_, _03244_);
  nor (_14766_, _14765_, _14706_);
  or (_14767_, _14766_, _02654_);
  nor (_14768_, _14767_, _14764_);
  nor (_14769_, _08981_, _06476_);
  nor (_14770_, _14769_, _14689_);
  and (_14771_, _14770_, _02654_);
  nor (_14772_, _14771_, _14768_);
  and (_14773_, _14772_, _05883_);
  nor (_14774_, _08828_, _06476_);
  nor (_14775_, _14774_, _14689_);
  nor (_14776_, _14775_, _05883_);
  or (_14777_, _14776_, _14773_);
  and (_14778_, _14777_, _03124_);
  nor (_14779_, _14703_, _03124_);
  or (_14780_, _14779_, _02650_);
  or (_14781_, _14780_, _14778_);
  nand (_14782_, _14722_, _02650_);
  and (_14783_, _14782_, _14781_);
  nor (_14784_, _14783_, _03121_);
  and (_14785_, _09037_, _04597_);
  nor (_14786_, _14785_, _14689_);
  and (_14787_, _14786_, _03121_);
  nor (_14788_, _14787_, _14784_);
  or (_14789_, _14788_, _27789_);
  or (_14790_, _27788_, \oc8051_golden_model_1.TCON [4]);
  and (_14791_, _14790_, _27053_);
  and (_28909_, _14791_, _14789_);
  not (_14792_, \oc8051_golden_model_1.TCON [5]);
  nor (_14793_, _04597_, _14792_);
  and (_14794_, _04597_, _06036_);
  nor (_14795_, _14794_, _14793_);
  and (_14796_, _14795_, _02575_);
  nor (_14797_, _06476_, _04480_);
  nor (_14798_, _14797_, _14793_);
  and (_14799_, _14798_, _05949_);
  and (_14800_, _04597_, \oc8051_golden_model_1.ACC [5]);
  nor (_14801_, _14800_, _14793_);
  and (_14802_, _14801_, _03168_);
  nor (_14803_, _09087_, _06476_);
  nor (_14804_, _14803_, _14793_);
  and (_14805_, _14804_, _02661_);
  nor (_14806_, _14801_, _05903_);
  nor (_14807_, _04505_, _14792_);
  or (_14808_, _14807_, _02661_);
  nor (_14809_, _14808_, _14806_);
  or (_14810_, _14809_, _06504_);
  nor (_14811_, _14810_, _14805_);
  nor (_14812_, _14798_, _03365_);
  nor (_14813_, _14812_, _14811_);
  nor (_14814_, _05440_, _14792_);
  and (_14815_, _09072_, _05440_);
  nor (_14816_, _14815_, _14814_);
  nor (_14817_, _14816_, _03390_);
  nor (_14818_, _14817_, _03168_);
  and (_14819_, _14818_, _14813_);
  nor (_14820_, _14819_, _14802_);
  and (_14821_, _14820_, _03177_);
  and (_14822_, _09099_, _05440_);
  nor (_14823_, _14822_, _14814_);
  nor (_14824_, _14823_, _03177_);
  or (_14825_, _14824_, _14821_);
  and (_14826_, _14825_, _05168_);
  nor (_14827_, _14814_, _09107_);
  or (_14828_, _14816_, _05168_);
  nor (_14829_, _14828_, _14827_);
  nor (_14830_, _14829_, _14826_);
  nor (_14831_, _14830_, _03140_);
  nor (_14832_, _09059_, _06529_);
  nor (_14833_, _14832_, _14814_);
  nor (_14834_, _14833_, _03141_);
  nor (_14835_, _14834_, _05949_);
  not (_14836_, _14835_);
  nor (_14837_, _14836_, _14831_);
  nor (_14838_, _14837_, _14799_);
  nor (_14839_, _14838_, _05959_);
  and (_14840_, _04597_, _03904_);
  nor (_14841_, _14793_, _05963_);
  not (_14842_, _14841_);
  nor (_14843_, _14842_, _14840_);
  or (_14844_, _14843_, _02024_);
  nor (_14845_, _14844_, _14839_);
  nor (_14846_, _09180_, _06476_);
  nor (_14847_, _14846_, _14793_);
  nor (_14848_, _14847_, _03139_);
  or (_14849_, _14848_, _02575_);
  nor (_14850_, _14849_, _14845_);
  nor (_14851_, _14850_, _14796_);
  or (_14852_, _14851_, _02656_);
  and (_14853_, _09195_, _04597_);
  or (_14854_, _14853_, _14793_);
  or (_14855_, _14854_, _05305_);
  and (_14856_, _14855_, _03252_);
  and (_14857_, _14856_, _14852_);
  and (_14858_, _09055_, _04597_);
  nor (_14859_, _14858_, _14793_);
  nor (_14860_, _14859_, _03252_);
  nor (_14861_, _14860_, _14857_);
  nor (_14862_, _14861_, _02669_);
  not (_14863_, _14793_);
  and (_14864_, _14863_, _04787_);
  not (_14865_, _14864_);
  nor (_14866_, _14795_, _05332_);
  and (_14867_, _14866_, _14865_);
  nor (_14868_, _14867_, _14862_);
  nor (_14869_, _14868_, _03243_);
  or (_14870_, _14864_, _03244_);
  nor (_14871_, _14870_, _14801_);
  or (_14872_, _14871_, _02654_);
  nor (_14873_, _14872_, _14869_);
  nor (_14874_, _09194_, _06476_);
  nor (_14875_, _14874_, _14793_);
  and (_14876_, _14875_, _02654_);
  nor (_14877_, _14876_, _14873_);
  and (_14878_, _14877_, _05883_);
  nor (_14879_, _09054_, _06476_);
  nor (_14880_, _14879_, _14793_);
  nor (_14881_, _14880_, _05883_);
  or (_14882_, _14881_, _14878_);
  and (_14883_, _14882_, _03124_);
  nor (_14884_, _14804_, _03124_);
  or (_14885_, _14884_, _02650_);
  or (_14886_, _14885_, _14883_);
  nand (_14887_, _14823_, _02650_);
  and (_14888_, _14887_, _14886_);
  nor (_14889_, _14888_, _03121_);
  and (_14890_, _09248_, _04597_);
  nor (_14891_, _14890_, _14793_);
  and (_14892_, _14891_, _03121_);
  nor (_14893_, _14892_, _14889_);
  or (_14894_, _14893_, _27789_);
  or (_14895_, _27788_, \oc8051_golden_model_1.TCON [5]);
  and (_14896_, _14895_, _27053_);
  and (_28910_, _14896_, _14894_);
  not (_14897_, \oc8051_golden_model_1.TCON [6]);
  nor (_14898_, _04597_, _14897_);
  and (_14899_, _04597_, _03960_);
  or (_14900_, _14899_, _14898_);
  and (_14901_, _14900_, _05959_);
  nor (_14902_, _05440_, _14897_);
  not (_14903_, _14902_);
  and (_14904_, _14903_, _09320_);
  and (_14905_, _09305_, _05440_);
  nor (_14906_, _14905_, _14902_);
  or (_14907_, _14906_, _05168_);
  nor (_14908_, _14907_, _14904_);
  nor (_14909_, _09301_, _06476_);
  nor (_14910_, _14909_, _14898_);
  and (_14911_, _14910_, _02661_);
  and (_14912_, _04597_, \oc8051_golden_model_1.ACC [6]);
  nor (_14913_, _14912_, _14898_);
  nor (_14914_, _14913_, _05903_);
  nor (_14915_, _04505_, _14897_);
  or (_14916_, _14915_, _02661_);
  nor (_14917_, _14916_, _14914_);
  or (_14918_, _14917_, _06504_);
  nor (_14919_, _14918_, _14911_);
  nor (_14920_, _06476_, _04373_);
  nor (_14921_, _14920_, _14898_);
  nor (_14922_, _14921_, _03365_);
  nor (_14923_, _14906_, _03390_);
  nor (_14924_, _14923_, _14922_);
  nand (_14925_, _14924_, _03179_);
  or (_14926_, _14925_, _14919_);
  nand (_14927_, _14913_, _03168_);
  and (_14928_, _14927_, _14926_);
  and (_14929_, _14928_, _03177_);
  and (_14930_, _09286_, _05440_);
  nor (_14931_, _14930_, _14902_);
  nor (_14932_, _14931_, _03177_);
  or (_14933_, _14932_, _14929_);
  and (_14934_, _14933_, _05168_);
  nor (_14935_, _14934_, _14908_);
  nor (_14936_, _14935_, _03140_);
  nor (_14937_, _09272_, _06529_);
  nor (_14938_, _14937_, _14902_);
  nor (_14939_, _14938_, _03141_);
  nor (_14940_, _14939_, _05949_);
  not (_14941_, _14940_);
  nor (_14942_, _14941_, _14936_);
  and (_14943_, _14921_, _05949_);
  or (_14944_, _14943_, _05959_);
  nor (_14945_, _14944_, _14942_);
  or (_14946_, _14945_, _14901_);
  and (_14947_, _14946_, _03139_);
  and (_14948_, _09388_, _04597_);
  nor (_14949_, _14948_, _14898_);
  nor (_14950_, _14949_, _03139_);
  or (_14951_, _14950_, _06549_);
  or (_14952_, _14951_, _14947_);
  and (_14953_, _09404_, _04597_);
  or (_14954_, _14898_, _05305_);
  or (_14955_, _14954_, _14953_);
  and (_14956_, _04597_, _09395_);
  nor (_14957_, _14956_, _14898_);
  and (_14958_, _14957_, _02575_);
  nor (_14959_, _14958_, _03251_);
  and (_14960_, _14959_, _14955_);
  and (_14961_, _14960_, _14952_);
  and (_14962_, _09268_, _04597_);
  nor (_14963_, _14962_, _14898_);
  nor (_14964_, _14963_, _03252_);
  nor (_14965_, _14964_, _14961_);
  nor (_14966_, _14965_, _02669_);
  nor (_14967_, _14898_, _06119_);
  not (_14968_, _14967_);
  nor (_14969_, _14957_, _05332_);
  and (_14970_, _14969_, _14968_);
  nor (_14971_, _14970_, _14966_);
  nor (_14972_, _14971_, _03243_);
  or (_14973_, _14967_, _03244_);
  nor (_14974_, _14973_, _14913_);
  or (_14975_, _14974_, _02654_);
  nor (_14976_, _14975_, _14972_);
  nor (_14977_, _09403_, _06476_);
  nor (_14978_, _14977_, _14898_);
  and (_14979_, _14978_, _02654_);
  nor (_14980_, _14979_, _14976_);
  and (_14981_, _14980_, _05883_);
  nor (_14982_, _09267_, _06476_);
  nor (_14983_, _14982_, _14898_);
  nor (_14984_, _14983_, _05883_);
  or (_14985_, _14984_, _14981_);
  and (_14986_, _14985_, _03124_);
  nor (_14987_, _14910_, _03124_);
  or (_14988_, _14987_, _02650_);
  or (_14989_, _14988_, _14986_);
  nand (_14990_, _14931_, _02650_);
  and (_14991_, _14990_, _14989_);
  nor (_14992_, _14991_, _03121_);
  and (_14993_, _09456_, _04597_);
  nor (_14994_, _14993_, _14898_);
  and (_14995_, _14994_, _03121_);
  nor (_14996_, _14995_, _14992_);
  or (_14997_, _14996_, _27789_);
  or (_14998_, _27788_, \oc8051_golden_model_1.TCON [6]);
  and (_14999_, _14998_, _27053_);
  and (_28912_, _14999_, _14997_);
  not (_15000_, \oc8051_golden_model_1.TH0 [0]);
  nor (_15001_, _04612_, _15000_);
  nor (_15002_, _08109_, _06402_);
  nor (_15003_, _15002_, _15001_);
  nor (_15004_, _15003_, _05883_);
  and (_15005_, _04612_, \oc8051_golden_model_1.ACC [0]);
  nor (_15006_, _15005_, _15001_);
  nor (_15007_, _15006_, _03179_);
  nor (_15008_, _15007_, _05949_);
  nor (_15009_, _04888_, _06402_);
  nor (_15010_, _15009_, _15001_);
  nor (_15011_, _15010_, _02662_);
  nor (_15012_, _04505_, _15000_);
  nor (_15013_, _15006_, _05903_);
  nor (_15014_, _15013_, _15012_);
  nor (_15015_, _15014_, _02661_);
  or (_15016_, _15015_, _03162_);
  nor (_15017_, _15016_, _15011_);
  or (_15018_, _15017_, _03168_);
  and (_15019_, _15018_, _15008_);
  and (_15020_, _04612_, _03716_);
  or (_15021_, _15001_, _12270_);
  nor (_15022_, _15021_, _15020_);
  nor (_15023_, _15022_, _15019_);
  nor (_15024_, _15023_, _05959_);
  and (_15025_, _04612_, _04268_);
  nor (_15026_, _15001_, _05963_);
  not (_15027_, _15026_);
  nor (_15028_, _15027_, _15025_);
  nor (_15029_, _15028_, _15024_);
  nor (_15030_, _15029_, _02024_);
  nor (_15031_, _08093_, _06402_);
  or (_15032_, _15001_, _03139_);
  nor (_15033_, _15032_, _15031_);
  or (_15034_, _15033_, _02575_);
  nor (_15035_, _15034_, _15030_);
  and (_15036_, _04612_, _05996_);
  nor (_15037_, _15036_, _15001_);
  nand (_15038_, _15037_, _05305_);
  and (_15039_, _15038_, _06549_);
  nor (_15040_, _15039_, _15035_);
  and (_15041_, _07968_, _04612_);
  nor (_15042_, _15041_, _15001_);
  and (_15043_, _15042_, _02656_);
  nor (_15044_, _15043_, _15040_);
  and (_15045_, _15044_, _03252_);
  and (_15046_, _08110_, _04612_);
  nor (_15047_, _15046_, _15001_);
  nor (_15048_, _15047_, _03252_);
  or (_15049_, _15048_, _15045_);
  and (_15050_, _15049_, _05332_);
  or (_15051_, _15037_, _05332_);
  nor (_15052_, _15051_, _15009_);
  nor (_15053_, _15052_, _15050_);
  nor (_15054_, _15053_, _03243_);
  and (_15055_, _08108_, _04612_);
  or (_15056_, _15055_, _15001_);
  and (_15057_, _15056_, _03243_);
  or (_15058_, _15057_, _15054_);
  and (_15059_, _15058_, _05357_);
  nor (_15060_, _07967_, _06402_);
  nor (_15061_, _15060_, _15001_);
  nor (_15062_, _15061_, _05357_);
  or (_15063_, _15062_, _15059_);
  and (_15064_, _15063_, _05883_);
  or (_15065_, _15064_, _11672_);
  nor (_15066_, _15065_, _15004_);
  and (_15067_, _15010_, _11672_);
  nor (_15068_, _15067_, _15066_);
  or (_15069_, _15068_, _27789_);
  or (_15070_, _27788_, \oc8051_golden_model_1.TH0 [0]);
  and (_15071_, _15070_, _27053_);
  and (_28913_, _15071_, _15069_);
  nor (_15072_, _04612_, \oc8051_golden_model_1.TH0 [1]);
  and (_15073_, _08209_, _04612_);
  nor (_15074_, _15073_, _15072_);
  nor (_15075_, _15074_, _03124_);
  not (_15076_, _15072_);
  nor (_15077_, _08184_, _06402_);
  nor (_15078_, _15077_, _05332_);
  and (_15079_, _15078_, _15076_);
  nor (_15080_, _08325_, _06402_);
  nor (_15081_, _15080_, _03252_);
  and (_15082_, _15081_, _15076_);
  and (_15083_, _04612_, _04218_);
  not (_15084_, \oc8051_golden_model_1.TH0 [1]);
  nor (_15085_, _04612_, _15084_);
  nor (_15086_, _15085_, _05963_);
  not (_15087_, _15086_);
  nor (_15088_, _15087_, _15083_);
  not (_15089_, _15088_);
  and (_15090_, _04612_, _08322_);
  nor (_15091_, _15090_, _15072_);
  and (_15092_, _15091_, _03168_);
  and (_15093_, _15091_, _04505_);
  nor (_15094_, _04505_, _15084_);
  or (_15095_, _15094_, _15093_);
  and (_15096_, _15095_, _02662_);
  and (_15097_, _15074_, _02661_);
  or (_15098_, _15097_, _15096_);
  and (_15099_, _15098_, _03365_);
  nor (_15100_, _06402_, _03777_);
  nor (_15101_, _15100_, _15085_);
  nor (_15102_, _15101_, _03365_);
  nor (_15103_, _15102_, _15099_);
  nor (_15104_, _15103_, _03168_);
  or (_15105_, _15104_, _05949_);
  nor (_15106_, _15105_, _15092_);
  and (_15107_, _15101_, _05949_);
  nor (_15108_, _15107_, _15106_);
  nor (_15109_, _15108_, _05959_);
  nor (_15110_, _15109_, _02024_);
  and (_15111_, _15110_, _15089_);
  and (_15112_, _08307_, _04612_);
  nor (_15113_, _15112_, _03139_);
  and (_15114_, _15113_, _15076_);
  nor (_15115_, _15114_, _15111_);
  nor (_15116_, _15115_, _06549_);
  nor (_15117_, _08185_, _06402_);
  nor (_15118_, _15117_, _05305_);
  and (_15119_, _04612_, _03016_);
  nor (_15120_, _15119_, _05245_);
  or (_15121_, _15120_, _15118_);
  and (_15122_, _15121_, _15076_);
  nor (_15123_, _15122_, _15116_);
  nor (_15124_, _15123_, _03251_);
  nor (_15125_, _15124_, _15082_);
  nor (_15126_, _15125_, _02669_);
  nor (_15127_, _15126_, _15079_);
  nor (_15128_, _15127_, _03243_);
  nor (_15129_, _15085_, _06122_);
  nor (_15130_, _15129_, _03244_);
  and (_15131_, _15130_, _15091_);
  nor (_15132_, _15131_, _15128_);
  nor (_15133_, _15132_, _03241_);
  and (_15134_, _15119_, _04835_);
  nor (_15135_, _15134_, _05357_);
  nand (_15136_, _15090_, _04835_);
  and (_15137_, _15136_, _03239_);
  or (_15138_, _15137_, _15135_);
  and (_15139_, _15138_, _15076_);
  or (_15140_, _15139_, _03123_);
  nor (_15141_, _15140_, _15133_);
  nor (_15142_, _15141_, _15075_);
  nor (_15143_, _15142_, _03121_);
  nor (_15144_, _15085_, _15073_);
  and (_15145_, _15144_, _03121_);
  nor (_15146_, _15145_, _15143_);
  or (_15147_, _15146_, _27789_);
  or (_15148_, _27788_, \oc8051_golden_model_1.TH0 [1]);
  and (_15149_, _15148_, _27053_);
  and (_28914_, _15149_, _15147_);
  not (_15150_, \oc8051_golden_model_1.TH0 [2]);
  nor (_15151_, _04612_, _15150_);
  nor (_15152_, _15151_, _06121_);
  not (_15153_, _15152_);
  and (_15154_, _04612_, _06009_);
  nor (_15155_, _15154_, _15151_);
  nor (_15156_, _15155_, _05332_);
  and (_15157_, _15156_, _15153_);
  and (_15158_, _04612_, _04170_);
  nor (_15159_, _15158_, _15151_);
  or (_15160_, _15159_, _05963_);
  and (_15161_, _04612_, \oc8051_golden_model_1.ACC [2]);
  nor (_15162_, _15161_, _15151_);
  nor (_15163_, _15162_, _03179_);
  nor (_15164_, _15162_, _05903_);
  nor (_15165_, _04505_, _15150_);
  or (_15166_, _15165_, _15164_);
  and (_15167_, _15166_, _02662_);
  nor (_15168_, _08420_, _06402_);
  nor (_15169_, _15168_, _15151_);
  nor (_15170_, _15169_, _02662_);
  or (_15171_, _15170_, _15167_);
  and (_15172_, _15171_, _03365_);
  nor (_15173_, _06402_, _03644_);
  nor (_15174_, _15173_, _15151_);
  nor (_15175_, _15174_, _03365_);
  nor (_15176_, _15175_, _15172_);
  nor (_15177_, _15176_, _03168_);
  or (_15178_, _15177_, _05949_);
  nor (_15179_, _15178_, _15163_);
  and (_15180_, _15174_, _05949_);
  or (_15181_, _15180_, _05959_);
  or (_15182_, _15181_, _15179_);
  and (_15183_, _15182_, _03139_);
  and (_15184_, _15183_, _15160_);
  nor (_15185_, _08522_, _06402_);
  or (_15186_, _15151_, _03139_);
  nor (_15187_, _15186_, _15185_);
  or (_15188_, _15187_, _02575_);
  nor (_15189_, _15188_, _15184_);
  nand (_15190_, _15155_, _05305_);
  and (_15191_, _15190_, _06549_);
  nor (_15192_, _15191_, _15189_);
  and (_15193_, _08537_, _04612_);
  nor (_15194_, _15193_, _15151_);
  and (_15195_, _15194_, _02656_);
  nor (_15196_, _15195_, _15192_);
  and (_15197_, _15196_, _03252_);
  and (_15198_, _08387_, _04612_);
  nor (_15199_, _15198_, _15151_);
  nor (_15200_, _15199_, _03252_);
  or (_15201_, _15200_, _15197_);
  and (_15202_, _15201_, _05332_);
  nor (_15203_, _15202_, _15157_);
  nor (_15204_, _15203_, _03243_);
  or (_15205_, _15152_, _03244_);
  nor (_15206_, _15205_, _15162_);
  or (_15207_, _15206_, _02654_);
  nor (_15208_, _15207_, _15204_);
  nor (_15209_, _08536_, _06402_);
  nor (_15210_, _15209_, _15151_);
  and (_15211_, _15210_, _02654_);
  nor (_15212_, _15211_, _15208_);
  and (_15213_, _15212_, _05883_);
  nor (_15214_, _08386_, _06402_);
  nor (_15215_, _15214_, _15151_);
  nor (_15216_, _15215_, _05883_);
  or (_15217_, _15216_, _15213_);
  and (_15218_, _15217_, _03124_);
  nor (_15219_, _15169_, _03124_);
  or (_15220_, _15219_, _15218_);
  and (_15221_, _15220_, _03513_);
  and (_15222_, _08596_, _04612_);
  nor (_15223_, _15222_, _15151_);
  nor (_15224_, _15223_, _03513_);
  or (_15225_, _15224_, _15221_);
  or (_15226_, _15225_, _27789_);
  or (_15227_, _27788_, \oc8051_golden_model_1.TH0 [2]);
  and (_15228_, _15227_, _27053_);
  and (_28915_, _15228_, _15226_);
  not (_15229_, \oc8051_golden_model_1.TH0 [3]);
  nor (_15230_, _04612_, _15229_);
  nor (_15231_, _15230_, _06120_);
  not (_15232_, _15231_);
  and (_15233_, _04612_, _05986_);
  nor (_15234_, _15233_, _15230_);
  nor (_15235_, _15234_, _05332_);
  and (_15236_, _15235_, _15232_);
  and (_15237_, _04612_, \oc8051_golden_model_1.ACC [3]);
  nor (_15238_, _15237_, _15230_);
  nor (_15239_, _15238_, _05903_);
  nor (_15240_, _04505_, _15229_);
  or (_15241_, _15240_, _15239_);
  and (_15242_, _15241_, _02662_);
  nor (_15243_, _08646_, _06402_);
  nor (_15244_, _15243_, _15230_);
  nor (_15245_, _15244_, _02662_);
  or (_15246_, _15245_, _15242_);
  and (_15247_, _15246_, _03365_);
  nor (_15248_, _06402_, _03859_);
  nor (_15249_, _15248_, _15230_);
  nor (_15250_, _15249_, _03365_);
  nor (_15251_, _15250_, _15247_);
  nor (_15252_, _15251_, _03168_);
  nor (_15253_, _15238_, _03179_);
  nor (_15254_, _15253_, _05949_);
  not (_15255_, _15254_);
  nor (_15256_, _15255_, _15252_);
  and (_15257_, _15249_, _05949_);
  or (_15258_, _15257_, _05959_);
  or (_15259_, _15258_, _15256_);
  and (_15260_, _04612_, _04120_);
  nor (_15261_, _15260_, _15230_);
  or (_15262_, _15261_, _05963_);
  and (_15263_, _15262_, _03139_);
  and (_15264_, _15263_, _15259_);
  nor (_15265_, _08744_, _06402_);
  or (_15266_, _15230_, _03139_);
  nor (_15267_, _15266_, _15265_);
  or (_15268_, _15267_, _02575_);
  nor (_15269_, _15268_, _15264_);
  nand (_15270_, _15234_, _05305_);
  and (_15271_, _15270_, _06549_);
  nor (_15272_, _15271_, _15269_);
  and (_15273_, _08622_, _04612_);
  nor (_15274_, _15273_, _15230_);
  and (_15275_, _15274_, _02656_);
  nor (_15276_, _15275_, _15272_);
  and (_15277_, _15276_, _03252_);
  and (_15278_, _08618_, _04612_);
  nor (_15279_, _15278_, _15230_);
  nor (_15280_, _15279_, _03252_);
  or (_15281_, _15280_, _15277_);
  and (_15282_, _15281_, _05332_);
  nor (_15283_, _15282_, _15236_);
  nor (_15284_, _15283_, _03243_);
  or (_15285_, _15231_, _03244_);
  nor (_15286_, _15285_, _15238_);
  or (_15287_, _15286_, _02654_);
  nor (_15288_, _15287_, _15284_);
  nor (_15289_, _08621_, _06402_);
  nor (_15290_, _15289_, _15230_);
  and (_15291_, _15290_, _02654_);
  nor (_15292_, _15291_, _15288_);
  and (_15293_, _15292_, _05883_);
  nor (_15294_, _08617_, _06402_);
  nor (_15295_, _15294_, _15230_);
  nor (_15296_, _15295_, _05883_);
  or (_15297_, _15296_, _15293_);
  and (_15298_, _15297_, _03124_);
  nor (_15299_, _15244_, _03124_);
  or (_15300_, _15299_, _15298_);
  and (_15301_, _15300_, _03513_);
  and (_15302_, _08807_, _04612_);
  nor (_15303_, _15302_, _15230_);
  nor (_15304_, _15303_, _03513_);
  or (_15305_, _15304_, _15301_);
  or (_15306_, _15305_, _27789_);
  or (_15307_, _27788_, \oc8051_golden_model_1.TH0 [3]);
  and (_15308_, _15307_, _27053_);
  and (_28916_, _15308_, _15306_);
  not (_15309_, \oc8051_golden_model_1.TH0 [4]);
  nor (_15310_, _04612_, _15309_);
  and (_15311_, _08830_, _04612_);
  nor (_15312_, _15311_, _15310_);
  nor (_15313_, _15312_, _03252_);
  and (_15314_, _04612_, _05974_);
  nor (_15315_, _15314_, _15310_);
  and (_15316_, _15315_, _02575_);
  and (_15317_, _04612_, \oc8051_golden_model_1.ACC [4]);
  nor (_15318_, _15317_, _15310_);
  nor (_15319_, _15318_, _03179_);
  nor (_15320_, _15318_, _05903_);
  nor (_15321_, _04505_, _15309_);
  or (_15322_, _15321_, _15320_);
  and (_15323_, _15322_, _02662_);
  nor (_15324_, _08838_, _06402_);
  nor (_15325_, _15324_, _15310_);
  nor (_15326_, _15325_, _02662_);
  or (_15327_, _15326_, _15323_);
  and (_15328_, _15327_, _03365_);
  nor (_15329_, _06402_, _04325_);
  nor (_15330_, _15329_, _15310_);
  nor (_15331_, _15330_, _03365_);
  nor (_15332_, _15331_, _15328_);
  nor (_15333_, _15332_, _03168_);
  or (_15334_, _15333_, _05949_);
  nor (_15335_, _15334_, _15319_);
  and (_15336_, _15330_, _05949_);
  nor (_15337_, _15336_, _15335_);
  nor (_15338_, _15337_, _05959_);
  and (_15339_, _04612_, _04012_);
  nor (_15340_, _15310_, _05963_);
  not (_15341_, _15340_);
  nor (_15342_, _15341_, _15339_);
  or (_15343_, _15342_, _02024_);
  nor (_15344_, _15343_, _15338_);
  nor (_15345_, _08967_, _06402_);
  nor (_15346_, _15345_, _15310_);
  nor (_15347_, _15346_, _03139_);
  or (_15348_, _15347_, _02575_);
  nor (_15349_, _15348_, _15344_);
  nor (_15350_, _15349_, _15316_);
  or (_15351_, _15350_, _02656_);
  and (_15352_, _08982_, _04612_);
  or (_15353_, _15352_, _15310_);
  or (_15354_, _15353_, _05305_);
  and (_15355_, _15354_, _03252_);
  and (_15356_, _15355_, _15351_);
  nor (_15357_, _15356_, _15313_);
  nor (_15358_, _15357_, _02669_);
  nor (_15359_, _15310_, _09034_);
  not (_15360_, _15359_);
  nor (_15361_, _15315_, _05332_);
  and (_15362_, _15361_, _15360_);
  nor (_15363_, _15362_, _15358_);
  nor (_15364_, _15363_, _03243_);
  or (_15365_, _15359_, _03244_);
  nor (_15366_, _15365_, _15318_);
  or (_15367_, _15366_, _02654_);
  nor (_15368_, _15367_, _15364_);
  nor (_15369_, _08981_, _06402_);
  nor (_15370_, _15369_, _15310_);
  and (_15371_, _15370_, _02654_);
  nor (_15372_, _15371_, _15368_);
  and (_15373_, _15372_, _05883_);
  nor (_15374_, _08828_, _06402_);
  nor (_15375_, _15374_, _15310_);
  nor (_15376_, _15375_, _05883_);
  or (_15377_, _15376_, _15373_);
  and (_15378_, _15377_, _03124_);
  nor (_15379_, _15325_, _03124_);
  or (_15380_, _15379_, _15378_);
  and (_15381_, _15380_, _03513_);
  and (_15382_, _09037_, _04612_);
  nor (_15383_, _15382_, _15310_);
  nor (_15384_, _15383_, _03513_);
  or (_15385_, _15384_, _15381_);
  or (_15386_, _15385_, _27789_);
  or (_15387_, _27788_, \oc8051_golden_model_1.TH0 [4]);
  and (_15388_, _15387_, _27053_);
  and (_28917_, _15388_, _15386_);
  not (_15389_, \oc8051_golden_model_1.TH0 [5]);
  nor (_15390_, _04612_, _15389_);
  and (_15391_, _09055_, _04612_);
  nor (_15392_, _15391_, _15390_);
  nor (_15393_, _15392_, _03252_);
  and (_15394_, _04612_, _06036_);
  nor (_15395_, _15394_, _15390_);
  and (_15396_, _15395_, _02575_);
  nor (_15397_, _06402_, _04480_);
  nor (_15398_, _15397_, _15390_);
  and (_15399_, _15398_, _05949_);
  and (_15400_, _04612_, \oc8051_golden_model_1.ACC [5]);
  nor (_15401_, _15400_, _15390_);
  nor (_15402_, _15401_, _05903_);
  nor (_15403_, _04505_, _15389_);
  or (_15404_, _15403_, _15402_);
  and (_15405_, _15404_, _02662_);
  nor (_15406_, _09087_, _06402_);
  nor (_15407_, _15406_, _15390_);
  nor (_15408_, _15407_, _02662_);
  or (_15409_, _15408_, _15405_);
  and (_15410_, _15409_, _03365_);
  nor (_15411_, _15398_, _03365_);
  nor (_15412_, _15411_, _15410_);
  nor (_15413_, _15412_, _03168_);
  nor (_15414_, _15401_, _03179_);
  nor (_15415_, _15414_, _05949_);
  not (_15416_, _15415_);
  nor (_15417_, _15416_, _15413_);
  nor (_15418_, _15417_, _15399_);
  nor (_15419_, _15418_, _05959_);
  and (_15420_, _04612_, _03904_);
  nor (_15421_, _15390_, _05963_);
  not (_15422_, _15421_);
  nor (_15423_, _15422_, _15420_);
  or (_15424_, _15423_, _02024_);
  nor (_15425_, _15424_, _15419_);
  nor (_15426_, _09180_, _06402_);
  nor (_15427_, _15426_, _15390_);
  nor (_15428_, _15427_, _03139_);
  or (_15429_, _15428_, _02575_);
  nor (_15430_, _15429_, _15425_);
  nor (_15431_, _15430_, _15396_);
  or (_15432_, _15431_, _02656_);
  and (_15433_, _09195_, _04612_);
  or (_15434_, _15433_, _15390_);
  or (_15435_, _15434_, _05305_);
  and (_15436_, _15435_, _03252_);
  and (_15437_, _15436_, _15432_);
  nor (_15438_, _15437_, _15393_);
  nor (_15439_, _15438_, _02669_);
  not (_15440_, _15390_);
  and (_15441_, _15440_, _04787_);
  not (_15442_, _15441_);
  nor (_15443_, _15395_, _05332_);
  and (_15444_, _15443_, _15442_);
  nor (_15445_, _15444_, _15439_);
  nor (_15446_, _15445_, _03243_);
  or (_15447_, _15441_, _03244_);
  nor (_15448_, _15447_, _15401_);
  or (_15449_, _15448_, _02654_);
  nor (_15450_, _15449_, _15446_);
  nor (_15451_, _09194_, _06402_);
  nor (_15452_, _15451_, _15390_);
  and (_15453_, _15452_, _02654_);
  nor (_15454_, _15453_, _15450_);
  and (_15455_, _15454_, _05883_);
  nor (_15456_, _09054_, _06402_);
  nor (_15457_, _15456_, _15390_);
  nor (_15458_, _15457_, _05883_);
  or (_15459_, _15458_, _15455_);
  and (_15460_, _15459_, _03124_);
  nor (_15461_, _15407_, _03124_);
  or (_15462_, _15461_, _15460_);
  and (_15463_, _15462_, _03513_);
  and (_15464_, _09248_, _04612_);
  nor (_15465_, _15464_, _15390_);
  nor (_15466_, _15465_, _03513_);
  or (_15467_, _15466_, _15463_);
  or (_15468_, _15467_, _27789_);
  or (_15469_, _27788_, \oc8051_golden_model_1.TH0 [5]);
  and (_15470_, _15469_, _27053_);
  and (_28918_, _15470_, _15468_);
  not (_15471_, \oc8051_golden_model_1.TH0 [6]);
  nor (_15472_, _04612_, _15471_);
  nor (_15473_, _15472_, _06119_);
  not (_15474_, _15473_);
  and (_15475_, _04612_, _09395_);
  nor (_15476_, _15475_, _15472_);
  nor (_15477_, _15476_, _05332_);
  and (_15478_, _15477_, _15474_);
  and (_15479_, _09268_, _04612_);
  nor (_15480_, _15479_, _15472_);
  nor (_15481_, _15480_, _03252_);
  and (_15482_, _04612_, _03960_);
  or (_15483_, _15482_, _15472_);
  and (_15484_, _15483_, _05959_);
  and (_15485_, _04612_, \oc8051_golden_model_1.ACC [6]);
  nor (_15486_, _15485_, _15472_);
  nor (_15487_, _15486_, _03179_);
  nor (_15488_, _15486_, _05903_);
  nor (_15489_, _04505_, _15471_);
  or (_15490_, _15489_, _15488_);
  and (_15491_, _15490_, _02662_);
  nor (_15492_, _09301_, _06402_);
  nor (_15493_, _15492_, _15472_);
  nor (_15494_, _15493_, _02662_);
  or (_15495_, _15494_, _15491_);
  and (_15496_, _15495_, _03365_);
  nor (_15497_, _06402_, _04373_);
  nor (_15498_, _15497_, _15472_);
  nor (_15499_, _15498_, _03365_);
  nor (_15500_, _15499_, _15496_);
  nor (_15501_, _15500_, _03168_);
  or (_15502_, _15501_, _05949_);
  nor (_15503_, _15502_, _15487_);
  and (_15504_, _15498_, _05949_);
  or (_15505_, _15504_, _05959_);
  nor (_15506_, _15505_, _15503_);
  or (_15507_, _15506_, _15484_);
  and (_15508_, _15507_, _03139_);
  and (_15509_, _09388_, _04612_);
  nor (_15510_, _15509_, _15472_);
  nor (_15511_, _15510_, _03139_);
  or (_15512_, _15511_, _06549_);
  or (_15513_, _15512_, _15508_);
  and (_15514_, _09404_, _04612_);
  or (_15515_, _15472_, _05305_);
  or (_15516_, _15515_, _15514_);
  and (_15517_, _15476_, _02575_);
  nor (_15518_, _15517_, _03251_);
  and (_15519_, _15518_, _15516_);
  and (_15520_, _15519_, _15513_);
  nor (_15521_, _15520_, _15481_);
  nor (_15522_, _15521_, _02669_);
  nor (_15523_, _15522_, _15478_);
  nor (_15524_, _15523_, _03243_);
  or (_15525_, _15473_, _03244_);
  nor (_15526_, _15525_, _15486_);
  or (_15527_, _15526_, _02654_);
  nor (_15528_, _15527_, _15524_);
  nor (_15529_, _09403_, _06402_);
  nor (_15530_, _15529_, _15472_);
  and (_15531_, _15530_, _02654_);
  nor (_15532_, _15531_, _15528_);
  and (_15533_, _15532_, _05883_);
  nor (_15534_, _09267_, _06402_);
  nor (_15535_, _15534_, _15472_);
  nor (_15536_, _15535_, _05883_);
  or (_15537_, _15536_, _15533_);
  and (_15538_, _15537_, _03124_);
  nor (_15539_, _15493_, _03124_);
  or (_15540_, _15539_, _15538_);
  and (_15541_, _15540_, _03513_);
  and (_15542_, _09456_, _04612_);
  nor (_15543_, _15542_, _15472_);
  nor (_15544_, _15543_, _03513_);
  or (_15545_, _15544_, _15541_);
  or (_15546_, _15545_, _27789_);
  or (_15547_, _27788_, \oc8051_golden_model_1.TH0 [6]);
  and (_15548_, _15547_, _27053_);
  and (_28919_, _15548_, _15546_);
  not (_15549_, \oc8051_golden_model_1.TH1 [0]);
  nor (_15550_, _04594_, _15549_);
  nor (_15551_, _04888_, _06316_);
  nor (_15552_, _15551_, _15550_);
  and (_15553_, _15552_, _11672_);
  and (_15554_, _04594_, _03716_);
  nor (_15555_, _15554_, _15550_);
  and (_15556_, _15555_, _05949_);
  and (_15557_, _04594_, \oc8051_golden_model_1.ACC [0]);
  nor (_15558_, _15557_, _15550_);
  nor (_15559_, _15558_, _05903_);
  nor (_15560_, _04505_, _15549_);
  or (_15561_, _15560_, _15559_);
  and (_15562_, _15561_, _02662_);
  nor (_15563_, _15552_, _02662_);
  or (_15564_, _15563_, _15562_);
  and (_15565_, _15564_, _03365_);
  nor (_15566_, _15555_, _03365_);
  nor (_15567_, _15566_, _15565_);
  nor (_15568_, _15567_, _03168_);
  nor (_15569_, _15558_, _03179_);
  nor (_15570_, _15569_, _05949_);
  not (_15571_, _15570_);
  nor (_15572_, _15571_, _15568_);
  nor (_15573_, _15572_, _15556_);
  nor (_15574_, _15573_, _05959_);
  and (_15575_, _04594_, _04268_);
  nor (_15576_, _15550_, _05963_);
  not (_15577_, _15576_);
  nor (_15578_, _15577_, _15575_);
  nor (_15579_, _15578_, _15574_);
  nor (_15580_, _15579_, _02024_);
  nor (_15581_, _08093_, _06316_);
  or (_15582_, _15550_, _03139_);
  nor (_15583_, _15582_, _15581_);
  or (_15584_, _15583_, _02575_);
  nor (_15585_, _15584_, _15580_);
  and (_15586_, _04594_, _05996_);
  nor (_15587_, _15586_, _15550_);
  nand (_15588_, _15587_, _05305_);
  and (_15589_, _15588_, _06549_);
  nor (_15590_, _15589_, _15585_);
  and (_15591_, _07968_, _04594_);
  nor (_15592_, _15591_, _15550_);
  and (_15593_, _15592_, _02656_);
  nor (_15594_, _15593_, _15590_);
  and (_15595_, _15594_, _03252_);
  and (_15596_, _08110_, _04594_);
  nor (_15597_, _15596_, _15550_);
  nor (_15598_, _15597_, _03252_);
  or (_15599_, _15598_, _15595_);
  and (_15600_, _15599_, _05332_);
  or (_15601_, _15587_, _05332_);
  nor (_15602_, _15601_, _15551_);
  nor (_15603_, _15602_, _15600_);
  nor (_15604_, _15603_, _03243_);
  and (_15605_, _08108_, _04594_);
  or (_15606_, _15605_, _15550_);
  and (_15607_, _15606_, _03243_);
  or (_15608_, _15607_, _15604_);
  and (_15609_, _15608_, _05357_);
  nor (_15610_, _07967_, _06316_);
  nor (_15611_, _15610_, _15550_);
  nor (_15612_, _15611_, _05357_);
  or (_15613_, _15612_, _15609_);
  and (_15614_, _15613_, _05883_);
  nor (_15615_, _08109_, _06316_);
  nor (_15616_, _15615_, _15550_);
  nor (_15617_, _15616_, _05883_);
  nor (_15618_, _15617_, _11672_);
  not (_15619_, _15618_);
  nor (_15620_, _15619_, _15614_);
  nor (_15621_, _15620_, _15553_);
  or (_15622_, _15621_, _27789_);
  or (_15623_, _27788_, \oc8051_golden_model_1.TH1 [0]);
  and (_15624_, _15623_, _27053_);
  and (_28922_, _15624_, _15622_);
  nor (_15625_, _04594_, \oc8051_golden_model_1.TH1 [1]);
  and (_15626_, _08209_, _04594_);
  nor (_15627_, _15626_, _15625_);
  nor (_15628_, _15627_, _03124_);
  not (_15629_, _15625_);
  nor (_15630_, _08184_, _06316_);
  nor (_15631_, _15630_, _05332_);
  and (_15632_, _15631_, _15629_);
  nor (_15633_, _08325_, _06316_);
  nor (_15634_, _15633_, _03252_);
  and (_15635_, _15634_, _15629_);
  and (_15636_, _04594_, _04218_);
  not (_15637_, \oc8051_golden_model_1.TH1 [1]);
  nor (_15638_, _04594_, _15637_);
  nor (_15639_, _15638_, _05963_);
  not (_15640_, _15639_);
  nor (_15641_, _15640_, _15636_);
  not (_15642_, _15641_);
  nor (_15643_, _06316_, _03777_);
  nor (_15644_, _15643_, _15638_);
  and (_15645_, _15644_, _05949_);
  and (_15646_, _04594_, _08322_);
  nor (_15647_, _15646_, _15625_);
  and (_15648_, _15647_, _03168_);
  and (_15649_, _15647_, _04505_);
  nor (_15650_, _04505_, _15637_);
  or (_15651_, _15650_, _15649_);
  and (_15652_, _15651_, _02662_);
  and (_15653_, _15627_, _02661_);
  or (_15654_, _15653_, _15652_);
  and (_15655_, _15654_, _03365_);
  nor (_15656_, _15644_, _03365_);
  nor (_15657_, _15656_, _15655_);
  nor (_15658_, _15657_, _03168_);
  or (_15659_, _15658_, _05949_);
  nor (_15660_, _15659_, _15648_);
  nor (_15661_, _15660_, _15645_);
  nor (_15662_, _15661_, _05959_);
  nor (_15663_, _15662_, _02024_);
  and (_15664_, _15663_, _15642_);
  and (_15665_, _08307_, _04594_);
  nor (_15666_, _15665_, _03139_);
  and (_15667_, _15666_, _15629_);
  nor (_15668_, _15667_, _15664_);
  nor (_15669_, _15668_, _06549_);
  nor (_15670_, _08185_, _06316_);
  nor (_15671_, _15670_, _05305_);
  and (_15672_, _04594_, _03016_);
  nor (_15673_, _15672_, _05245_);
  or (_15674_, _15673_, _15671_);
  and (_15675_, _15674_, _15629_);
  nor (_15676_, _15675_, _15669_);
  nor (_15677_, _15676_, _03251_);
  nor (_15678_, _15677_, _15635_);
  nor (_15679_, _15678_, _02669_);
  nor (_15680_, _15679_, _15632_);
  nor (_15681_, _15680_, _03243_);
  nor (_15682_, _15638_, _06122_);
  nor (_15683_, _15682_, _03244_);
  and (_15684_, _15683_, _15647_);
  nor (_15685_, _15684_, _15681_);
  nor (_15686_, _15685_, _03241_);
  and (_15687_, _15672_, _04835_);
  nor (_15688_, _15687_, _05357_);
  nand (_15689_, _15646_, _04835_);
  and (_15690_, _15689_, _03239_);
  or (_15691_, _15690_, _15688_);
  and (_15692_, _15691_, _15629_);
  or (_15693_, _15692_, _03123_);
  nor (_15694_, _15693_, _15686_);
  nor (_15695_, _15694_, _15628_);
  nor (_15696_, _15695_, _03121_);
  nor (_15697_, _15638_, _15626_);
  and (_15698_, _15697_, _03121_);
  nor (_15699_, _15698_, _15696_);
  or (_15700_, _15699_, _27789_);
  or (_15701_, _27788_, \oc8051_golden_model_1.TH1 [1]);
  and (_15702_, _15701_, _27053_);
  and (_28923_, _15702_, _15700_);
  not (_15703_, \oc8051_golden_model_1.TH1 [2]);
  nor (_15704_, _04594_, _15703_);
  and (_15705_, _04594_, _04170_);
  nor (_15706_, _15705_, _15704_);
  or (_15707_, _15706_, _05963_);
  and (_15708_, _04594_, \oc8051_golden_model_1.ACC [2]);
  nor (_15709_, _15708_, _15704_);
  nor (_15710_, _15709_, _05903_);
  nor (_15711_, _04505_, _15703_);
  or (_15712_, _15711_, _15710_);
  and (_15713_, _15712_, _02662_);
  nor (_15714_, _08420_, _06316_);
  nor (_15715_, _15714_, _15704_);
  nor (_15716_, _15715_, _02662_);
  or (_15717_, _15716_, _15713_);
  and (_15718_, _15717_, _03365_);
  nor (_15719_, _06316_, _03644_);
  nor (_15720_, _15719_, _15704_);
  nor (_15721_, _15720_, _03365_);
  nor (_15722_, _15721_, _15718_);
  nor (_15723_, _15722_, _03168_);
  nor (_15724_, _15709_, _03179_);
  nor (_15725_, _15724_, _05949_);
  not (_15726_, _15725_);
  nor (_15727_, _15726_, _15723_);
  and (_15728_, _15720_, _05949_);
  or (_15729_, _15728_, _05959_);
  or (_15730_, _15729_, _15727_);
  and (_15731_, _15730_, _03139_);
  and (_15732_, _15731_, _15707_);
  nor (_15733_, _08522_, _06316_);
  or (_15734_, _15704_, _03139_);
  nor (_15735_, _15734_, _15733_);
  or (_15736_, _15735_, _02575_);
  nor (_15737_, _15736_, _15732_);
  and (_15738_, _04594_, _06009_);
  nor (_15739_, _15738_, _15704_);
  nand (_15740_, _15739_, _05305_);
  and (_15741_, _15740_, _06549_);
  nor (_15742_, _15741_, _15737_);
  and (_15743_, _08537_, _04594_);
  nor (_15744_, _15743_, _15704_);
  and (_15745_, _15744_, _02656_);
  nor (_15746_, _15745_, _15742_);
  and (_15747_, _15746_, _03252_);
  and (_15748_, _08387_, _04594_);
  nor (_15749_, _15748_, _15704_);
  nor (_15750_, _15749_, _03252_);
  or (_15751_, _15750_, _15747_);
  and (_15752_, _15751_, _05332_);
  nor (_15753_, _15704_, _06121_);
  not (_15754_, _15753_);
  nor (_15755_, _15739_, _05332_);
  and (_15756_, _15755_, _15754_);
  nor (_15757_, _15756_, _15752_);
  nor (_15758_, _15757_, _03243_);
  or (_15759_, _15753_, _03244_);
  nor (_15760_, _15759_, _15709_);
  or (_15761_, _15760_, _02654_);
  nor (_15762_, _15761_, _15758_);
  nor (_15763_, _08536_, _06316_);
  nor (_15764_, _15763_, _15704_);
  and (_15765_, _15764_, _02654_);
  nor (_15766_, _15765_, _15762_);
  and (_15767_, _15766_, _05883_);
  nor (_15768_, _08386_, _06316_);
  nor (_15769_, _15768_, _15704_);
  nor (_15770_, _15769_, _05883_);
  or (_15771_, _15770_, _15767_);
  and (_15772_, _15771_, _03124_);
  nor (_15773_, _15715_, _03124_);
  or (_15774_, _15773_, _15772_);
  and (_15775_, _15774_, _03513_);
  and (_15776_, _08596_, _04594_);
  nor (_15777_, _15776_, _15704_);
  nor (_15778_, _15777_, _03513_);
  or (_15779_, _15778_, _15775_);
  or (_15780_, _15779_, _27789_);
  or (_15781_, _27788_, \oc8051_golden_model_1.TH1 [2]);
  and (_15782_, _15781_, _27053_);
  and (_28924_, _15782_, _15780_);
  not (_15783_, \oc8051_golden_model_1.TH1 [3]);
  nor (_15784_, _04594_, _15783_);
  and (_15785_, _04594_, \oc8051_golden_model_1.ACC [3]);
  nor (_15786_, _15785_, _15784_);
  nor (_15787_, _15786_, _05903_);
  nor (_15788_, _04505_, _15783_);
  or (_15789_, _15788_, _15787_);
  and (_15790_, _15789_, _02662_);
  nor (_15791_, _08646_, _06316_);
  nor (_15792_, _15791_, _15784_);
  nor (_15793_, _15792_, _02662_);
  or (_15794_, _15793_, _15790_);
  and (_15795_, _15794_, _03365_);
  nor (_15796_, _06316_, _03859_);
  nor (_15797_, _15796_, _15784_);
  nor (_15798_, _15797_, _03365_);
  nor (_15799_, _15798_, _15795_);
  nor (_15800_, _15799_, _03168_);
  nor (_15801_, _15786_, _03179_);
  nor (_15802_, _15801_, _05949_);
  not (_15803_, _15802_);
  nor (_15804_, _15803_, _15800_);
  and (_15805_, _15797_, _05949_);
  or (_15806_, _15805_, _05959_);
  or (_15807_, _15806_, _15804_);
  and (_15808_, _04594_, _04120_);
  nor (_15809_, _15808_, _15784_);
  or (_15810_, _15809_, _05963_);
  and (_15811_, _15810_, _03139_);
  and (_15812_, _15811_, _15807_);
  nor (_15813_, _08744_, _06316_);
  or (_15814_, _15784_, _03139_);
  nor (_15815_, _15814_, _15813_);
  or (_15816_, _15815_, _02575_);
  nor (_15817_, _15816_, _15812_);
  and (_15818_, _04594_, _05986_);
  nor (_15819_, _15818_, _15784_);
  nand (_15820_, _15819_, _05305_);
  and (_15821_, _15820_, _06549_);
  nor (_15822_, _15821_, _15817_);
  and (_15823_, _08622_, _04594_);
  nor (_15824_, _15823_, _15784_);
  and (_15825_, _15824_, _02656_);
  nor (_15826_, _15825_, _15822_);
  and (_15827_, _15826_, _03252_);
  and (_15828_, _08618_, _04594_);
  nor (_15829_, _15828_, _15784_);
  nor (_15830_, _15829_, _03252_);
  or (_15831_, _15830_, _15827_);
  and (_15832_, _15831_, _05332_);
  nor (_15833_, _15784_, _06120_);
  not (_15834_, _15833_);
  nor (_15835_, _15819_, _05332_);
  and (_15836_, _15835_, _15834_);
  nor (_15837_, _15836_, _15832_);
  nor (_15838_, _15837_, _03243_);
  or (_15839_, _15833_, _03244_);
  nor (_15840_, _15839_, _15786_);
  or (_15841_, _15840_, _02654_);
  nor (_15842_, _15841_, _15838_);
  nor (_15843_, _08621_, _06316_);
  nor (_15844_, _15843_, _15784_);
  and (_15845_, _15844_, _02654_);
  nor (_15846_, _15845_, _15842_);
  and (_15847_, _15846_, _05883_);
  nor (_15848_, _08617_, _06316_);
  nor (_15849_, _15848_, _15784_);
  nor (_15850_, _15849_, _05883_);
  or (_15851_, _15850_, _15847_);
  and (_15852_, _15851_, _03124_);
  nor (_15853_, _15792_, _03124_);
  or (_15854_, _15853_, _15852_);
  and (_15855_, _15854_, _03513_);
  and (_15856_, _08807_, _04594_);
  nor (_15857_, _15856_, _15784_);
  nor (_15858_, _15857_, _03513_);
  or (_15859_, _15858_, _15855_);
  or (_15860_, _15859_, _27789_);
  or (_15861_, _27788_, \oc8051_golden_model_1.TH1 [3]);
  and (_15862_, _15861_, _27053_);
  and (_28925_, _15862_, _15860_);
  not (_15863_, \oc8051_golden_model_1.TH1 [4]);
  nor (_15864_, _04594_, _15863_);
  and (_15865_, _08830_, _04594_);
  nor (_15866_, _15865_, _15864_);
  nor (_15867_, _15866_, _03252_);
  and (_15868_, _04594_, _05974_);
  nor (_15869_, _15868_, _15864_);
  and (_15870_, _15869_, _02575_);
  nor (_15871_, _06316_, _04325_);
  nor (_15872_, _15871_, _15864_);
  and (_15873_, _15872_, _05949_);
  and (_15874_, _04594_, \oc8051_golden_model_1.ACC [4]);
  nor (_15875_, _15874_, _15864_);
  nor (_15876_, _15875_, _05903_);
  nor (_15877_, _04505_, _15863_);
  or (_15878_, _15877_, _15876_);
  and (_15879_, _15878_, _02662_);
  nor (_15880_, _08838_, _06316_);
  nor (_15881_, _15880_, _15864_);
  nor (_15882_, _15881_, _02662_);
  or (_15883_, _15882_, _15879_);
  and (_15884_, _15883_, _03365_);
  nor (_15885_, _15872_, _03365_);
  nor (_15886_, _15885_, _15884_);
  nor (_15887_, _15886_, _03168_);
  nor (_15888_, _15875_, _03179_);
  nor (_15889_, _15888_, _05949_);
  not (_15890_, _15889_);
  nor (_15891_, _15890_, _15887_);
  nor (_15892_, _15891_, _15873_);
  nor (_15893_, _15892_, _05959_);
  and (_15894_, _04594_, _04012_);
  nor (_15895_, _15864_, _05963_);
  not (_15896_, _15895_);
  nor (_15897_, _15896_, _15894_);
  or (_15898_, _15897_, _02024_);
  nor (_15899_, _15898_, _15893_);
  nor (_15900_, _08967_, _06316_);
  nor (_15901_, _15900_, _15864_);
  nor (_15902_, _15901_, _03139_);
  or (_15903_, _15902_, _02575_);
  nor (_15904_, _15903_, _15899_);
  nor (_15905_, _15904_, _15870_);
  or (_15906_, _15905_, _02656_);
  and (_15907_, _08982_, _04594_);
  or (_15908_, _15907_, _15864_);
  or (_15909_, _15908_, _05305_);
  and (_15910_, _15909_, _03252_);
  and (_15911_, _15910_, _15906_);
  nor (_15912_, _15911_, _15867_);
  nor (_15913_, _15912_, _02669_);
  nor (_15914_, _15864_, _09034_);
  not (_15915_, _15914_);
  nor (_15916_, _15869_, _05332_);
  and (_15917_, _15916_, _15915_);
  nor (_15918_, _15917_, _15913_);
  nor (_15919_, _15918_, _03243_);
  or (_15920_, _15914_, _03244_);
  nor (_15921_, _15920_, _15875_);
  or (_15922_, _15921_, _02654_);
  nor (_15923_, _15922_, _15919_);
  nor (_15924_, _08981_, _06316_);
  nor (_15925_, _15924_, _15864_);
  and (_15926_, _15925_, _02654_);
  nor (_15927_, _15926_, _15923_);
  and (_15928_, _15927_, _05883_);
  nor (_15929_, _08828_, _06316_);
  nor (_15930_, _15929_, _15864_);
  nor (_15931_, _15930_, _05883_);
  or (_15932_, _15931_, _15928_);
  and (_15933_, _15932_, _03124_);
  nor (_15934_, _15881_, _03124_);
  or (_15935_, _15934_, _15933_);
  and (_15936_, _15935_, _03513_);
  and (_15937_, _09037_, _04594_);
  nor (_15938_, _15937_, _15864_);
  nor (_15939_, _15938_, _03513_);
  or (_15940_, _15939_, _15936_);
  or (_15941_, _15940_, _27789_);
  or (_15942_, _27788_, \oc8051_golden_model_1.TH1 [4]);
  and (_15943_, _15942_, _27053_);
  and (_28926_, _15943_, _15941_);
  not (_15944_, \oc8051_golden_model_1.TH1 [5]);
  nor (_15945_, _04594_, _15944_);
  and (_15946_, _09055_, _04594_);
  nor (_15947_, _15946_, _15945_);
  nor (_15948_, _15947_, _03252_);
  and (_15949_, _04594_, _06036_);
  nor (_15950_, _15949_, _15945_);
  and (_15951_, _15950_, _02575_);
  nor (_15952_, _06316_, _04480_);
  nor (_15953_, _15952_, _15945_);
  and (_15954_, _15953_, _05949_);
  and (_15955_, _04594_, \oc8051_golden_model_1.ACC [5]);
  nor (_15956_, _15955_, _15945_);
  nor (_15957_, _15956_, _03179_);
  nor (_15958_, _15956_, _05903_);
  nor (_15959_, _04505_, _15944_);
  or (_15960_, _15959_, _15958_);
  and (_15961_, _15960_, _02662_);
  nor (_15962_, _09087_, _06316_);
  nor (_15963_, _15962_, _15945_);
  nor (_15964_, _15963_, _02662_);
  or (_15965_, _15964_, _15961_);
  and (_15966_, _15965_, _03365_);
  nor (_15967_, _15953_, _03365_);
  nor (_15968_, _15967_, _15966_);
  nor (_15969_, _15968_, _03168_);
  or (_15970_, _15969_, _05949_);
  nor (_15971_, _15970_, _15957_);
  nor (_15972_, _15971_, _15954_);
  nor (_15973_, _15972_, _05959_);
  and (_15974_, _04594_, _03904_);
  nor (_15975_, _15945_, _05963_);
  not (_15976_, _15975_);
  nor (_15977_, _15976_, _15974_);
  or (_15978_, _15977_, _02024_);
  nor (_15979_, _15978_, _15973_);
  nor (_15980_, _09180_, _06316_);
  nor (_15981_, _15980_, _15945_);
  nor (_15982_, _15981_, _03139_);
  or (_15983_, _15982_, _02575_);
  nor (_15984_, _15983_, _15979_);
  nor (_15985_, _15984_, _15951_);
  or (_15986_, _15985_, _02656_);
  and (_15987_, _09195_, _04594_);
  or (_15988_, _15987_, _15945_);
  or (_15989_, _15988_, _05305_);
  and (_15990_, _15989_, _03252_);
  and (_15991_, _15990_, _15986_);
  nor (_15992_, _15991_, _15948_);
  nor (_15993_, _15992_, _02669_);
  not (_15994_, _15945_);
  and (_15995_, _15994_, _04787_);
  not (_15996_, _15995_);
  nor (_15997_, _15950_, _05332_);
  and (_15998_, _15997_, _15996_);
  nor (_15999_, _15998_, _15993_);
  nor (_16000_, _15999_, _03243_);
  or (_16001_, _15995_, _03244_);
  nor (_16002_, _16001_, _15956_);
  or (_16003_, _16002_, _02654_);
  nor (_16004_, _16003_, _16000_);
  nor (_16005_, _09194_, _06316_);
  nor (_16006_, _16005_, _15945_);
  and (_16007_, _16006_, _02654_);
  nor (_16008_, _16007_, _16004_);
  and (_16009_, _16008_, _05883_);
  nor (_16010_, _09054_, _06316_);
  nor (_16011_, _16010_, _15945_);
  nor (_16012_, _16011_, _05883_);
  or (_16013_, _16012_, _16009_);
  and (_16014_, _16013_, _03124_);
  nor (_16015_, _15963_, _03124_);
  or (_16016_, _16015_, _16014_);
  and (_16017_, _16016_, _03513_);
  and (_16018_, _09248_, _04594_);
  nor (_16019_, _16018_, _15945_);
  nor (_16020_, _16019_, _03513_);
  or (_16021_, _16020_, _16017_);
  or (_16022_, _16021_, _27789_);
  or (_16023_, _27788_, \oc8051_golden_model_1.TH1 [5]);
  and (_16024_, _16023_, _27053_);
  and (_28927_, _16024_, _16022_);
  not (_16025_, \oc8051_golden_model_1.TH1 [6]);
  nor (_16026_, _04594_, _16025_);
  and (_16027_, _09268_, _04594_);
  nor (_16028_, _16027_, _16026_);
  nor (_16029_, _16028_, _03252_);
  and (_16030_, _04594_, _03960_);
  or (_16031_, _16030_, _16026_);
  and (_16032_, _16031_, _05959_);
  and (_16033_, _04594_, \oc8051_golden_model_1.ACC [6]);
  nor (_16034_, _16033_, _16026_);
  nor (_16035_, _16034_, _05903_);
  nor (_16036_, _04505_, _16025_);
  or (_16037_, _16036_, _16035_);
  and (_16038_, _16037_, _02662_);
  nor (_16039_, _09301_, _06316_);
  nor (_16040_, _16039_, _16026_);
  nor (_16041_, _16040_, _02662_);
  or (_16042_, _16041_, _16038_);
  and (_16043_, _16042_, _03365_);
  nor (_16044_, _06316_, _04373_);
  nor (_16045_, _16044_, _16026_);
  nor (_16046_, _16045_, _03365_);
  nor (_16047_, _16046_, _16043_);
  nor (_16048_, _16047_, _03168_);
  nor (_16049_, _16034_, _03179_);
  nor (_16050_, _16049_, _05949_);
  not (_16051_, _16050_);
  nor (_16052_, _16051_, _16048_);
  and (_16053_, _16045_, _05949_);
  or (_16054_, _16053_, _05959_);
  nor (_16055_, _16054_, _16052_);
  or (_16056_, _16055_, _16032_);
  and (_16057_, _16056_, _03139_);
  and (_16058_, _09388_, _04594_);
  nor (_16059_, _16058_, _16026_);
  nor (_16060_, _16059_, _03139_);
  or (_16061_, _16060_, _06549_);
  or (_16062_, _16061_, _16057_);
  and (_16063_, _09404_, _04594_);
  or (_16064_, _16026_, _05305_);
  or (_16065_, _16064_, _16063_);
  and (_16066_, _04594_, _09395_);
  nor (_16067_, _16066_, _16026_);
  and (_16068_, _16067_, _02575_);
  nor (_16069_, _16068_, _03251_);
  and (_16070_, _16069_, _16065_);
  and (_16071_, _16070_, _16062_);
  nor (_16072_, _16071_, _16029_);
  nor (_16073_, _16072_, _02669_);
  nor (_16074_, _16026_, _06119_);
  not (_16075_, _16074_);
  nor (_16076_, _16067_, _05332_);
  and (_16077_, _16076_, _16075_);
  nor (_16078_, _16077_, _16073_);
  nor (_16079_, _16078_, _03243_);
  or (_16080_, _16074_, _03244_);
  nor (_16081_, _16080_, _16034_);
  or (_16082_, _16081_, _02654_);
  nor (_16083_, _16082_, _16079_);
  nor (_16084_, _09403_, _06316_);
  nor (_16085_, _16084_, _16026_);
  and (_16086_, _16085_, _02654_);
  nor (_16087_, _16086_, _16083_);
  and (_16088_, _16087_, _05883_);
  nor (_16089_, _09267_, _06316_);
  nor (_16090_, _16089_, _16026_);
  nor (_16091_, _16090_, _05883_);
  or (_16092_, _16091_, _16088_);
  and (_16093_, _16092_, _03124_);
  nor (_16094_, _16040_, _03124_);
  or (_16095_, _16094_, _16093_);
  and (_16096_, _16095_, _03513_);
  and (_16097_, _09456_, _04594_);
  nor (_16098_, _16097_, _16026_);
  nor (_16099_, _16098_, _03513_);
  or (_16100_, _16099_, _16096_);
  or (_16101_, _16100_, _27789_);
  or (_16102_, _27788_, \oc8051_golden_model_1.TH1 [6]);
  and (_16103_, _16102_, _27053_);
  and (_28928_, _16103_, _16101_);
  not (_16104_, \oc8051_golden_model_1.TL0 [0]);
  nor (_16105_, _04608_, _16104_);
  nor (_16106_, _04888_, _06226_);
  nor (_16107_, _16106_, _16105_);
  and (_16108_, _16107_, _11672_);
  and (_16109_, _04608_, \oc8051_golden_model_1.ACC [0]);
  nor (_16110_, _16109_, _16105_);
  nor (_16111_, _16110_, _03179_);
  nor (_16112_, _16110_, _05903_);
  nor (_16113_, _04505_, _16104_);
  or (_16114_, _16113_, _16112_);
  and (_16115_, _16114_, _02662_);
  nor (_16116_, _16107_, _02662_);
  or (_16117_, _16116_, _16115_);
  and (_16118_, _16117_, _03365_);
  and (_16119_, _04608_, _03716_);
  nor (_16120_, _16119_, _16105_);
  nor (_16121_, _16120_, _03365_);
  nor (_16122_, _16121_, _16118_);
  nor (_16123_, _16122_, _03168_);
  or (_16124_, _16123_, _05949_);
  nor (_16125_, _16124_, _16111_);
  and (_16126_, _16120_, _05949_);
  nor (_16127_, _16126_, _16125_);
  nor (_16128_, _16127_, _05959_);
  and (_16129_, _04608_, _04268_);
  nor (_16130_, _16105_, _05963_);
  not (_16131_, _16130_);
  nor (_16132_, _16131_, _16129_);
  nor (_16133_, _16132_, _16128_);
  nor (_16134_, _16133_, _02024_);
  nor (_16135_, _08093_, _06226_);
  or (_16136_, _16105_, _03139_);
  nor (_16137_, _16136_, _16135_);
  or (_16138_, _16137_, _02575_);
  nor (_16139_, _16138_, _16134_);
  and (_16140_, _04608_, _05996_);
  nor (_16141_, _16140_, _16105_);
  nand (_16142_, _16141_, _05305_);
  and (_16143_, _16142_, _06549_);
  nor (_16144_, _16143_, _16139_);
  and (_16145_, _07968_, _04608_);
  nor (_16146_, _16145_, _16105_);
  and (_16147_, _16146_, _02656_);
  nor (_16148_, _16147_, _16144_);
  and (_16149_, _16148_, _03252_);
  and (_16150_, _08110_, _04608_);
  nor (_16151_, _16150_, _16105_);
  nor (_16152_, _16151_, _03252_);
  or (_16153_, _16152_, _16149_);
  and (_16154_, _16153_, _05332_);
  or (_16155_, _16141_, _05332_);
  nor (_16156_, _16155_, _16106_);
  nor (_16157_, _16156_, _16154_);
  nor (_16158_, _16157_, _03243_);
  and (_16159_, _08108_, _04608_);
  or (_16160_, _16159_, _16105_);
  and (_16161_, _16160_, _03243_);
  or (_16162_, _16161_, _16158_);
  and (_16163_, _16162_, _05357_);
  nor (_16164_, _07967_, _06226_);
  nor (_16165_, _16164_, _16105_);
  nor (_16166_, _16165_, _05357_);
  or (_16167_, _16166_, _16163_);
  and (_16168_, _16167_, _05883_);
  nor (_16169_, _08109_, _06226_);
  nor (_16170_, _16169_, _16105_);
  nor (_16171_, _16170_, _05883_);
  nor (_16172_, _16171_, _11672_);
  not (_16173_, _16172_);
  nor (_16174_, _16173_, _16168_);
  nor (_16175_, _16174_, _16108_);
  or (_16176_, _16175_, _27789_);
  or (_16177_, _27788_, \oc8051_golden_model_1.TL0 [0]);
  and (_16178_, _16177_, _27053_);
  and (_28931_, _16178_, _16176_);
  nor (_16179_, _04608_, \oc8051_golden_model_1.TL0 [1]);
  and (_16180_, _08209_, _04608_);
  nor (_16181_, _16180_, _16179_);
  nor (_16182_, _16181_, _03124_);
  not (_16183_, _16179_);
  nor (_16184_, _08325_, _06226_);
  nor (_16185_, _16184_, _03252_);
  and (_16186_, _16185_, _16183_);
  and (_16187_, _04608_, _04218_);
  not (_16188_, \oc8051_golden_model_1.TL0 [1]);
  nor (_16189_, _04608_, _16188_);
  nor (_16190_, _16189_, _05963_);
  not (_16191_, _16190_);
  nor (_16192_, _16191_, _16187_);
  not (_16193_, _16192_);
  and (_16194_, _04608_, _08322_);
  nor (_16195_, _16194_, _16179_);
  and (_16196_, _16195_, _03168_);
  and (_16197_, _16195_, _04505_);
  nor (_16198_, _04505_, _16188_);
  or (_16199_, _16198_, _16197_);
  and (_16200_, _16199_, _02662_);
  and (_16201_, _16181_, _02661_);
  or (_16202_, _16201_, _16200_);
  and (_16203_, _16202_, _03365_);
  nor (_16204_, _06226_, _03777_);
  nor (_16205_, _16204_, _16189_);
  nor (_16206_, _16205_, _03365_);
  nor (_16207_, _16206_, _16203_);
  nor (_16208_, _16207_, _03168_);
  or (_16209_, _16208_, _05949_);
  nor (_16210_, _16209_, _16196_);
  and (_16211_, _16205_, _05949_);
  nor (_16212_, _16211_, _16210_);
  nor (_16213_, _16212_, _05959_);
  nor (_16214_, _16213_, _02024_);
  and (_16215_, _16214_, _16193_);
  and (_16216_, _08307_, _04608_);
  nor (_16217_, _16216_, _03139_);
  and (_16218_, _16217_, _16183_);
  nor (_16219_, _16218_, _16215_);
  nor (_16220_, _16219_, _06549_);
  nor (_16221_, _08185_, _06226_);
  nor (_16222_, _16221_, _05305_);
  and (_16223_, _04608_, _03016_);
  nor (_16224_, _16223_, _05245_);
  or (_16225_, _16224_, _16222_);
  and (_16226_, _16225_, _16183_);
  nor (_16227_, _16226_, _16220_);
  nor (_16228_, _16227_, _03251_);
  nor (_16229_, _16228_, _16186_);
  nor (_16230_, _16229_, _02669_);
  nor (_16231_, _08184_, _06226_);
  nor (_16232_, _16231_, _05332_);
  and (_16233_, _16232_, _16183_);
  nor (_16234_, _16233_, _16230_);
  nor (_16235_, _16234_, _03243_);
  nor (_16236_, _16189_, _06122_);
  nor (_16237_, _16236_, _03244_);
  and (_16238_, _16237_, _16195_);
  nor (_16239_, _16238_, _16235_);
  nor (_16240_, _16239_, _03241_);
  and (_16241_, _16223_, _04835_);
  nor (_16242_, _16241_, _05357_);
  and (_16243_, _16194_, _04835_);
  nor (_16244_, _16243_, _05883_);
  or (_16245_, _16244_, _16242_);
  and (_16246_, _16245_, _16183_);
  or (_16247_, _16246_, _03123_);
  nor (_16248_, _16247_, _16240_);
  nor (_16249_, _16248_, _16182_);
  nor (_16250_, _16249_, _03121_);
  nor (_16251_, _16189_, _16180_);
  and (_16252_, _16251_, _03121_);
  nor (_16253_, _16252_, _16250_);
  or (_16254_, _16253_, _27789_);
  or (_16255_, _27788_, \oc8051_golden_model_1.TL0 [1]);
  and (_16256_, _16255_, _27053_);
  and (_28932_, _16256_, _16254_);
  not (_16257_, \oc8051_golden_model_1.TL0 [2]);
  nor (_16258_, _04608_, _16257_);
  and (_16259_, _04608_, _04170_);
  nor (_16260_, _16259_, _16258_);
  or (_16261_, _16260_, _05963_);
  and (_16262_, _04608_, \oc8051_golden_model_1.ACC [2]);
  nor (_16263_, _16262_, _16258_);
  nor (_16264_, _16263_, _03179_);
  nor (_16265_, _16263_, _05903_);
  nor (_16266_, _04505_, _16257_);
  or (_16267_, _16266_, _16265_);
  and (_16268_, _16267_, _02662_);
  nor (_16269_, _08420_, _06226_);
  nor (_16270_, _16269_, _16258_);
  nor (_16271_, _16270_, _02662_);
  or (_16272_, _16271_, _16268_);
  and (_16273_, _16272_, _03365_);
  nor (_16274_, _06226_, _03644_);
  nor (_16275_, _16274_, _16258_);
  nor (_16276_, _16275_, _03365_);
  nor (_16277_, _16276_, _16273_);
  nor (_16278_, _16277_, _03168_);
  or (_16279_, _16278_, _05949_);
  nor (_16280_, _16279_, _16264_);
  and (_16281_, _16275_, _05949_);
  or (_16282_, _16281_, _05959_);
  or (_16283_, _16282_, _16280_);
  and (_16284_, _16283_, _03139_);
  and (_16285_, _16284_, _16261_);
  nor (_16286_, _08522_, _06226_);
  or (_16287_, _16258_, _03139_);
  nor (_16288_, _16287_, _16286_);
  or (_16289_, _16288_, _02575_);
  nor (_16290_, _16289_, _16285_);
  and (_16291_, _04608_, _06009_);
  nor (_16292_, _16291_, _16258_);
  nand (_16293_, _16292_, _05305_);
  and (_16294_, _16293_, _06549_);
  nor (_16295_, _16294_, _16290_);
  and (_16296_, _08537_, _04608_);
  nor (_16297_, _16296_, _16258_);
  and (_16298_, _16297_, _02656_);
  nor (_16299_, _16298_, _16295_);
  and (_16300_, _16299_, _03252_);
  and (_16301_, _08387_, _04608_);
  nor (_16302_, _16301_, _16258_);
  nor (_16303_, _16302_, _03252_);
  or (_16304_, _16303_, _16300_);
  and (_16305_, _16304_, _05332_);
  nor (_16306_, _16258_, _06121_);
  not (_16307_, _16306_);
  nor (_16308_, _16292_, _05332_);
  and (_16309_, _16308_, _16307_);
  nor (_16310_, _16309_, _16305_);
  nor (_16311_, _16310_, _03243_);
  or (_16312_, _16306_, _03244_);
  nor (_16313_, _16312_, _16263_);
  or (_16314_, _16313_, _02654_);
  nor (_16315_, _16314_, _16311_);
  nor (_16316_, _08536_, _06226_);
  nor (_16317_, _16316_, _16258_);
  and (_16318_, _16317_, _02654_);
  nor (_16319_, _16318_, _16315_);
  and (_16320_, _16319_, _05883_);
  nor (_16321_, _08386_, _06226_);
  nor (_16322_, _16321_, _16258_);
  nor (_16323_, _16322_, _05883_);
  or (_16324_, _16323_, _16320_);
  and (_16325_, _16324_, _03124_);
  nor (_16326_, _16270_, _03124_);
  or (_16327_, _16326_, _16325_);
  and (_16328_, _16327_, _03513_);
  and (_16329_, _08596_, _04608_);
  nor (_16330_, _16329_, _16258_);
  nor (_16331_, _16330_, _03513_);
  or (_16332_, _16331_, _16328_);
  or (_16333_, _16332_, _27789_);
  or (_16334_, _27788_, \oc8051_golden_model_1.TL0 [2]);
  and (_16335_, _16334_, _27053_);
  and (_28933_, _16335_, _16333_);
  not (_16336_, \oc8051_golden_model_1.TL0 [3]);
  nor (_16337_, _04608_, _16336_);
  and (_16338_, _08618_, _04608_);
  nor (_16339_, _16338_, _16337_);
  nor (_16340_, _16339_, _03252_);
  and (_16341_, _04608_, _04120_);
  or (_16342_, _16341_, _16337_);
  and (_16343_, _16342_, _05959_);
  and (_16344_, _04608_, \oc8051_golden_model_1.ACC [3]);
  nor (_16345_, _16344_, _16337_);
  nor (_16346_, _16345_, _03179_);
  nor (_16347_, _16345_, _05903_);
  nor (_16348_, _04505_, _16336_);
  or (_16349_, _16348_, _16347_);
  and (_16350_, _16349_, _02662_);
  nor (_16351_, _08646_, _06226_);
  nor (_16352_, _16351_, _16337_);
  nor (_16353_, _16352_, _02662_);
  or (_16354_, _16353_, _16350_);
  and (_16355_, _16354_, _03365_);
  nor (_16356_, _06226_, _03859_);
  nor (_16357_, _16356_, _16337_);
  nor (_16358_, _16357_, _03365_);
  nor (_16359_, _16358_, _16355_);
  nor (_16360_, _16359_, _03168_);
  or (_16361_, _16360_, _05949_);
  nor (_16362_, _16361_, _16346_);
  and (_16363_, _16357_, _05949_);
  or (_16364_, _16363_, _05959_);
  nor (_16365_, _16364_, _16362_);
  or (_16366_, _16365_, _16343_);
  and (_16367_, _16366_, _03139_);
  nor (_16368_, _08744_, _06226_);
  nor (_16369_, _16368_, _16337_);
  nor (_16370_, _16369_, _03139_);
  or (_16371_, _16370_, _06549_);
  or (_16372_, _16371_, _16367_);
  and (_16373_, _08622_, _04608_);
  or (_16374_, _16337_, _05305_);
  or (_16375_, _16374_, _16373_);
  and (_16376_, _04608_, _05986_);
  nor (_16377_, _16376_, _16337_);
  and (_16378_, _16377_, _02575_);
  nor (_16379_, _16378_, _03251_);
  and (_16380_, _16379_, _16375_);
  and (_16381_, _16380_, _16372_);
  nor (_16382_, _16381_, _16340_);
  nor (_16383_, _16382_, _02669_);
  nor (_16384_, _16337_, _06120_);
  not (_16385_, _16384_);
  nor (_16386_, _16377_, _05332_);
  and (_16387_, _16386_, _16385_);
  nor (_16388_, _16387_, _16383_);
  nor (_16389_, _16388_, _03243_);
  or (_16390_, _16384_, _03244_);
  nor (_16391_, _16390_, _16345_);
  or (_16392_, _16391_, _02654_);
  nor (_16393_, _16392_, _16389_);
  nor (_16394_, _08621_, _06226_);
  nor (_16395_, _16394_, _16337_);
  and (_16396_, _16395_, _02654_);
  nor (_16397_, _16396_, _16393_);
  and (_16398_, _16397_, _05883_);
  nor (_16399_, _08617_, _06226_);
  nor (_16400_, _16399_, _16337_);
  nor (_16401_, _16400_, _05883_);
  or (_16402_, _16401_, _16398_);
  and (_16403_, _16402_, _03124_);
  nor (_16404_, _16352_, _03124_);
  or (_16405_, _16404_, _16403_);
  and (_16406_, _16405_, _03513_);
  and (_16407_, _08807_, _04608_);
  nor (_16408_, _16407_, _16337_);
  nor (_16409_, _16408_, _03513_);
  or (_16410_, _16409_, _16406_);
  or (_16411_, _16410_, _27789_);
  or (_16412_, _27788_, \oc8051_golden_model_1.TL0 [3]);
  and (_16413_, _16412_, _27053_);
  and (_28934_, _16413_, _16411_);
  not (_16414_, \oc8051_golden_model_1.TL0 [4]);
  nor (_16415_, _04608_, _16414_);
  and (_16416_, _08830_, _04608_);
  nor (_16417_, _16416_, _16415_);
  nor (_16418_, _16417_, _03252_);
  and (_16419_, _04608_, _05974_);
  nor (_16420_, _16419_, _16415_);
  and (_16421_, _16420_, _02575_);
  nor (_16422_, _06226_, _04325_);
  nor (_16423_, _16422_, _16415_);
  and (_16424_, _16423_, _05949_);
  and (_16425_, _04608_, \oc8051_golden_model_1.ACC [4]);
  nor (_16426_, _16425_, _16415_);
  nor (_16427_, _16426_, _05903_);
  nor (_16428_, _04505_, _16414_);
  or (_16429_, _16428_, _16427_);
  and (_16430_, _16429_, _02662_);
  nor (_16431_, _08838_, _06226_);
  nor (_16432_, _16431_, _16415_);
  nor (_16433_, _16432_, _02662_);
  or (_16434_, _16433_, _16430_);
  and (_16435_, _16434_, _03365_);
  nor (_16436_, _16423_, _03365_);
  nor (_16437_, _16436_, _16435_);
  nor (_16438_, _16437_, _03168_);
  nor (_16439_, _16426_, _03179_);
  nor (_16440_, _16439_, _05949_);
  not (_16441_, _16440_);
  nor (_16442_, _16441_, _16438_);
  nor (_16443_, _16442_, _16424_);
  nor (_16444_, _16443_, _05959_);
  and (_16445_, _04608_, _04012_);
  nor (_16446_, _16415_, _05963_);
  not (_16447_, _16446_);
  nor (_16448_, _16447_, _16445_);
  or (_16449_, _16448_, _02024_);
  nor (_16450_, _16449_, _16444_);
  nor (_16451_, _08967_, _06226_);
  nor (_16452_, _16451_, _16415_);
  nor (_16453_, _16452_, _03139_);
  or (_16454_, _16453_, _02575_);
  nor (_16455_, _16454_, _16450_);
  nor (_16456_, _16455_, _16421_);
  or (_16457_, _16456_, _02656_);
  and (_16458_, _08982_, _04608_);
  or (_16459_, _16458_, _16415_);
  or (_16460_, _16459_, _05305_);
  and (_16461_, _16460_, _03252_);
  and (_16462_, _16461_, _16457_);
  nor (_16463_, _16462_, _16418_);
  nor (_16464_, _16463_, _02669_);
  nor (_16465_, _16415_, _09034_);
  not (_16466_, _16465_);
  nor (_16467_, _16420_, _05332_);
  and (_16468_, _16467_, _16466_);
  nor (_16469_, _16468_, _16464_);
  nor (_16470_, _16469_, _03243_);
  or (_16471_, _16465_, _03244_);
  nor (_16472_, _16471_, _16426_);
  or (_16473_, _16472_, _02654_);
  nor (_16474_, _16473_, _16470_);
  nor (_16475_, _08981_, _06226_);
  nor (_16476_, _16475_, _16415_);
  and (_16477_, _16476_, _02654_);
  nor (_16478_, _16477_, _16474_);
  and (_16479_, _16478_, _05883_);
  nor (_16480_, _08828_, _06226_);
  nor (_16481_, _16480_, _16415_);
  nor (_16482_, _16481_, _05883_);
  or (_16483_, _16482_, _16479_);
  and (_16484_, _16483_, _03124_);
  nor (_16485_, _16432_, _03124_);
  or (_16486_, _16485_, _16484_);
  and (_16487_, _16486_, _03513_);
  and (_16488_, _09037_, _04608_);
  nor (_16489_, _16488_, _16415_);
  nor (_16490_, _16489_, _03513_);
  or (_16491_, _16490_, _16487_);
  or (_16492_, _16491_, _27789_);
  or (_16493_, _27788_, \oc8051_golden_model_1.TL0 [4]);
  and (_16494_, _16493_, _27053_);
  and (_28935_, _16494_, _16492_);
  not (_16495_, \oc8051_golden_model_1.TL0 [5]);
  nor (_16496_, _04608_, _16495_);
  not (_16497_, _16496_);
  and (_16498_, _16497_, _04787_);
  not (_16499_, _16498_);
  and (_16500_, _04608_, _06036_);
  nor (_16501_, _16500_, _16496_);
  nor (_16502_, _16501_, _05332_);
  and (_16503_, _16502_, _16499_);
  and (_16504_, _09055_, _04608_);
  nor (_16505_, _16504_, _16496_);
  nor (_16506_, _16505_, _03252_);
  nor (_16507_, _09180_, _06226_);
  or (_16508_, _16496_, _03139_);
  or (_16509_, _16508_, _16507_);
  nor (_16510_, _09087_, _06226_);
  nor (_16511_, _16510_, _16496_);
  nor (_16512_, _16511_, _02662_);
  nor (_16513_, _04505_, _16495_);
  and (_16514_, _04608_, \oc8051_golden_model_1.ACC [5]);
  nor (_16515_, _16514_, _16496_);
  nor (_16516_, _16515_, _05903_);
  nor (_16517_, _16516_, _16513_);
  nor (_16518_, _16517_, _02661_);
  or (_16519_, _16518_, _16512_);
  and (_16520_, _16519_, _03365_);
  nor (_16521_, _06226_, _04480_);
  nor (_16522_, _16521_, _16496_);
  nor (_16523_, _16522_, _03365_);
  or (_16524_, _16523_, _16520_);
  and (_16525_, _16524_, _03179_);
  nor (_16526_, _16515_, _03179_);
  nor (_16527_, _16526_, _05949_);
  not (_16528_, _16527_);
  nor (_16529_, _16528_, _16525_);
  and (_16530_, _16522_, _05949_);
  or (_16531_, _16530_, _05959_);
  nor (_16532_, _16531_, _16529_);
  and (_16533_, _04608_, _03904_);
  or (_16534_, _16533_, _16496_);
  and (_16535_, _16534_, _05959_);
  or (_16536_, _16535_, _02024_);
  or (_16537_, _16536_, _16532_);
  and (_16538_, _16537_, _16509_);
  and (_16539_, _16538_, _05245_);
  nor (_16540_, _16501_, _05245_);
  or (_16541_, _16540_, _16539_);
  or (_16542_, _16541_, _02656_);
  and (_16543_, _09195_, _04608_);
  or (_16544_, _16543_, _16496_);
  or (_16545_, _16544_, _05305_);
  and (_16546_, _16545_, _03252_);
  and (_16547_, _16546_, _16542_);
  nor (_16548_, _16547_, _16506_);
  nor (_16549_, _16548_, _02669_);
  nor (_16550_, _16549_, _16503_);
  nor (_16551_, _16550_, _03243_);
  or (_16552_, _16498_, _03244_);
  nor (_16553_, _16552_, _16515_);
  or (_16554_, _16553_, _02654_);
  nor (_16555_, _16554_, _16551_);
  nor (_16556_, _09194_, _06226_);
  nor (_16557_, _16556_, _16496_);
  and (_16558_, _16557_, _02654_);
  nor (_16559_, _16558_, _16555_);
  and (_16560_, _16559_, _05883_);
  nor (_16561_, _09054_, _06226_);
  nor (_16562_, _16561_, _16496_);
  nor (_16563_, _16562_, _05883_);
  or (_16564_, _16563_, _16560_);
  and (_16565_, _16564_, _03124_);
  nor (_16566_, _16511_, _03124_);
  or (_16567_, _16566_, _16565_);
  and (_16568_, _16567_, _03513_);
  and (_16569_, _09248_, _04608_);
  nor (_16570_, _16569_, _16496_);
  nor (_16571_, _16570_, _03513_);
  or (_16572_, _16571_, _16568_);
  or (_16573_, _16572_, _27789_);
  or (_16574_, _27788_, \oc8051_golden_model_1.TL0 [5]);
  and (_16575_, _16574_, _27053_);
  and (_28936_, _16575_, _16573_);
  not (_16576_, \oc8051_golden_model_1.TL0 [6]);
  nor (_16577_, _04608_, _16576_);
  nor (_16578_, _16577_, _06119_);
  not (_16579_, _16578_);
  and (_16580_, _04608_, _09395_);
  nor (_16581_, _16580_, _16577_);
  nor (_16582_, _16581_, _05332_);
  and (_16583_, _16582_, _16579_);
  and (_16584_, _09268_, _04608_);
  nor (_16585_, _16584_, _16577_);
  nor (_16586_, _16585_, _03252_);
  and (_16587_, _04608_, _03960_);
  or (_16588_, _16587_, _16577_);
  and (_16589_, _16588_, _05959_);
  and (_16590_, _04608_, \oc8051_golden_model_1.ACC [6]);
  nor (_16591_, _16590_, _16577_);
  nor (_16592_, _16591_, _03179_);
  nor (_16593_, _16591_, _05903_);
  nor (_16594_, _04505_, _16576_);
  or (_16595_, _16594_, _16593_);
  and (_16596_, _16595_, _02662_);
  nor (_16597_, _09301_, _06226_);
  nor (_16598_, _16597_, _16577_);
  nor (_16599_, _16598_, _02662_);
  or (_16600_, _16599_, _16596_);
  and (_16601_, _16600_, _03365_);
  nor (_16602_, _06226_, _04373_);
  nor (_16603_, _16602_, _16577_);
  nor (_16604_, _16603_, _03365_);
  nor (_16605_, _16604_, _16601_);
  nor (_16606_, _16605_, _03168_);
  or (_16607_, _16606_, _05949_);
  nor (_16608_, _16607_, _16592_);
  and (_16609_, _16603_, _05949_);
  or (_16610_, _16609_, _05959_);
  nor (_16611_, _16610_, _16608_);
  or (_16612_, _16611_, _16589_);
  and (_16613_, _16612_, _03139_);
  and (_16614_, _09388_, _04608_);
  nor (_16615_, _16614_, _16577_);
  nor (_16616_, _16615_, _03139_);
  or (_16617_, _16616_, _06549_);
  or (_16618_, _16617_, _16613_);
  and (_16619_, _09404_, _04608_);
  or (_16620_, _16577_, _05305_);
  or (_16621_, _16620_, _16619_);
  and (_16622_, _16581_, _02575_);
  nor (_16623_, _16622_, _03251_);
  and (_16624_, _16623_, _16621_);
  and (_16625_, _16624_, _16618_);
  nor (_16626_, _16625_, _16586_);
  nor (_16627_, _16626_, _02669_);
  nor (_16628_, _16627_, _16583_);
  nor (_16629_, _16628_, _03243_);
  or (_16630_, _16578_, _03244_);
  nor (_16631_, _16630_, _16591_);
  or (_16632_, _16631_, _02654_);
  nor (_16633_, _16632_, _16629_);
  nor (_16634_, _09403_, _06226_);
  nor (_16635_, _16634_, _16577_);
  and (_16636_, _16635_, _02654_);
  nor (_16637_, _16636_, _16633_);
  and (_16638_, _16637_, _05883_);
  nor (_16639_, _09267_, _06226_);
  nor (_16640_, _16639_, _16577_);
  nor (_16641_, _16640_, _05883_);
  or (_16642_, _16641_, _16638_);
  and (_16643_, _16642_, _03124_);
  nor (_16644_, _16598_, _03124_);
  or (_16645_, _16644_, _16643_);
  and (_16646_, _16645_, _03513_);
  and (_16647_, _09456_, _04608_);
  nor (_16648_, _16647_, _16577_);
  nor (_16649_, _16648_, _03513_);
  or (_16650_, _16649_, _16646_);
  or (_16651_, _16650_, _27789_);
  or (_16652_, _27788_, \oc8051_golden_model_1.TL0 [6]);
  and (_16653_, _16652_, _27053_);
  and (_28937_, _16653_, _16651_);
  not (_16654_, \oc8051_golden_model_1.TL1 [0]);
  nor (_16655_, _04590_, _16654_);
  nor (_16656_, _04888_, _06151_);
  nor (_16657_, _16656_, _16655_);
  and (_16658_, _16657_, _11672_);
  and (_16659_, _04590_, _03716_);
  nor (_16660_, _16659_, _16655_);
  and (_16661_, _16660_, _05949_);
  and (_16662_, _04590_, \oc8051_golden_model_1.ACC [0]);
  nor (_16663_, _16662_, _16655_);
  nor (_16664_, _16663_, _03179_);
  nor (_16665_, _16663_, _05903_);
  nor (_16666_, _04505_, _16654_);
  or (_16667_, _16666_, _16665_);
  and (_16668_, _16667_, _02662_);
  nor (_16669_, _16657_, _02662_);
  or (_16670_, _16669_, _16668_);
  and (_16671_, _16670_, _03365_);
  nor (_16672_, _16660_, _03365_);
  nor (_16673_, _16672_, _16671_);
  nor (_16674_, _16673_, _03168_);
  or (_16675_, _16674_, _05949_);
  nor (_16676_, _16675_, _16664_);
  nor (_16677_, _16676_, _16661_);
  nor (_16678_, _16677_, _05959_);
  and (_16679_, _04590_, _04268_);
  nor (_16680_, _16655_, _05963_);
  not (_16681_, _16680_);
  nor (_16682_, _16681_, _16679_);
  nor (_16683_, _16682_, _16678_);
  nor (_16684_, _16683_, _02024_);
  nor (_16685_, _08093_, _06151_);
  or (_16686_, _16655_, _03139_);
  nor (_16687_, _16686_, _16685_);
  or (_16688_, _16687_, _02575_);
  nor (_16689_, _16688_, _16684_);
  and (_16690_, _04590_, _05996_);
  nor (_16691_, _16690_, _16655_);
  nand (_16692_, _16691_, _05305_);
  and (_16693_, _16692_, _06549_);
  nor (_16694_, _16693_, _16689_);
  and (_16695_, _07968_, _04590_);
  nor (_16696_, _16695_, _16655_);
  and (_16697_, _16696_, _02656_);
  nor (_16698_, _16697_, _16694_);
  and (_16699_, _16698_, _03252_);
  and (_16700_, _08110_, _04590_);
  nor (_16701_, _16700_, _16655_);
  nor (_16702_, _16701_, _03252_);
  or (_16703_, _16702_, _16699_);
  and (_16704_, _16703_, _05332_);
  or (_16705_, _16691_, _05332_);
  nor (_16706_, _16705_, _16656_);
  nor (_16707_, _16706_, _16704_);
  nor (_16708_, _16707_, _03243_);
  and (_16709_, _08108_, _04590_);
  or (_16710_, _16709_, _16655_);
  and (_16711_, _16710_, _03243_);
  or (_16712_, _16711_, _16708_);
  and (_16713_, _16712_, _05357_);
  nor (_16714_, _07967_, _06151_);
  nor (_16715_, _16714_, _16655_);
  nor (_16716_, _16715_, _05357_);
  or (_16717_, _16716_, _16713_);
  and (_16718_, _16717_, _05883_);
  nor (_16719_, _08109_, _06151_);
  nor (_16720_, _16719_, _16655_);
  nor (_16721_, _16720_, _05883_);
  nor (_16722_, _16721_, _11672_);
  not (_16723_, _16722_);
  nor (_16724_, _16723_, _16718_);
  nor (_16725_, _16724_, _16658_);
  or (_16726_, _16725_, _27789_);
  or (_16727_, _27788_, \oc8051_golden_model_1.TL1 [0]);
  and (_16728_, _16727_, _27053_);
  and (_28940_, _16728_, _16726_);
  nor (_16729_, _04590_, \oc8051_golden_model_1.TL1 [1]);
  and (_16730_, _08209_, _04590_);
  nor (_16731_, _16730_, _16729_);
  nor (_16732_, _16731_, _03124_);
  not (_16733_, _16729_);
  nor (_16734_, _08325_, _06151_);
  nor (_16735_, _16734_, _03252_);
  and (_16736_, _16735_, _16733_);
  and (_16737_, _04590_, _04218_);
  not (_16738_, \oc8051_golden_model_1.TL1 [1]);
  nor (_16739_, _04590_, _16738_);
  nor (_16740_, _16739_, _05963_);
  not (_16741_, _16740_);
  nor (_16742_, _16741_, _16737_);
  not (_16743_, _16742_);
  and (_16744_, _04590_, _08322_);
  nor (_16745_, _16744_, _16729_);
  and (_16746_, _16745_, _03168_);
  and (_16747_, _16745_, _04505_);
  nor (_16748_, _04505_, _16738_);
  or (_16749_, _16748_, _16747_);
  and (_16750_, _16749_, _02662_);
  and (_16751_, _16731_, _02661_);
  or (_16752_, _16751_, _16750_);
  and (_16753_, _16752_, _03365_);
  nor (_16754_, _06151_, _03777_);
  nor (_16755_, _16754_, _16739_);
  nor (_16756_, _16755_, _03365_);
  nor (_16757_, _16756_, _16753_);
  nor (_16758_, _16757_, _03168_);
  or (_16759_, _16758_, _05949_);
  nor (_16760_, _16759_, _16746_);
  and (_16761_, _16755_, _05949_);
  nor (_16762_, _16761_, _16760_);
  nor (_16763_, _16762_, _05959_);
  nor (_16764_, _16763_, _02024_);
  and (_16765_, _16764_, _16743_);
  and (_16766_, _08307_, _04590_);
  nor (_16767_, _16766_, _03139_);
  and (_16768_, _16767_, _16733_);
  nor (_16769_, _16768_, _16765_);
  nor (_16770_, _16769_, _06549_);
  nor (_16771_, _08185_, _06151_);
  nor (_16772_, _16771_, _05305_);
  and (_16773_, _04590_, _03016_);
  nor (_16774_, _16773_, _05245_);
  or (_16775_, _16774_, _16772_);
  and (_16776_, _16775_, _16733_);
  nor (_16777_, _16776_, _16770_);
  nor (_16778_, _16777_, _03251_);
  nor (_16779_, _16778_, _16736_);
  nor (_16780_, _16779_, _02669_);
  nor (_16781_, _08184_, _06151_);
  nor (_16782_, _16781_, _05332_);
  and (_16783_, _16782_, _16733_);
  nor (_16784_, _16783_, _16780_);
  nor (_16785_, _16784_, _03243_);
  nor (_16786_, _16739_, _06122_);
  nor (_16787_, _16786_, _03244_);
  and (_16788_, _16787_, _16745_);
  nor (_16789_, _16788_, _16785_);
  nor (_16790_, _16789_, _03241_);
  and (_16791_, _16773_, _04835_);
  nor (_16792_, _16791_, _05357_);
  nand (_16793_, _16744_, _04835_);
  and (_16794_, _16793_, _03239_);
  or (_16795_, _16794_, _16792_);
  and (_16796_, _16795_, _16733_);
  or (_16797_, _16796_, _03123_);
  nor (_16798_, _16797_, _16790_);
  nor (_16799_, _16798_, _16732_);
  nor (_16800_, _16799_, _03121_);
  nor (_16801_, _16739_, _16730_);
  and (_16802_, _16801_, _03121_);
  nor (_16803_, _16802_, _16800_);
  or (_16804_, _16803_, _27789_);
  or (_16805_, _27788_, \oc8051_golden_model_1.TL1 [1]);
  and (_16806_, _16805_, _27053_);
  and (_28941_, _16806_, _16804_);
  not (_16807_, \oc8051_golden_model_1.TL1 [2]);
  nor (_16808_, _04590_, _16807_);
  nor (_16809_, _16808_, _06121_);
  not (_16810_, _16809_);
  and (_16811_, _04590_, _06009_);
  nor (_16812_, _16811_, _16808_);
  nor (_16813_, _16812_, _05332_);
  and (_16814_, _16813_, _16810_);
  and (_16815_, _04590_, _04170_);
  nor (_16816_, _16815_, _16808_);
  or (_16817_, _16816_, _05963_);
  and (_16818_, _04590_, \oc8051_golden_model_1.ACC [2]);
  nor (_16819_, _16818_, _16808_);
  nor (_16820_, _16819_, _05903_);
  nor (_16821_, _04505_, _16807_);
  or (_16822_, _16821_, _16820_);
  and (_16823_, _16822_, _02662_);
  nor (_16824_, _08420_, _06151_);
  nor (_16825_, _16824_, _16808_);
  nor (_16826_, _16825_, _02662_);
  or (_16827_, _16826_, _16823_);
  and (_16828_, _16827_, _03365_);
  nor (_16829_, _06151_, _03644_);
  nor (_16830_, _16829_, _16808_);
  nor (_16831_, _16830_, _03365_);
  nor (_16832_, _16831_, _16828_);
  nor (_16833_, _16832_, _03168_);
  nor (_16834_, _16819_, _03179_);
  nor (_16835_, _16834_, _05949_);
  not (_16836_, _16835_);
  nor (_16837_, _16836_, _16833_);
  and (_16838_, _16830_, _05949_);
  or (_16839_, _16838_, _05959_);
  or (_16840_, _16839_, _16837_);
  and (_16841_, _16840_, _03139_);
  and (_16842_, _16841_, _16817_);
  nor (_16843_, _08522_, _06151_);
  or (_16844_, _16808_, _03139_);
  nor (_16845_, _16844_, _16843_);
  or (_16846_, _16845_, _02575_);
  nor (_16847_, _16846_, _16842_);
  nand (_16848_, _16812_, _05305_);
  and (_16849_, _16848_, _06549_);
  nor (_16850_, _16849_, _16847_);
  and (_16851_, _08537_, _04590_);
  nor (_16852_, _16851_, _16808_);
  and (_16853_, _16852_, _02656_);
  nor (_16854_, _16853_, _16850_);
  and (_16855_, _16854_, _03252_);
  and (_16856_, _08387_, _04590_);
  nor (_16857_, _16856_, _16808_);
  nor (_16858_, _16857_, _03252_);
  or (_16859_, _16858_, _16855_);
  and (_16860_, _16859_, _05332_);
  nor (_16861_, _16860_, _16814_);
  nor (_16862_, _16861_, _03243_);
  or (_16863_, _16809_, _03244_);
  nor (_16864_, _16863_, _16819_);
  or (_16865_, _16864_, _02654_);
  nor (_16866_, _16865_, _16862_);
  nor (_16867_, _08536_, _06151_);
  nor (_16868_, _16867_, _16808_);
  and (_16869_, _16868_, _02654_);
  nor (_16870_, _16869_, _16866_);
  and (_16871_, _16870_, _05883_);
  nor (_16872_, _08386_, _06151_);
  nor (_16873_, _16872_, _16808_);
  nor (_16874_, _16873_, _05883_);
  or (_16875_, _16874_, _16871_);
  and (_16876_, _16875_, _03124_);
  nor (_16877_, _16825_, _03124_);
  or (_16878_, _16877_, _16876_);
  and (_16879_, _16878_, _03513_);
  and (_16880_, _08596_, _04590_);
  nor (_16881_, _16880_, _16808_);
  nor (_16882_, _16881_, _03513_);
  or (_16884_, _16882_, _16879_);
  or (_16885_, _16884_, _27789_);
  or (_16886_, _27788_, \oc8051_golden_model_1.TL1 [2]);
  and (_16887_, _16886_, _27053_);
  and (_28942_, _16887_, _16885_);
  not (_16888_, \oc8051_golden_model_1.TL1 [3]);
  nor (_16889_, _04590_, _16888_);
  nor (_16890_, _16889_, _06120_);
  not (_16891_, _16890_);
  and (_16892_, _04590_, _05986_);
  nor (_16894_, _16892_, _16889_);
  nor (_16895_, _16894_, _05332_);
  and (_16896_, _16895_, _16891_);
  and (_16897_, _08618_, _04590_);
  nor (_16898_, _16897_, _16889_);
  nor (_16899_, _16898_, _03252_);
  and (_16900_, _04590_, _04120_);
  or (_16901_, _16900_, _16889_);
  and (_16902_, _16901_, _05959_);
  and (_16903_, _04590_, \oc8051_golden_model_1.ACC [3]);
  nor (_16905_, _16903_, _16889_);
  nor (_16906_, _16905_, _03179_);
  nor (_16907_, _16905_, _05903_);
  nor (_16908_, _04505_, _16888_);
  or (_16909_, _16908_, _16907_);
  and (_16910_, _16909_, _02662_);
  nor (_16911_, _08646_, _06151_);
  nor (_16912_, _16911_, _16889_);
  nor (_16913_, _16912_, _02662_);
  or (_16914_, _16913_, _16910_);
  and (_16916_, _16914_, _03365_);
  nor (_16917_, _06151_, _03859_);
  nor (_16918_, _16917_, _16889_);
  nor (_16919_, _16918_, _03365_);
  nor (_16920_, _16919_, _16916_);
  nor (_16921_, _16920_, _03168_);
  or (_16922_, _16921_, _05949_);
  nor (_16923_, _16922_, _16906_);
  and (_16924_, _16918_, _05949_);
  or (_16925_, _16924_, _05959_);
  nor (_16927_, _16925_, _16923_);
  or (_16928_, _16927_, _16902_);
  and (_16929_, _16928_, _03139_);
  nor (_16930_, _08744_, _06151_);
  nor (_16931_, _16930_, _16889_);
  nor (_16932_, _16931_, _03139_);
  or (_16933_, _16932_, _06549_);
  or (_16934_, _16933_, _16929_);
  and (_16935_, _08622_, _04590_);
  or (_16936_, _16889_, _05305_);
  or (_16938_, _16936_, _16935_);
  and (_16939_, _16894_, _02575_);
  nor (_16940_, _16939_, _03251_);
  and (_16941_, _16940_, _16938_);
  and (_16942_, _16941_, _16934_);
  nor (_16943_, _16942_, _16899_);
  nor (_16944_, _16943_, _02669_);
  nor (_16945_, _16944_, _16896_);
  nor (_16946_, _16945_, _03243_);
  or (_16947_, _16890_, _03244_);
  nor (_16949_, _16947_, _16905_);
  or (_16950_, _16949_, _02654_);
  nor (_16951_, _16950_, _16946_);
  nor (_16952_, _08621_, _06151_);
  nor (_16953_, _16952_, _16889_);
  and (_16954_, _16953_, _02654_);
  nor (_16955_, _16954_, _16951_);
  and (_16956_, _16955_, _05883_);
  nor (_16957_, _08617_, _06151_);
  nor (_16958_, _16957_, _16889_);
  nor (_16960_, _16958_, _05883_);
  or (_16961_, _16960_, _16956_);
  and (_16962_, _16961_, _03124_);
  nor (_16963_, _16912_, _03124_);
  or (_16964_, _16963_, _16962_);
  and (_16965_, _16964_, _03513_);
  and (_16966_, _08807_, _04590_);
  nor (_16967_, _16966_, _16889_);
  nor (_16968_, _16967_, _03513_);
  or (_16969_, _16968_, _16965_);
  or (_16971_, _16969_, _27789_);
  or (_16972_, _27788_, \oc8051_golden_model_1.TL1 [3]);
  and (_16973_, _16972_, _27053_);
  and (_28943_, _16973_, _16971_);
  not (_16974_, \oc8051_golden_model_1.TL1 [4]);
  nor (_16975_, _04590_, _16974_);
  and (_16976_, _08830_, _04590_);
  nor (_16977_, _16976_, _16975_);
  nor (_16978_, _16977_, _03252_);
  and (_16979_, _04590_, _05974_);
  nor (_16981_, _16979_, _16975_);
  and (_16982_, _16981_, _02575_);
  nor (_16983_, _06151_, _04325_);
  nor (_16984_, _16983_, _16975_);
  and (_16985_, _16984_, _05949_);
  and (_16986_, _04590_, \oc8051_golden_model_1.ACC [4]);
  nor (_16987_, _16986_, _16975_);
  nor (_16988_, _16987_, _05903_);
  nor (_16989_, _04505_, _16974_);
  or (_16990_, _16989_, _16988_);
  and (_16992_, _16990_, _02662_);
  nor (_16993_, _08838_, _06151_);
  nor (_16994_, _16993_, _16975_);
  nor (_16995_, _16994_, _02662_);
  or (_16996_, _16995_, _16992_);
  and (_16997_, _16996_, _03365_);
  nor (_16998_, _16984_, _03365_);
  nor (_16999_, _16998_, _16997_);
  nor (_17000_, _16999_, _03168_);
  nor (_17001_, _16987_, _03179_);
  nor (_17003_, _17001_, _05949_);
  not (_17004_, _17003_);
  nor (_17005_, _17004_, _17000_);
  nor (_17006_, _17005_, _16985_);
  nor (_17007_, _17006_, _05959_);
  and (_17008_, _04590_, _04012_);
  nor (_17009_, _16975_, _05963_);
  not (_17010_, _17009_);
  nor (_17011_, _17010_, _17008_);
  or (_17012_, _17011_, _02024_);
  nor (_17014_, _17012_, _17007_);
  nor (_17015_, _08967_, _06151_);
  nor (_17016_, _17015_, _16975_);
  nor (_17017_, _17016_, _03139_);
  or (_17018_, _17017_, _02575_);
  nor (_17019_, _17018_, _17014_);
  nor (_17020_, _17019_, _16982_);
  or (_17021_, _17020_, _02656_);
  and (_17022_, _08982_, _04590_);
  or (_17023_, _17022_, _16975_);
  or (_17025_, _17023_, _05305_);
  and (_17026_, _17025_, _03252_);
  and (_17027_, _17026_, _17021_);
  nor (_17028_, _17027_, _16978_);
  nor (_17029_, _17028_, _02669_);
  nor (_17030_, _16975_, _09034_);
  not (_17031_, _17030_);
  nor (_17032_, _16981_, _05332_);
  and (_17033_, _17032_, _17031_);
  nor (_17034_, _17033_, _17029_);
  nor (_17036_, _17034_, _03243_);
  or (_17037_, _17030_, _03244_);
  nor (_17038_, _17037_, _16987_);
  or (_17039_, _17038_, _02654_);
  nor (_17040_, _17039_, _17036_);
  nor (_17041_, _08981_, _06151_);
  nor (_17042_, _17041_, _16975_);
  and (_17043_, _17042_, _02654_);
  nor (_17044_, _17043_, _17040_);
  and (_17045_, _17044_, _05883_);
  nor (_17047_, _08828_, _06151_);
  nor (_17048_, _17047_, _16975_);
  nor (_17049_, _17048_, _05883_);
  or (_17050_, _17049_, _17045_);
  and (_17051_, _17050_, _03124_);
  nor (_17052_, _16994_, _03124_);
  or (_17053_, _17052_, _17051_);
  and (_17054_, _17053_, _03513_);
  and (_17055_, _09037_, _04590_);
  nor (_17056_, _17055_, _16975_);
  nor (_17058_, _17056_, _03513_);
  or (_17059_, _17058_, _17054_);
  or (_17060_, _17059_, _27789_);
  or (_17061_, _27788_, \oc8051_golden_model_1.TL1 [4]);
  and (_17062_, _17061_, _27053_);
  and (_28944_, _17062_, _17060_);
  not (_17063_, \oc8051_golden_model_1.TL1 [5]);
  nor (_17064_, _04590_, _17063_);
  and (_17065_, _09055_, _04590_);
  nor (_17066_, _17065_, _17064_);
  nor (_17068_, _17066_, _03252_);
  and (_17069_, _04590_, _06036_);
  nor (_17070_, _17069_, _17064_);
  and (_17071_, _17070_, _02575_);
  nor (_17072_, _06151_, _04480_);
  nor (_17073_, _17072_, _17064_);
  and (_17074_, _17073_, _05949_);
  and (_17075_, _04590_, \oc8051_golden_model_1.ACC [5]);
  nor (_17076_, _17075_, _17064_);
  nor (_17077_, _17076_, _03179_);
  nor (_17079_, _17076_, _05903_);
  nor (_17080_, _04505_, _17063_);
  or (_17081_, _17080_, _17079_);
  and (_17082_, _17081_, _02662_);
  nor (_17083_, _09087_, _06151_);
  nor (_17084_, _17083_, _17064_);
  nor (_17085_, _17084_, _02662_);
  or (_17086_, _17085_, _17082_);
  and (_17087_, _17086_, _03365_);
  nor (_17088_, _17073_, _03365_);
  nor (_17090_, _17088_, _17087_);
  nor (_17091_, _17090_, _03168_);
  or (_17092_, _17091_, _05949_);
  nor (_17093_, _17092_, _17077_);
  nor (_17094_, _17093_, _17074_);
  nor (_17095_, _17094_, _05959_);
  and (_17096_, _04590_, _03904_);
  nor (_17097_, _17064_, _05963_);
  not (_17098_, _17097_);
  nor (_17099_, _17098_, _17096_);
  or (_17101_, _17099_, _02024_);
  nor (_17102_, _17101_, _17095_);
  nor (_17103_, _09180_, _06151_);
  nor (_17104_, _17103_, _17064_);
  nor (_17105_, _17104_, _03139_);
  or (_17106_, _17105_, _02575_);
  nor (_17107_, _17106_, _17102_);
  nor (_17108_, _17107_, _17071_);
  or (_17109_, _17108_, _02656_);
  and (_17110_, _09195_, _04590_);
  or (_17112_, _17110_, _17064_);
  or (_17113_, _17112_, _05305_);
  and (_17114_, _17113_, _03252_);
  and (_17115_, _17114_, _17109_);
  nor (_17116_, _17115_, _17068_);
  nor (_17117_, _17116_, _02669_);
  not (_17118_, _17064_);
  and (_17119_, _17118_, _04787_);
  not (_17120_, _17119_);
  nor (_17121_, _17070_, _05332_);
  and (_17123_, _17121_, _17120_);
  nor (_17124_, _17123_, _17117_);
  nor (_17125_, _17124_, _03243_);
  or (_17126_, _17119_, _03244_);
  nor (_17127_, _17126_, _17076_);
  or (_17128_, _17127_, _02654_);
  nor (_17129_, _17128_, _17125_);
  nor (_17130_, _09194_, _06151_);
  nor (_17131_, _17130_, _17064_);
  and (_17132_, _17131_, _02654_);
  nor (_17134_, _17132_, _17129_);
  and (_17135_, _17134_, _05883_);
  nor (_17136_, _09054_, _06151_);
  nor (_17137_, _17136_, _17064_);
  nor (_17138_, _17137_, _05883_);
  or (_17139_, _17138_, _17135_);
  and (_17140_, _17139_, _03124_);
  nor (_17141_, _17084_, _03124_);
  or (_17142_, _17141_, _17140_);
  and (_17143_, _17142_, _03513_);
  and (_17145_, _09248_, _04590_);
  nor (_17146_, _17145_, _17064_);
  nor (_17147_, _17146_, _03513_);
  or (_17148_, _17147_, _17143_);
  or (_17149_, _17148_, _27789_);
  or (_17150_, _27788_, \oc8051_golden_model_1.TL1 [5]);
  and (_17151_, _17150_, _27053_);
  and (_28945_, _17151_, _17149_);
  not (_17152_, \oc8051_golden_model_1.TL1 [6]);
  nor (_17153_, _04590_, _17152_);
  and (_17155_, _09268_, _04590_);
  nor (_17156_, _17155_, _17153_);
  nor (_17157_, _17156_, _03252_);
  and (_17158_, _04590_, _03960_);
  or (_17159_, _17158_, _17153_);
  and (_17160_, _17159_, _05959_);
  and (_17161_, _04590_, \oc8051_golden_model_1.ACC [6]);
  nor (_17162_, _17161_, _17153_);
  nor (_17163_, _17162_, _03179_);
  nor (_17164_, _17162_, _05903_);
  nor (_17166_, _04505_, _17152_);
  or (_17167_, _17166_, _17164_);
  and (_17168_, _17167_, _02662_);
  nor (_17169_, _09301_, _06151_);
  nor (_17170_, _17169_, _17153_);
  nor (_17171_, _17170_, _02662_);
  or (_17172_, _17171_, _17168_);
  and (_17173_, _17172_, _03365_);
  nor (_17174_, _06151_, _04373_);
  nor (_17175_, _17174_, _17153_);
  nor (_17177_, _17175_, _03365_);
  nor (_17178_, _17177_, _17173_);
  nor (_17179_, _17178_, _03168_);
  or (_17180_, _17179_, _05949_);
  nor (_17181_, _17180_, _17163_);
  and (_17182_, _17175_, _05949_);
  or (_17183_, _17182_, _05959_);
  nor (_17184_, _17183_, _17181_);
  or (_17185_, _17184_, _17160_);
  and (_17186_, _17185_, _03139_);
  and (_17188_, _09388_, _04590_);
  nor (_17189_, _17188_, _17153_);
  nor (_17190_, _17189_, _03139_);
  or (_17191_, _17190_, _06549_);
  or (_17192_, _17191_, _17186_);
  and (_17193_, _09404_, _04590_);
  or (_17194_, _17153_, _05305_);
  or (_17195_, _17194_, _17193_);
  and (_17196_, _04590_, _09395_);
  nor (_17197_, _17196_, _17153_);
  and (_17199_, _17197_, _02575_);
  nor (_17200_, _17199_, _03251_);
  and (_17201_, _17200_, _17195_);
  and (_17202_, _17201_, _17192_);
  nor (_17203_, _17202_, _17157_);
  nor (_17204_, _17203_, _02669_);
  nor (_17205_, _17153_, _06119_);
  not (_17206_, _17205_);
  nor (_17207_, _17197_, _05332_);
  and (_17208_, _17207_, _17206_);
  nor (_17210_, _17208_, _17204_);
  nor (_17211_, _17210_, _03243_);
  or (_17212_, _17205_, _03244_);
  nor (_17213_, _17212_, _17162_);
  or (_17214_, _17213_, _02654_);
  nor (_17215_, _17214_, _17211_);
  nor (_17216_, _09403_, _06151_);
  nor (_17217_, _17216_, _17153_);
  and (_17218_, _17217_, _02654_);
  nor (_17219_, _17218_, _17215_);
  and (_17221_, _17219_, _05883_);
  nor (_17222_, _09267_, _06151_);
  nor (_17223_, _17222_, _17153_);
  nor (_17224_, _17223_, _05883_);
  or (_17225_, _17224_, _17221_);
  and (_17226_, _17225_, _03124_);
  nor (_17227_, _17170_, _03124_);
  or (_17228_, _17227_, _17226_);
  and (_17229_, _17228_, _03513_);
  and (_17230_, _09456_, _04590_);
  nor (_17232_, _17230_, _17153_);
  nor (_17233_, _17232_, _03513_);
  or (_17234_, _17233_, _17229_);
  or (_17235_, _17234_, _27789_);
  or (_17236_, _27788_, \oc8051_golden_model_1.TL1 [6]);
  and (_17237_, _17236_, _27053_);
  and (_28946_, _17237_, _17235_);
  not (_17238_, \oc8051_golden_model_1.TMOD [0]);
  nor (_17239_, _04605_, _17238_);
  nor (_17240_, _04888_, _05913_);
  nor (_17242_, _17240_, _17239_);
  and (_17243_, _17242_, _11672_);
  and (_17244_, _04605_, _05996_);
  nor (_17245_, _17244_, _17239_);
  nor (_17246_, _17245_, _05332_);
  not (_17247_, _17246_);
  nor (_17248_, _17247_, _17240_);
  and (_17249_, _04605_, \oc8051_golden_model_1.ACC [0]);
  nor (_17250_, _17249_, _17239_);
  nor (_17251_, _17250_, _03179_);
  nor (_17253_, _17251_, _05949_);
  nor (_17254_, _17242_, _02662_);
  nor (_17255_, _04505_, _17238_);
  nor (_17256_, _17250_, _05903_);
  nor (_17257_, _17256_, _17255_);
  nor (_17258_, _17257_, _02661_);
  or (_17259_, _17258_, _03162_);
  nor (_17260_, _17259_, _17254_);
  or (_17261_, _17260_, _03168_);
  and (_17262_, _17261_, _17253_);
  and (_17264_, _04605_, _03716_);
  or (_17265_, _17239_, _12270_);
  nor (_17266_, _17265_, _17264_);
  nor (_17267_, _17266_, _17262_);
  nor (_17268_, _17267_, _05959_);
  and (_17269_, _04605_, _04268_);
  nor (_17270_, _17239_, _05963_);
  not (_17271_, _17270_);
  nor (_17272_, _17271_, _17269_);
  nor (_17273_, _17272_, _17268_);
  nor (_17275_, _17273_, _02024_);
  nor (_17276_, _08093_, _05913_);
  or (_17277_, _17239_, _03139_);
  nor (_17278_, _17277_, _17276_);
  or (_17279_, _17278_, _02575_);
  nor (_17280_, _17279_, _17275_);
  nor (_17281_, _17245_, _05245_);
  or (_17282_, _17281_, _17280_);
  and (_17283_, _17282_, _05305_);
  and (_17284_, _07968_, _04605_);
  nor (_17286_, _17284_, _17239_);
  nor (_17287_, _17286_, _05305_);
  or (_17288_, _17287_, _17283_);
  and (_17289_, _17288_, _03252_);
  and (_17290_, _08110_, _04605_);
  nor (_17291_, _17290_, _17239_);
  nor (_17292_, _17291_, _03252_);
  or (_17293_, _17292_, _17289_);
  and (_17294_, _17293_, _05332_);
  nor (_17295_, _17294_, _17248_);
  nor (_17297_, _17295_, _03243_);
  and (_17298_, _08108_, _04605_);
  or (_17299_, _17298_, _17239_);
  and (_17300_, _17299_, _03243_);
  or (_17301_, _17300_, _17297_);
  and (_17302_, _17301_, _05357_);
  nor (_17303_, _07967_, _05913_);
  nor (_17304_, _17303_, _17239_);
  nor (_17305_, _17304_, _05357_);
  or (_17306_, _17305_, _17302_);
  and (_17308_, _17306_, _05883_);
  nor (_17309_, _08109_, _05913_);
  nor (_17310_, _17309_, _17239_);
  nor (_17311_, _17310_, _05883_);
  nor (_17312_, _17311_, _11672_);
  not (_17313_, _17312_);
  nor (_17314_, _17313_, _17308_);
  nor (_17315_, _17314_, _17243_);
  or (_17316_, _17315_, _27789_);
  or (_17317_, _27788_, \oc8051_golden_model_1.TMOD [0]);
  and (_17319_, _17317_, _27053_);
  and (_28949_, _17319_, _17316_);
  nor (_17320_, _04605_, \oc8051_golden_model_1.TMOD [1]);
  and (_17321_, _08209_, _04605_);
  nor (_17322_, _17321_, _17320_);
  nor (_17323_, _17322_, _03124_);
  not (_17324_, _17320_);
  nor (_17325_, _08325_, _05913_);
  nor (_17326_, _17325_, _03252_);
  and (_17327_, _17326_, _17324_);
  and (_17329_, _04605_, _04218_);
  not (_17330_, \oc8051_golden_model_1.TMOD [1]);
  nor (_17331_, _04605_, _17330_);
  nor (_17332_, _17331_, _05963_);
  not (_17333_, _17332_);
  nor (_17334_, _17333_, _17329_);
  not (_17335_, _17334_);
  nor (_17336_, _05913_, _03777_);
  nor (_17337_, _17336_, _17331_);
  and (_17338_, _17337_, _05949_);
  and (_17340_, _04605_, _08322_);
  nor (_17341_, _17340_, _17320_);
  and (_17342_, _17341_, _04505_);
  nor (_17343_, _04505_, _17330_);
  or (_17344_, _17343_, _17342_);
  and (_17345_, _17344_, _02662_);
  and (_17346_, _17322_, _02661_);
  or (_17347_, _17346_, _17345_);
  and (_17348_, _17347_, _03365_);
  nor (_17349_, _17337_, _03365_);
  nor (_17351_, _17349_, _17348_);
  nor (_17352_, _17351_, _03168_);
  and (_17353_, _17341_, _03168_);
  nor (_17354_, _17353_, _05949_);
  not (_17355_, _17354_);
  nor (_17356_, _17355_, _17352_);
  nor (_17357_, _17356_, _17338_);
  nor (_17358_, _17357_, _05959_);
  nor (_17359_, _17358_, _02024_);
  and (_17360_, _17359_, _17335_);
  and (_17362_, _08307_, _04605_);
  nor (_17363_, _17362_, _03139_);
  and (_17364_, _17363_, _17324_);
  nor (_17365_, _17364_, _17360_);
  nor (_17366_, _17365_, _06549_);
  nor (_17367_, _08185_, _05913_);
  nor (_17368_, _17367_, _05305_);
  and (_17369_, _04605_, _03016_);
  nor (_17370_, _17369_, _05245_);
  or (_17371_, _17370_, _17368_);
  and (_17373_, _17371_, _17324_);
  nor (_17374_, _17373_, _17366_);
  nor (_17375_, _17374_, _03251_);
  nor (_17376_, _17375_, _17327_);
  nor (_17377_, _17376_, _02669_);
  nor (_17378_, _08184_, _05913_);
  nor (_17379_, _17378_, _05332_);
  and (_17380_, _17379_, _17324_);
  nor (_17381_, _17380_, _17377_);
  nor (_17382_, _17381_, _03243_);
  nor (_17384_, _17331_, _06122_);
  nor (_17385_, _17384_, _03244_);
  and (_17386_, _17385_, _17341_);
  nor (_17387_, _17386_, _17382_);
  nor (_17388_, _17387_, _03241_);
  and (_17389_, _17369_, _04835_);
  nor (_17390_, _17389_, _05357_);
  nand (_17391_, _17340_, _04835_);
  and (_17392_, _17391_, _03239_);
  or (_17393_, _17392_, _17390_);
  and (_17395_, _17393_, _17324_);
  or (_17396_, _17395_, _03123_);
  nor (_17397_, _17396_, _17388_);
  nor (_17398_, _17397_, _17323_);
  nor (_17399_, _17398_, _03121_);
  nor (_17400_, _17331_, _17321_);
  and (_17401_, _17400_, _03121_);
  nor (_17402_, _17401_, _17399_);
  or (_17403_, _17402_, _27789_);
  or (_17404_, _27788_, \oc8051_golden_model_1.TMOD [1]);
  and (_17406_, _17404_, _27053_);
  and (_28950_, _17406_, _17403_);
  not (_17407_, \oc8051_golden_model_1.TMOD [2]);
  nor (_17408_, _04605_, _17407_);
  and (_17409_, _04605_, _04170_);
  nor (_17410_, _17409_, _17408_);
  or (_17411_, _17410_, _05963_);
  and (_17412_, _04605_, \oc8051_golden_model_1.ACC [2]);
  nor (_17413_, _17412_, _17408_);
  nor (_17414_, _17413_, _05903_);
  nor (_17416_, _04505_, _17407_);
  or (_17417_, _17416_, _17414_);
  and (_17418_, _17417_, _02662_);
  nor (_17419_, _08420_, _05913_);
  nor (_17420_, _17419_, _17408_);
  nor (_17421_, _17420_, _02662_);
  or (_17422_, _17421_, _17418_);
  and (_17423_, _17422_, _03365_);
  nor (_17424_, _05913_, _03644_);
  nor (_17425_, _17424_, _17408_);
  nor (_17427_, _17425_, _03365_);
  nor (_17428_, _17427_, _17423_);
  nor (_17429_, _17428_, _03168_);
  nor (_17430_, _17413_, _03179_);
  nor (_17431_, _17430_, _05949_);
  not (_17432_, _17431_);
  nor (_17433_, _17432_, _17429_);
  and (_17434_, _17425_, _05949_);
  or (_17435_, _17434_, _05959_);
  or (_17436_, _17435_, _17433_);
  and (_17438_, _17436_, _03139_);
  and (_17439_, _17438_, _17411_);
  nor (_17440_, _08522_, _05913_);
  or (_17441_, _17408_, _03139_);
  nor (_17442_, _17441_, _17440_);
  or (_17443_, _17442_, _02575_);
  nor (_17444_, _17443_, _17439_);
  and (_17445_, _04605_, _06009_);
  nor (_17446_, _17445_, _17408_);
  nor (_17447_, _17446_, _05245_);
  or (_17449_, _17447_, _17444_);
  and (_17450_, _17449_, _05305_);
  and (_17451_, _08537_, _04605_);
  nor (_17452_, _17451_, _17408_);
  nor (_17453_, _17452_, _05305_);
  or (_17454_, _17453_, _17450_);
  and (_17455_, _17454_, _03252_);
  and (_17456_, _08387_, _04605_);
  nor (_17457_, _17456_, _17408_);
  nor (_17458_, _17457_, _03252_);
  or (_17459_, _17458_, _17455_);
  and (_17460_, _17459_, _05332_);
  nor (_17461_, _17408_, _06121_);
  or (_17462_, _17446_, _05332_);
  nor (_17463_, _17462_, _17461_);
  nor (_17464_, _17463_, _17460_);
  nor (_17465_, _17464_, _03243_);
  or (_17466_, _17461_, _03244_);
  nor (_17467_, _17466_, _17413_);
  or (_17468_, _17467_, _02654_);
  nor (_17471_, _17468_, _17465_);
  nor (_17472_, _08536_, _05913_);
  nor (_17473_, _17472_, _17408_);
  and (_17474_, _17473_, _02654_);
  nor (_17475_, _17474_, _17471_);
  and (_17476_, _17475_, _05883_);
  nor (_17477_, _08386_, _05913_);
  nor (_17478_, _17477_, _17408_);
  nor (_17479_, _17478_, _05883_);
  or (_17480_, _17479_, _17476_);
  and (_17482_, _17480_, _03124_);
  nor (_17483_, _17420_, _03124_);
  or (_17484_, _17483_, _17482_);
  and (_17485_, _17484_, _03513_);
  and (_17486_, _08596_, _04605_);
  nor (_17487_, _17486_, _17408_);
  nor (_17488_, _17487_, _03513_);
  or (_17489_, _17488_, _17485_);
  or (_17490_, _17489_, _27789_);
  or (_17491_, _27788_, \oc8051_golden_model_1.TMOD [2]);
  and (_17493_, _17491_, _27053_);
  and (_28951_, _17493_, _17490_);
  not (_17494_, \oc8051_golden_model_1.TMOD [3]);
  nor (_17495_, _04605_, _17494_);
  and (_17496_, _08618_, _04605_);
  nor (_17497_, _17496_, _17495_);
  nor (_17498_, _17497_, _03252_);
  and (_17499_, _04605_, _04120_);
  or (_17500_, _17499_, _17495_);
  and (_17501_, _17500_, _05959_);
  and (_17503_, _04605_, \oc8051_golden_model_1.ACC [3]);
  nor (_17504_, _17503_, _17495_);
  nor (_17505_, _17504_, _03179_);
  nor (_17506_, _17504_, _05903_);
  nor (_17507_, _04505_, _17494_);
  or (_17508_, _17507_, _17506_);
  and (_17509_, _17508_, _02662_);
  nor (_17510_, _08646_, _05913_);
  nor (_17511_, _17510_, _17495_);
  nor (_17512_, _17511_, _02662_);
  or (_17514_, _17512_, _17509_);
  and (_17515_, _17514_, _03365_);
  nor (_17516_, _05913_, _03859_);
  nor (_17517_, _17516_, _17495_);
  nor (_17518_, _17517_, _03365_);
  nor (_17519_, _17518_, _17515_);
  nor (_17520_, _17519_, _03168_);
  or (_17521_, _17520_, _05949_);
  nor (_17522_, _17521_, _17505_);
  and (_17523_, _17517_, _05949_);
  or (_17525_, _17523_, _05959_);
  nor (_17526_, _17525_, _17522_);
  or (_17527_, _17526_, _17501_);
  and (_17528_, _17527_, _03139_);
  nor (_17529_, _08744_, _05913_);
  nor (_17530_, _17529_, _17495_);
  nor (_17531_, _17530_, _03139_);
  or (_17532_, _17531_, _06549_);
  or (_17533_, _17532_, _17528_);
  and (_17534_, _08622_, _04605_);
  or (_17536_, _17495_, _05305_);
  or (_17537_, _17536_, _17534_);
  and (_17538_, _04605_, _05986_);
  nor (_17539_, _17538_, _17495_);
  and (_17540_, _17539_, _02575_);
  nor (_17541_, _17540_, _03251_);
  and (_17542_, _17541_, _17537_);
  and (_17543_, _17542_, _17533_);
  nor (_17544_, _17543_, _17498_);
  nor (_17545_, _17544_, _02669_);
  nor (_17547_, _17495_, _06120_);
  not (_17548_, _17547_);
  nor (_17549_, _17539_, _05332_);
  and (_17550_, _17549_, _17548_);
  nor (_17551_, _17550_, _17545_);
  nor (_17552_, _17551_, _03243_);
  or (_17553_, _17547_, _03244_);
  nor (_17554_, _17553_, _17504_);
  or (_17555_, _17554_, _02654_);
  nor (_17556_, _17555_, _17552_);
  nor (_17558_, _08621_, _05913_);
  nor (_17559_, _17558_, _17495_);
  and (_17560_, _17559_, _02654_);
  nor (_17561_, _17560_, _17556_);
  and (_17562_, _17561_, _05883_);
  nor (_17563_, _08617_, _05913_);
  nor (_17564_, _17563_, _17495_);
  nor (_17565_, _17564_, _05883_);
  or (_17566_, _17565_, _17562_);
  and (_17567_, _17566_, _03124_);
  nor (_17569_, _17511_, _03124_);
  or (_17570_, _17569_, _17567_);
  and (_17571_, _17570_, _03513_);
  and (_17572_, _08807_, _04605_);
  nor (_17573_, _17572_, _17495_);
  nor (_17574_, _17573_, _03513_);
  or (_17575_, _17574_, _17571_);
  or (_17576_, _17575_, _27789_);
  or (_17577_, _27788_, \oc8051_golden_model_1.TMOD [3]);
  and (_17578_, _17577_, _27053_);
  and (_28952_, _17578_, _17576_);
  not (_17580_, \oc8051_golden_model_1.TMOD [4]);
  nor (_17581_, _04605_, _17580_);
  and (_17582_, _08830_, _04605_);
  nor (_17583_, _17582_, _17581_);
  nor (_17584_, _17583_, _03252_);
  and (_17585_, _04605_, _05974_);
  nor (_17586_, _17585_, _17581_);
  and (_17587_, _17586_, _02575_);
  nor (_17588_, _05913_, _04325_);
  nor (_17590_, _17588_, _17581_);
  and (_17591_, _17590_, _05949_);
  and (_17592_, _04605_, \oc8051_golden_model_1.ACC [4]);
  nor (_17593_, _17592_, _17581_);
  nor (_17594_, _17593_, _03179_);
  nor (_17595_, _17593_, _05903_);
  nor (_17596_, _04505_, _17580_);
  or (_17597_, _17596_, _17595_);
  and (_17598_, _17597_, _02662_);
  nor (_17599_, _08838_, _05913_);
  nor (_17601_, _17599_, _17581_);
  nor (_17602_, _17601_, _02662_);
  or (_17603_, _17602_, _17598_);
  and (_17604_, _17603_, _03365_);
  nor (_17605_, _17590_, _03365_);
  nor (_17606_, _17605_, _17604_);
  nor (_17607_, _17606_, _03168_);
  or (_17608_, _17607_, _05949_);
  nor (_17609_, _17608_, _17594_);
  nor (_17610_, _17609_, _17591_);
  nor (_17612_, _17610_, _05959_);
  and (_17613_, _04605_, _04012_);
  nor (_17614_, _17581_, _05963_);
  not (_17615_, _17614_);
  nor (_17616_, _17615_, _17613_);
  or (_17617_, _17616_, _02024_);
  nor (_17618_, _17617_, _17612_);
  nor (_17619_, _08967_, _05913_);
  nor (_17620_, _17619_, _17581_);
  nor (_17621_, _17620_, _03139_);
  or (_17623_, _17621_, _02575_);
  nor (_17624_, _17623_, _17618_);
  nor (_17625_, _17624_, _17587_);
  or (_17626_, _17625_, _02656_);
  and (_17627_, _08982_, _04605_);
  or (_17628_, _17627_, _17581_);
  or (_17629_, _17628_, _05305_);
  and (_17630_, _17629_, _03252_);
  and (_17631_, _17630_, _17626_);
  nor (_17632_, _17631_, _17584_);
  nor (_17634_, _17632_, _02669_);
  nor (_17635_, _17581_, _09034_);
  not (_17636_, _17635_);
  nor (_17637_, _17586_, _05332_);
  and (_17638_, _17637_, _17636_);
  nor (_17639_, _17638_, _17634_);
  nor (_17640_, _17639_, _03243_);
  or (_17641_, _17635_, _03244_);
  nor (_17642_, _17641_, _17593_);
  or (_17643_, _17642_, _02654_);
  nor (_17645_, _17643_, _17640_);
  nor (_17646_, _08981_, _05913_);
  nor (_17647_, _17646_, _17581_);
  and (_17648_, _17647_, _02654_);
  nor (_17649_, _17648_, _17645_);
  and (_17650_, _17649_, _05883_);
  nor (_17651_, _08828_, _05913_);
  nor (_17652_, _17651_, _17581_);
  nor (_17653_, _17652_, _05883_);
  or (_17654_, _17653_, _17650_);
  and (_17656_, _17654_, _03124_);
  nor (_17657_, _17601_, _03124_);
  or (_17658_, _17657_, _17656_);
  and (_17659_, _17658_, _03513_);
  and (_17660_, _09037_, _04605_);
  nor (_17661_, _17660_, _17581_);
  nor (_17662_, _17661_, _03513_);
  or (_17663_, _17662_, _17659_);
  or (_17664_, _17663_, _27789_);
  or (_17665_, _27788_, \oc8051_golden_model_1.TMOD [4]);
  and (_17667_, _17665_, _27053_);
  and (_28953_, _17667_, _17664_);
  not (_17668_, \oc8051_golden_model_1.TMOD [5]);
  nor (_17669_, _04605_, _17668_);
  and (_17670_, _09055_, _04605_);
  nor (_17671_, _17670_, _17669_);
  nor (_17672_, _17671_, _03252_);
  and (_17673_, _04605_, _06036_);
  nor (_17674_, _17673_, _17669_);
  and (_17675_, _17674_, _02575_);
  and (_17677_, _04605_, \oc8051_golden_model_1.ACC [5]);
  nor (_17678_, _17677_, _17669_);
  nor (_17679_, _17678_, _03179_);
  nor (_17680_, _17678_, _05903_);
  nor (_17681_, _04505_, _17668_);
  or (_17682_, _17681_, _17680_);
  and (_17683_, _17682_, _02662_);
  nor (_17684_, _09087_, _05913_);
  nor (_17685_, _17684_, _17669_);
  nor (_17686_, _17685_, _02662_);
  or (_17688_, _17686_, _17683_);
  and (_17689_, _17688_, _03365_);
  nor (_17690_, _05913_, _04480_);
  nor (_17691_, _17690_, _17669_);
  nor (_17692_, _17691_, _03365_);
  nor (_17693_, _17692_, _17689_);
  nor (_17694_, _17693_, _03168_);
  or (_17695_, _17694_, _05949_);
  nor (_17696_, _17695_, _17679_);
  and (_17697_, _17691_, _05949_);
  nor (_17699_, _17697_, _17696_);
  nor (_17700_, _17699_, _05959_);
  and (_17701_, _04605_, _03904_);
  nor (_17702_, _17669_, _05963_);
  not (_17703_, _17702_);
  nor (_17704_, _17703_, _17701_);
  or (_17705_, _17704_, _02024_);
  nor (_17706_, _17705_, _17700_);
  nor (_17707_, _09180_, _05913_);
  nor (_17708_, _17707_, _17669_);
  nor (_17710_, _17708_, _03139_);
  or (_17711_, _17710_, _02575_);
  nor (_17712_, _17711_, _17706_);
  nor (_17713_, _17712_, _17675_);
  or (_17714_, _17713_, _02656_);
  and (_17715_, _09195_, _04605_);
  or (_17716_, _17715_, _17669_);
  or (_17717_, _17716_, _05305_);
  and (_17718_, _17717_, _03252_);
  and (_17719_, _17718_, _17714_);
  nor (_17721_, _17719_, _17672_);
  nor (_17722_, _17721_, _02669_);
  not (_17723_, _17669_);
  and (_17724_, _17723_, _04787_);
  not (_17725_, _17724_);
  nor (_17726_, _17674_, _05332_);
  and (_17727_, _17726_, _17725_);
  nor (_17728_, _17727_, _17722_);
  nor (_17729_, _17728_, _03243_);
  or (_17730_, _17724_, _03244_);
  nor (_17732_, _17730_, _17678_);
  or (_17733_, _17732_, _02654_);
  nor (_17734_, _17733_, _17729_);
  nor (_17735_, _09194_, _05913_);
  nor (_17736_, _17735_, _17669_);
  and (_17737_, _17736_, _02654_);
  nor (_17738_, _17737_, _17734_);
  and (_17739_, _17738_, _05883_);
  nor (_17740_, _09054_, _05913_);
  nor (_17741_, _17740_, _17669_);
  nor (_17743_, _17741_, _05883_);
  or (_17744_, _17743_, _17739_);
  and (_17745_, _17744_, _03124_);
  nor (_17746_, _17685_, _03124_);
  or (_17747_, _17746_, _17745_);
  and (_17748_, _17747_, _03513_);
  and (_17749_, _09248_, _04605_);
  nor (_17750_, _17749_, _17669_);
  nor (_17751_, _17750_, _03513_);
  or (_17752_, _17751_, _17748_);
  or (_17754_, _17752_, _27789_);
  or (_17755_, _27788_, \oc8051_golden_model_1.TMOD [5]);
  and (_17756_, _17755_, _27053_);
  and (_28954_, _17756_, _17754_);
  not (_17757_, \oc8051_golden_model_1.TMOD [6]);
  nor (_17758_, _04605_, _17757_);
  and (_17759_, _09268_, _04605_);
  nor (_17760_, _17759_, _17758_);
  nor (_17761_, _17760_, _03252_);
  and (_17762_, _04605_, _03960_);
  or (_17764_, _17762_, _17758_);
  and (_17765_, _17764_, _05959_);
  and (_17766_, _04605_, \oc8051_golden_model_1.ACC [6]);
  nor (_17767_, _17766_, _17758_);
  nor (_17768_, _17767_, _05903_);
  nor (_17769_, _04505_, _17757_);
  or (_17770_, _17769_, _17768_);
  and (_17771_, _17770_, _02662_);
  nor (_17772_, _09301_, _05913_);
  nor (_17773_, _17772_, _17758_);
  nor (_17775_, _17773_, _02662_);
  or (_17776_, _17775_, _17771_);
  and (_17777_, _17776_, _03365_);
  nor (_17778_, _05913_, _04373_);
  nor (_17779_, _17778_, _17758_);
  nor (_17780_, _17779_, _03365_);
  nor (_17781_, _17780_, _17777_);
  nor (_17782_, _17781_, _03168_);
  nor (_17783_, _17767_, _03179_);
  nor (_17784_, _17783_, _05949_);
  not (_17786_, _17784_);
  nor (_17787_, _17786_, _17782_);
  and (_17788_, _17779_, _05949_);
  or (_17789_, _17788_, _05959_);
  nor (_17790_, _17789_, _17787_);
  or (_17791_, _17790_, _17765_);
  and (_17792_, _17791_, _03139_);
  and (_17793_, _09388_, _04605_);
  nor (_17794_, _17793_, _17758_);
  nor (_17795_, _17794_, _03139_);
  or (_17797_, _17795_, _06549_);
  or (_17798_, _17797_, _17792_);
  and (_17799_, _09404_, _04605_);
  or (_17800_, _17758_, _05305_);
  or (_17801_, _17800_, _17799_);
  and (_17802_, _04605_, _09395_);
  nor (_17803_, _17802_, _17758_);
  and (_17804_, _17803_, _02575_);
  nor (_17805_, _17804_, _03251_);
  and (_17806_, _17805_, _17801_);
  and (_17808_, _17806_, _17798_);
  nor (_17809_, _17808_, _17761_);
  nor (_17810_, _17809_, _02669_);
  nor (_17811_, _17758_, _06119_);
  not (_17812_, _17811_);
  nor (_17813_, _17803_, _05332_);
  and (_17814_, _17813_, _17812_);
  nor (_17815_, _17814_, _17810_);
  nor (_17816_, _17815_, _03243_);
  or (_17817_, _17811_, _03244_);
  nor (_17819_, _17817_, _17767_);
  or (_17820_, _17819_, _02654_);
  nor (_17821_, _17820_, _17816_);
  nor (_17822_, _09403_, _05913_);
  nor (_17823_, _17822_, _17758_);
  and (_17824_, _17823_, _02654_);
  nor (_17825_, _17824_, _17821_);
  and (_17826_, _17825_, _05883_);
  nor (_17827_, _09267_, _05913_);
  nor (_17828_, _17827_, _17758_);
  nor (_17830_, _17828_, _05883_);
  or (_17831_, _17830_, _17826_);
  and (_17832_, _17831_, _03124_);
  nor (_17833_, _17773_, _03124_);
  or (_17834_, _17833_, _17832_);
  and (_17835_, _17834_, _03513_);
  and (_17836_, _09456_, _04605_);
  nor (_17837_, _17836_, _17758_);
  nor (_17838_, _17837_, _03513_);
  or (_17839_, _17838_, _17835_);
  or (_17841_, _17839_, _27789_);
  or (_17842_, _27788_, \oc8051_golden_model_1.TMOD [6]);
  and (_17843_, _17842_, _27053_);
  and (_28955_, _17843_, _17841_);
  and (_17844_, _05862_, _01647_);
  and (_17845_, _06742_, _03048_);
  and (_17846_, _05726_, _01930_);
  nor (_17847_, _17846_, _01647_);
  not (_17848_, _01957_);
  nor (_17849_, _02654_, _01944_);
  nor (_17851_, _17849_, _01647_);
  not (_17852_, _01965_);
  nor (_17853_, _05325_, _02669_);
  nor (_17854_, _17853_, _01647_);
  not (_17855_, _01974_);
  nor (_17856_, _05297_, _02656_);
  nor (_17857_, _17856_, _01647_);
  and (_17858_, _02575_, _01647_);
  nor (_17859_, _03048_, _01993_);
  and (_17860_, _03048_, \oc8051_golden_model_1.PC [0]);
  nor (_17862_, _17860_, _03049_);
  or (_17863_, _17862_, _04275_);
  or (_17864_, _04277_, _01647_);
  and (_17865_, _17864_, _02675_);
  and (_17866_, _17865_, _17863_);
  nor (_17867_, _03048_, _01990_);
  nor (_17868_, _04522_, _01647_);
  and (_17869_, _04521_, _01647_);
  nor (_17870_, _04521_, _01647_);
  nor (_17871_, _17870_, _17869_);
  and (_17873_, _17871_, _01988_);
  not (_17874_, _04522_);
  nor (_17875_, _03048_, _01988_);
  or (_17876_, _17875_, _17874_);
  nor (_17877_, _17876_, _17873_);
  or (_17878_, _17877_, _04527_);
  nor (_17879_, _17878_, _17868_);
  nor (_17880_, _03048_, _01998_);
  or (_17881_, _17880_, _03406_);
  nor (_17882_, _17881_, _17879_);
  and (_17883_, _04540_, \oc8051_golden_model_1.PC [0]);
  not (_17884_, _17883_);
  and (_17885_, _02503_, _01647_);
  nor (_17886_, _17885_, _02504_);
  and (_17887_, _17886_, _04537_);
  nor (_17888_, _17887_, _04539_);
  and (_17889_, _17888_, _17884_);
  nor (_17890_, _17889_, _17882_);
  nor (_17891_, _17890_, _04545_);
  and (_17892_, _04545_, \oc8051_golden_model_1.PC [0]);
  nor (_17895_, _17892_, _02661_);
  not (_17896_, _17895_);
  nor (_17897_, _17896_, _17891_);
  not (_17898_, _17897_);
  and (_17899_, _04985_, \oc8051_golden_model_1.PC [0]);
  not (_17900_, _17899_);
  not (_17901_, _17862_);
  and (_17902_, _17901_, _04987_);
  nor (_17903_, _17902_, _02662_);
  and (_17904_, _17903_, _17900_);
  nor (_17906_, _17904_, _04992_);
  and (_17907_, _17906_, _17898_);
  and (_17908_, _04992_, \oc8051_golden_model_1.PC [0]);
  nor (_17909_, _17908_, _07558_);
  not (_17910_, _17909_);
  nor (_17911_, _17910_, _17907_);
  nor (_17912_, _03048_, _01995_);
  nor (_17913_, _05009_, _05000_);
  not (_17914_, _17913_);
  nor (_17915_, _17914_, _17912_);
  not (_17917_, _17915_);
  nor (_17918_, _17917_, _17911_);
  not (_17919_, _01990_);
  nor (_17920_, _17913_, _01647_);
  nor (_17921_, _17920_, _17919_);
  not (_17922_, _17921_);
  nor (_17923_, _17922_, _17918_);
  or (_17924_, _17923_, _04498_);
  nor (_17925_, _17924_, _17867_);
  and (_17926_, _04494_, _01647_);
  nor (_17927_, _17901_, _04494_);
  or (_17928_, _17927_, _17926_);
  nor (_17929_, _17928_, _04499_);
  or (_17930_, _17929_, _02675_);
  nor (_17931_, _17930_, _17925_);
  or (_17932_, _17931_, _02664_);
  or (_17933_, _17932_, _17866_);
  and (_17934_, _05157_, _01647_);
  nor (_17935_, _17901_, _05157_);
  or (_17936_, _17935_, _03387_);
  or (_17939_, _17936_, _17934_);
  and (_17940_, _17939_, _05024_);
  and (_17941_, _17940_, _17933_);
  and (_17942_, _02630_, \oc8051_golden_model_1.PC [0]);
  nor (_17943_, _17862_, _02630_);
  or (_17944_, _17943_, _05024_);
  nor (_17945_, _17944_, _17942_);
  or (_17946_, _17945_, _17941_);
  and (_17947_, _17946_, _02599_);
  and (_17948_, _02598_, _01647_);
  or (_17950_, _17948_, _17947_);
  and (_17951_, _17950_, _02000_);
  nor (_17952_, _03048_, _02000_);
  nor (_17953_, _17952_, _05185_);
  not (_17954_, _17953_);
  nor (_17955_, _17954_, _17951_);
  not (_17956_, _01993_);
  and (_17957_, _05185_, \oc8051_golden_model_1.PC [0]);
  nor (_17958_, _17957_, _17956_);
  not (_17959_, _17958_);
  nor (_17961_, _17959_, _17955_);
  nor (_17962_, _05194_, _02047_);
  not (_17963_, _17962_);
  or (_17964_, _17963_, _17961_);
  nor (_17965_, _17964_, _17859_);
  nor (_17966_, _17962_, _01647_);
  nor (_17967_, _17966_, _02025_);
  not (_17968_, _17967_);
  nor (_17969_, _17968_, _17965_);
  nor (_17970_, _03048_, _07791_);
  or (_17972_, _05225_, _02024_);
  nor (_17973_, _17972_, _02670_);
  not (_17974_, _17973_);
  nor (_17975_, _17974_, _17970_);
  not (_17976_, _17975_);
  nor (_17977_, _17976_, _17969_);
  nor (_17978_, _17973_, _01647_);
  nor (_17979_, _17978_, _01960_);
  not (_17980_, _17979_);
  nor (_17981_, _17980_, _17977_);
  not (_17983_, _01960_);
  nor (_17984_, _03048_, _17983_);
  or (_17985_, _17984_, _05233_);
  nor (_17986_, _17985_, _17981_);
  nor (_17987_, _17886_, _05234_);
  nor (_17988_, _17987_, _17986_);
  and (_17989_, _17988_, _05245_);
  or (_17990_, _17989_, _17858_);
  and (_17991_, _17990_, _02574_);
  and (_17992_, _02573_, _02049_);
  or (_17994_, _17992_, _17991_);
  and (_17995_, _17994_, _13603_);
  nor (_17996_, _03048_, _13603_);
  or (_17997_, _17996_, _17995_);
  and (_17998_, _17997_, _05291_);
  not (_17999_, _17856_);
  nor (_18000_, _17886_, _01953_);
  and (_18001_, _01953_, _01647_);
  nor (_18002_, _18001_, _05291_);
  not (_18003_, _18002_);
  nor (_18005_, _18003_, _18000_);
  nor (_18006_, _18005_, _17999_);
  not (_18007_, _18006_);
  nor (_18008_, _18007_, _17998_);
  nor (_18009_, _18008_, _17857_);
  and (_18010_, _18009_, _17855_);
  nor (_18011_, _03048_, _17855_);
  or (_18012_, _18011_, _18010_);
  and (_18013_, _18012_, _05316_);
  not (_18014_, _17853_);
  nor (_18016_, _01953_, _01647_);
  and (_18017_, _17886_, _01953_);
  or (_18018_, _18017_, _18016_);
  and (_18019_, _18018_, _05315_);
  nor (_18020_, _18019_, _18014_);
  not (_18021_, _18020_);
  nor (_18022_, _18021_, _18013_);
  nor (_18023_, _18022_, _17854_);
  and (_18024_, _18023_, _17852_);
  nor (_18025_, _03048_, _17852_);
  or (_18027_, _18025_, _18024_);
  and (_18028_, _18027_, _05343_);
  not (_18029_, _17849_);
  nor (_18030_, _17886_, \oc8051_golden_model_1.PSW [7]);
  and (_18031_, \oc8051_golden_model_1.PSW [7], _01647_);
  nor (_18032_, _18031_, _05343_);
  not (_18033_, _18032_);
  nor (_18034_, _18033_, _18030_);
  nor (_18035_, _18034_, _18029_);
  not (_18036_, _18035_);
  nor (_18038_, _18036_, _18028_);
  nor (_18039_, _18038_, _17851_);
  and (_18040_, _18039_, _17848_);
  nor (_18041_, _03048_, _17848_);
  or (_18042_, _18041_, _18040_);
  and (_18043_, _18042_, _05368_);
  and (_18044_, _05348_, \oc8051_golden_model_1.PC [0]);
  and (_18045_, _17886_, \oc8051_golden_model_1.PSW [7]);
  or (_18046_, _18045_, _18044_);
  and (_18047_, _18046_, _05367_);
  and (_18049_, _05397_, _05389_);
  not (_18050_, _18049_);
  nor (_18051_, _18050_, _18047_);
  not (_18052_, _18051_);
  nor (_18053_, _18052_, _18043_);
  nor (_18054_, _18049_, _01647_);
  or (_18055_, _18054_, _03109_);
  nor (_18056_, _18055_, _18053_);
  and (_18057_, _04268_, _03109_);
  or (_18058_, _18057_, _18056_);
  and (_18060_, _18058_, _05408_);
  nor (_18061_, _03048_, _05408_);
  or (_18062_, _18061_, _18060_);
  and (_18063_, _18062_, _03267_);
  not (_18064_, _17846_);
  and (_18065_, _17901_, _05702_);
  nor (_18066_, _05702_, _01647_);
  or (_18067_, _18066_, _03267_);
  nor (_18068_, _18067_, _18065_);
  nor (_18069_, _18068_, _18064_);
  not (_18071_, _18069_);
  nor (_18072_, _18071_, _18063_);
  nor (_18073_, _18072_, _17847_);
  and (_18074_, _18073_, _03126_);
  and (_18075_, _04268_, _03108_);
  or (_18076_, _18075_, _18074_);
  and (_18077_, _18076_, _05748_);
  nor (_18078_, _03048_, _05748_);
  or (_18079_, _18078_, _02647_);
  or (_18080_, _18079_, _18077_);
  nor (_18082_, _05780_, _05764_);
  and (_18083_, _05702_, \oc8051_golden_model_1.PC [0]);
  nor (_18084_, _17862_, _05702_);
  nor (_18085_, _18084_, _18083_);
  or (_18086_, _18085_, _03125_);
  and (_18087_, _18086_, _18082_);
  and (_18088_, _18087_, _18080_);
  nor (_18089_, _18082_, \oc8051_golden_model_1.PC [0]);
  nor (_18090_, _18089_, _06742_);
  not (_18091_, _18090_);
  nor (_18093_, _18091_, _18088_);
  nor (_18094_, _18093_, _17845_);
  or (_18095_, _18094_, _02650_);
  and (_18096_, _05848_, _05824_);
  or (_18097_, _18085_, _03122_);
  and (_18098_, _18097_, _18096_);
  and (_18099_, _18098_, _18095_);
  nor (_18100_, _02649_, _01955_);
  not (_18101_, _18100_);
  nor (_18102_, _18096_, \oc8051_golden_model_1.PC [0]);
  nor (_18104_, _18102_, _18101_);
  not (_18105_, _18104_);
  nor (_18106_, _18105_, _18099_);
  and (_18107_, _18101_, _03048_);
  nor (_18108_, _18107_, _05862_);
  not (_18109_, _18108_);
  nor (_18110_, _18109_, _18106_);
  nor (_18111_, _18110_, _17844_);
  nand (_18112_, _18111_, _27788_);
  or (_18113_, _27788_, \oc8051_golden_model_1.PC [0]);
  and (_18115_, _18113_, _27053_);
  and (_28958_, _18115_, _18112_);
  nor (_18116_, _03051_, _03049_);
  nor (_18117_, _18116_, _03052_);
  nor (_18118_, _18117_, _05702_);
  and (_18119_, _05702_, _02006_);
  nor (_18120_, _18119_, _18118_);
  and (_18121_, _18120_, _02650_);
  and (_18122_, _03123_, _01620_);
  and (_18123_, _03016_, _01899_);
  and (_18125_, _01942_, _02639_);
  and (_18126_, _03251_, \oc8051_golden_model_1.PC [1]);
  and (_18127_, _02577_, \oc8051_golden_model_1.PC [1]);
  nor (_18128_, _05177_, _01620_);
  not (_18129_, _18117_);
  nor (_18130_, _18129_, _05157_);
  and (_18131_, _05157_, _02007_);
  nor (_18132_, _18131_, _18130_);
  nor (_18133_, _18132_, _03387_);
  not (_18134_, _04992_);
  and (_18136_, _04545_, _02007_);
  nor (_18137_, _02506_, _02504_);
  nor (_18138_, _18137_, _02507_);
  or (_18139_, _18138_, _04540_);
  or (_18140_, _04537_, _01620_);
  and (_18141_, _18140_, _03406_);
  nand (_18142_, _18141_, _18139_);
  and (_18143_, _03016_, _04527_);
  not (_18144_, _04502_);
  nor (_18145_, _02674_, _01917_);
  or (_18147_, _18145_, _01997_);
  nor (_18148_, _18147_, _02006_);
  and (_18149_, _03016_, _04504_);
  and (_18150_, _04512_, \oc8051_golden_model_1.PC [0]);
  not (_18151_, _04514_);
  and (_18152_, _04520_, _01647_);
  nor (_18153_, _18152_, _18151_);
  nor (_18154_, _18153_, _18150_);
  and (_18155_, _18154_, \oc8051_golden_model_1.PC [1]);
  nor (_18156_, _18154_, \oc8051_golden_model_1.PC [1]);
  nor (_18158_, _18156_, _18155_);
  and (_18159_, _18158_, _01988_);
  nor (_18160_, _03325_, _02007_);
  nor (_18161_, _18160_, _03328_);
  or (_18162_, _18161_, _18159_);
  nor (_18163_, _18162_, _18149_);
  not (_18164_, _18147_);
  nor (_18165_, _03328_, _02007_);
  nor (_18166_, _18165_, _18164_);
  not (_18167_, _18166_);
  nor (_18169_, _18167_, _18163_);
  nor (_18170_, _18169_, _18148_);
  and (_18171_, _18170_, _04503_);
  and (_18172_, _03154_, _01620_);
  or (_18173_, _18172_, _18171_);
  and (_18174_, _18173_, _18144_);
  and (_18175_, _04502_, _02006_);
  nor (_18176_, _18175_, _04527_);
  not (_18177_, _18176_);
  nor (_18178_, _18177_, _18174_);
  or (_18180_, _18178_, _03406_);
  nor (_18181_, _18180_, _18143_);
  nor (_18182_, _18181_, _04545_);
  and (_18183_, _18182_, _18142_);
  or (_18184_, _18183_, _18136_);
  nand (_18185_, _18184_, _02662_);
  and (_18186_, _18117_, _04987_);
  and (_18187_, _04985_, _02007_);
  nor (_18188_, _18187_, _18186_);
  nand (_18189_, _18188_, _02661_);
  nand (_18191_, _18189_, _18185_);
  nand (_18192_, _18191_, _18134_);
  and (_18193_, _04992_, _02007_);
  nor (_18194_, _18193_, _03150_);
  nand (_18195_, _18194_, _18192_);
  and (_18196_, _03150_, _01620_);
  nor (_18197_, _18196_, _07558_);
  nand (_18198_, _18197_, _18195_);
  and (_18199_, _03016_, _07558_);
  nor (_18200_, _18199_, _03162_);
  nand (_18202_, _18200_, _18198_);
  and (_18203_, _03162_, _01620_);
  nor (_18204_, _18203_, _05000_);
  nand (_18205_, _18204_, _18202_);
  and (_18206_, _05000_, _02007_);
  nor (_18207_, _18206_, _03168_);
  nand (_18208_, _18207_, _18205_);
  and (_18209_, _03168_, _01620_);
  nor (_18210_, _18209_, _05009_);
  and (_18211_, _18210_, _18208_);
  and (_18213_, _05009_, _02007_);
  or (_18214_, _18213_, _18211_);
  nand (_18215_, _18214_, _03177_);
  and (_18216_, _03176_, \oc8051_golden_model_1.PC [1]);
  nor (_18217_, _18216_, _17919_);
  and (_18218_, _18217_, _18215_);
  nor (_18219_, _03016_, _01990_);
  or (_18220_, _18219_, _18218_);
  nand (_18221_, _18220_, _03430_);
  and (_18222_, _03187_, _01620_);
  nor (_18224_, _18222_, _04498_);
  and (_18225_, _18224_, _18221_);
  and (_18226_, _04494_, _02007_);
  nor (_18227_, _18129_, _04494_);
  or (_18228_, _18227_, _18226_);
  nor (_18229_, _18228_, _04499_);
  or (_18230_, _18229_, _18225_);
  nand (_18231_, _18230_, _03107_);
  or (_18232_, _18129_, _04275_);
  or (_18233_, _04277_, _02006_);
  and (_18235_, _18233_, _02675_);
  nand (_18236_, _18235_, _18232_);
  and (_18237_, _18236_, _03387_);
  and (_18238_, _18237_, _18231_);
  or (_18239_, _18238_, _18133_);
  nand (_18240_, _18239_, _05024_);
  and (_18241_, _02630_, _02006_);
  nor (_18242_, _18117_, _02630_);
  or (_18243_, _18242_, _05024_);
  or (_18244_, _18243_, _18241_);
  and (_18246_, _18244_, _02599_);
  and (_18247_, _18246_, _18240_);
  and (_18248_, _02598_, _02007_);
  or (_18249_, _18248_, _18247_);
  nand (_18250_, _18249_, _05168_);
  and (_18251_, _03144_, \oc8051_golden_model_1.PC [1]);
  nor (_18252_, _18251_, _06664_);
  nand (_18253_, _18252_, _18250_);
  not (_18254_, _05177_);
  nor (_18255_, _03016_, _02000_);
  nor (_18257_, _18255_, _18254_);
  and (_18258_, _18257_, _18253_);
  or (_18259_, _18258_, _18128_);
  nand (_18260_, _18259_, _05186_);
  and (_18261_, _05185_, _02007_);
  nor (_18262_, _18261_, _03205_);
  nand (_18263_, _18262_, _18260_);
  and (_18264_, _03205_, _01620_);
  nor (_18265_, _18264_, _17956_);
  nand (_18266_, _18265_, _18263_);
  and (_18268_, _03016_, _17956_);
  nor (_18269_, _18268_, _03203_);
  nand (_18270_, _18269_, _18266_);
  and (_18271_, _03203_, _01620_);
  and (_18272_, _01983_, _01920_);
  nor (_18273_, _18272_, _18271_);
  nand (_18274_, _18273_, _18270_);
  and (_18275_, _18272_, _02007_);
  nor (_18276_, _18145_, _01984_);
  nor (_18277_, _18276_, _18275_);
  nand (_18279_, _18277_, _18274_);
  and (_18280_, _18276_, _02006_);
  nor (_18281_, _18280_, _05199_);
  nand (_18282_, _18281_, _18279_);
  and (_18283_, _05199_, \oc8051_golden_model_1.PC [1]);
  nor (_18284_, _18283_, _02047_);
  nand (_18285_, _18284_, _18282_);
  nor (_18286_, _02007_, _01985_);
  nor (_18287_, _18286_, _03140_);
  and (_18288_, _18287_, _18285_);
  and (_18290_, _03140_, \oc8051_golden_model_1.PC [1]);
  or (_18291_, _18290_, _18288_);
  nand (_18292_, _18291_, _07791_);
  and (_18293_, _03016_, _02025_);
  nor (_18294_, _18293_, _02670_);
  nand (_18295_, _18294_, _18292_);
  and (_18296_, _02670_, _02007_);
  nor (_18297_, _18296_, _05217_);
  nand (_18298_, _18297_, _18295_);
  and (_18299_, _05217_, \oc8051_golden_model_1.PC [1]);
  nor (_18301_, _18299_, _02024_);
  nand (_18302_, _18301_, _18298_);
  and (_18303_, _02024_, _02007_);
  nor (_18304_, _18303_, _05225_);
  and (_18305_, _18304_, _18302_);
  and (_18306_, _05225_, _02007_);
  or (_18307_, _18306_, _18305_);
  nand (_18308_, _18307_, _03462_);
  and (_18309_, _03135_, \oc8051_golden_model_1.PC [1]);
  nor (_18310_, _18309_, _01960_);
  and (_18312_, _18310_, _18308_);
  nor (_18313_, _03016_, _17983_);
  or (_18314_, _18313_, _18312_);
  nand (_18315_, _18314_, _05234_);
  and (_18316_, _18138_, _05233_);
  nor (_18317_, _18316_, _02577_);
  and (_18318_, _18317_, _18315_);
  or (_18319_, _18318_, _18127_);
  nand (_18320_, _18319_, _05245_);
  and (_18321_, _02575_, _02006_);
  nor (_18323_, _18321_, _05243_);
  nand (_18324_, _18323_, _18320_);
  and (_18325_, _05243_, _01620_);
  nor (_18326_, _18325_, _02573_);
  nand (_18327_, _18326_, _18324_);
  and (_18328_, _02573_, _02018_);
  nor (_18329_, _18328_, _03134_);
  nand (_18330_, _18329_, _18327_);
  and (_18331_, _03134_, _01620_);
  nor (_18332_, _18331_, _01967_);
  nand (_18334_, _18332_, _18330_);
  and (_18335_, _03016_, _01967_);
  nor (_18336_, _18335_, _02567_);
  nand (_18337_, _18336_, _18334_);
  nand (_18338_, _01953_, _01620_);
  nand (_18339_, _18138_, _02568_);
  and (_18340_, _18339_, _18338_);
  or (_18341_, _18340_, _05291_);
  and (_18342_, _18341_, _18337_);
  nor (_18343_, _05169_, _05296_);
  or (_18345_, _18343_, _18342_);
  and (_18346_, _03421_, _01916_);
  nor (_18347_, _05378_, _18346_);
  nor (_18348_, _18347_, _05296_);
  and (_18349_, _18343_, _02006_);
  nor (_18350_, _18349_, _18348_);
  nand (_18351_, _18350_, _18345_);
  and (_18352_, _18348_, _02007_);
  nor (_18353_, _18352_, _03469_);
  nand (_18354_, _18353_, _18351_);
  and (_18356_, _03469_, _02006_);
  nor (_18357_, _18356_, _05302_);
  nand (_18358_, _18357_, _18354_);
  and (_18359_, _05302_, \oc8051_golden_model_1.PC [1]);
  nor (_18360_, _18359_, _02656_);
  nand (_18361_, _18360_, _18358_);
  and (_18362_, _02656_, _02007_);
  nor (_18363_, _18362_, _03251_);
  and (_18364_, _18363_, _18361_);
  or (_18365_, _18364_, _18126_);
  nand (_18367_, _18365_, _17855_);
  and (_18368_, _03016_, _01974_);
  nor (_18369_, _18368_, _05315_);
  nand (_18370_, _18369_, _18367_);
  nor (_18371_, _01953_, \oc8051_golden_model_1.PC [1]);
  and (_18372_, _18138_, _01953_);
  or (_18373_, _18372_, _18371_);
  and (_18374_, _18373_, _05315_);
  and (_18375_, _01964_, _01920_);
  nor (_18376_, _18375_, _18374_);
  nand (_18378_, _18376_, _18370_);
  and (_18379_, _18375_, _02007_);
  nor (_18380_, _18145_, _03359_);
  nor (_18381_, _18380_, _18379_);
  nand (_18382_, _18381_, _18378_);
  and (_18383_, _18380_, _02006_);
  nor (_18384_, _18383_, _05329_);
  nand (_18385_, _18384_, _18382_);
  and (_18386_, _05329_, \oc8051_golden_model_1.PC [1]);
  nor (_18387_, _18386_, _02669_);
  nand (_18389_, _18387_, _18385_);
  and (_18390_, _02669_, _02007_);
  nor (_18391_, _18390_, _03243_);
  and (_18392_, _18391_, _18389_);
  and (_18393_, _03243_, \oc8051_golden_model_1.PC [1]);
  or (_18394_, _18393_, _18392_);
  nand (_18395_, _18394_, _17852_);
  and (_18396_, _03016_, _01965_);
  nor (_18397_, _18396_, _05342_);
  nand (_18398_, _18397_, _18395_);
  or (_18400_, _05348_, \oc8051_golden_model_1.PC [1]);
  nand (_18401_, _18138_, _05348_);
  and (_18402_, _18401_, _18400_);
  or (_18403_, _18402_, _05343_);
  and (_18404_, _18403_, _18398_);
  or (_18405_, _18404_, _18125_);
  and (_18406_, _18125_, _02006_);
  not (_18407_, _03326_);
  nand (_18408_, _07487_, _18407_);
  and (_18409_, _18408_, _01942_);
  nor (_18411_, _18409_, _18406_);
  nand (_18412_, _18411_, _18405_);
  and (_18413_, _18409_, _02007_);
  or (_18414_, _02640_, _02674_);
  and (_18415_, _01942_, _18414_);
  nor (_18416_, _18415_, _18413_);
  nand (_18417_, _18416_, _18412_);
  and (_18418_, _18415_, _02006_);
  nor (_18419_, _18418_, _05355_);
  nand (_18420_, _18419_, _18417_);
  and (_18422_, _05355_, \oc8051_golden_model_1.PC [1]);
  nor (_18423_, _18422_, _02654_);
  nand (_18424_, _18423_, _18420_);
  and (_18425_, _02654_, _02007_);
  nor (_18426_, _18425_, _03239_);
  and (_18427_, _18426_, _18424_);
  and (_18428_, _03239_, \oc8051_golden_model_1.PC [1]);
  or (_18429_, _18428_, _18427_);
  nand (_18430_, _18429_, _17848_);
  and (_18431_, _03016_, _01957_);
  nor (_18433_, _18431_, _05367_);
  nand (_18434_, _18433_, _18430_);
  nor (_18435_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_18436_, _18138_, \oc8051_golden_model_1.PSW [7]);
  or (_18437_, _18436_, _18435_);
  and (_18438_, _18437_, _05367_);
  nor (_18439_, _18438_, _05387_);
  and (_18440_, _18439_, _18434_);
  and (_18441_, _05387_, _02007_);
  or (_18442_, _18441_, _18440_);
  nand (_18444_, _18442_, _05385_);
  and (_18445_, _05384_, _02007_);
  nor (_18446_, _18445_, _05386_);
  nand (_18447_, _18446_, _18444_);
  and (_18448_, _05386_, _02006_);
  nor (_18449_, _18448_, _05393_);
  nand (_18450_, _18449_, _18447_);
  and (_18451_, _05393_, \oc8051_golden_model_1.PC [1]);
  nor (_18452_, _18451_, _05396_);
  and (_18453_, _18452_, _18450_);
  and (_18455_, _05396_, _02006_);
  or (_18456_, _18455_, _18453_);
  nand (_18457_, _18456_, _06612_);
  and (_18458_, _04218_, _03109_);
  nor (_18459_, _18458_, _01936_);
  nand (_18460_, _18459_, _18457_);
  and (_18461_, _03016_, _01936_);
  nor (_18462_, _18461_, _02653_);
  nand (_18463_, _18462_, _18460_);
  and (_18464_, _18129_, _05702_);
  not (_18466_, _18464_);
  nor (_18467_, _05702_, _02007_);
  nor (_18468_, _18467_, _03267_);
  and (_18469_, _18468_, _18466_);
  nor (_18470_, _18469_, _01923_);
  and (_18471_, _18470_, _18463_);
  nor (_18472_, _02007_, _01929_);
  nor (_18473_, _18472_, _01930_);
  or (_18474_, _18473_, _18471_);
  and (_18475_, _02006_, _01929_);
  nor (_18477_, _18475_, _05720_);
  nand (_18478_, _18477_, _18474_);
  and (_18479_, _05720_, \oc8051_golden_model_1.PC [1]);
  nor (_18480_, _18479_, _05724_);
  nand (_18481_, _18480_, _18478_);
  and (_18482_, _05724_, _02006_);
  nor (_18483_, _18482_, _03108_);
  and (_18484_, _18483_, _18481_);
  and (_18485_, _04221_, _03108_);
  or (_18486_, _18485_, _18484_);
  and (_18488_, _18486_, _05748_);
  or (_18489_, _18488_, _18123_);
  nand (_18490_, _18489_, _03125_);
  and (_18491_, _01970_, _01927_);
  nor (_18492_, _18120_, _03125_);
  nor (_18493_, _18492_, _18491_);
  nand (_18494_, _18493_, _18490_);
  and (_18495_, _18491_, _02006_);
  nor (_18496_, _18495_, _07491_);
  nand (_18497_, _18496_, _18494_);
  nor (_18499_, _07490_, _02006_);
  nor (_18500_, _18499_, _03123_);
  and (_18501_, _18500_, _18497_);
  or (_18502_, _18501_, _18122_);
  nand (_18503_, _18502_, _05788_);
  and (_18504_, _05780_, _02006_);
  nor (_18505_, _18504_, _06742_);
  nand (_18506_, _18505_, _18503_);
  and (_18507_, _06742_, _03016_);
  nor (_18508_, _18507_, _02650_);
  and (_18510_, _18508_, _18506_);
  or (_18511_, _18510_, _18121_);
  nand (_18512_, _18511_, _08578_);
  and (_18513_, _05820_, _02006_);
  nor (_18514_, _05812_, _05816_);
  not (_18515_, _18514_);
  nor (_18516_, _18515_, _18513_);
  nand (_18517_, _18516_, _18512_);
  nor (_18518_, _18514_, _02006_);
  nor (_18519_, _18518_, _03121_);
  nand (_18521_, _18519_, _18517_);
  and (_18522_, _03121_, _01620_);
  nor (_18523_, _18522_, _05840_);
  and (_18524_, _18523_, _18521_);
  and (_18525_, _05840_, _02007_);
  or (_18526_, _18525_, _18524_);
  nand (_18527_, _18526_, _18100_);
  and (_18528_, _18101_, _03016_);
  nor (_18529_, _18528_, _05862_);
  nand (_18530_, _18529_, _18527_);
  and (_18532_, _05862_, _02006_);
  not (_18533_, _18532_);
  nand (_18534_, _18533_, _18530_);
  or (_18535_, _18534_, _27789_);
  or (_18536_, _27788_, \oc8051_golden_model_1.PC [1]);
  and (_18537_, _18536_, _27053_);
  and (_28959_, _18537_, _18535_);
  and (_18538_, _05862_, _02080_);
  not (_18539_, _18538_);
  and (_18540_, _03121_, _02086_);
  and (_18542_, _03123_, _02086_);
  and (_18543_, _04168_, _03108_);
  nor (_18544_, _02080_, _01930_);
  and (_18545_, _04168_, _03109_);
  nor (_18546_, _05389_, _02080_);
  and (_18547_, _01966_, _02637_);
  and (_18548_, _01959_, _01928_);
  nand (_18549_, _05194_, _02682_);
  nand (_18550_, _02598_, _02682_);
  and (_18551_, _04494_, _02983_);
  and (_18553_, _03056_, _03053_);
  nor (_18554_, _18553_, _03057_);
  not (_18555_, _18554_);
  nor (_18556_, _18555_, _04494_);
  or (_18557_, _18556_, _18551_);
  or (_18558_, _18557_, _04499_);
  or (_18559_, _18554_, _04985_);
  or (_18560_, _04987_, _02983_);
  and (_18561_, _18560_, _18559_);
  or (_18562_, _18561_, _02662_);
  and (_18564_, _04540_, _02086_);
  and (_18565_, _02511_, _02508_);
  nor (_18566_, _18565_, _02512_);
  and (_18567_, _18566_, _04537_);
  or (_18568_, _18567_, _18564_);
  or (_18569_, _18568_, _04539_);
  nand (_18570_, _02981_, _04504_);
  and (_18571_, _04510_, _02682_);
  nor (_18572_, _18571_, _03154_);
  or (_18573_, _04521_, _02080_);
  nand (_18575_, _04505_, _02408_);
  or (_18576_, _04512_, \oc8051_golden_model_1.PC [2]);
  or (_18577_, _18576_, _04505_);
  and (_18578_, _18577_, _18575_);
  or (_18579_, _18578_, _04520_);
  and (_18580_, _18579_, _18573_);
  nor (_18581_, _04510_, _04504_);
  not (_18582_, _18581_);
  or (_18583_, _18582_, _18580_);
  and (_18584_, _18583_, _18572_);
  and (_18585_, _18584_, _18570_);
  and (_18586_, _03154_, _02086_);
  or (_18587_, _18586_, _04502_);
  or (_18588_, _18587_, _18585_);
  nand (_18589_, _04502_, _02682_);
  and (_18590_, _18589_, _01998_);
  and (_18591_, _18590_, _18588_);
  nor (_18592_, _02981_, _01998_);
  or (_18593_, _18592_, _03406_);
  or (_18594_, _18593_, _18591_);
  and (_18596_, _18594_, _07798_);
  and (_18597_, _18596_, _18569_);
  and (_18598_, _04545_, _02080_);
  or (_18599_, _18598_, _02661_);
  or (_18600_, _18599_, _18597_);
  and (_18601_, _18600_, _18562_);
  or (_18602_, _18601_, _04992_);
  nand (_18603_, _04992_, _02682_);
  and (_18604_, _18603_, _03390_);
  and (_18605_, _18604_, _18602_);
  and (_18607_, _03150_, _02086_);
  or (_18608_, _18607_, _07558_);
  or (_18609_, _18608_, _18605_);
  nand (_18610_, _02981_, _07558_);
  and (_18611_, _18610_, _03365_);
  and (_18612_, _18611_, _18609_);
  and (_18613_, _03162_, _02086_);
  or (_18614_, _18613_, _05000_);
  or (_18615_, _18614_, _18612_);
  and (_18616_, _05000_, _02682_);
  nor (_18618_, _18616_, _03168_);
  and (_18619_, _18618_, _18615_);
  and (_18620_, _03168_, _02086_);
  or (_18621_, _18620_, _05009_);
  or (_18622_, _18621_, _18619_);
  nand (_18623_, _05009_, _02682_);
  and (_18624_, _18623_, _03177_);
  and (_18625_, _18624_, _18622_);
  and (_18626_, _03176_, _02086_);
  or (_18627_, _18626_, _17919_);
  or (_18629_, _18627_, _18625_);
  nand (_18630_, _02981_, _17919_);
  and (_18631_, _18630_, _03430_);
  and (_18632_, _18631_, _18629_);
  and (_18633_, _03187_, _02086_);
  or (_18634_, _18633_, _04498_);
  or (_18635_, _18634_, _18632_);
  and (_18636_, _18635_, _18558_);
  or (_18637_, _18636_, _02675_);
  and (_18638_, _04275_, _02983_);
  and (_18640_, _18554_, _04277_);
  or (_18641_, _18640_, _03107_);
  or (_18642_, _18641_, _18638_);
  and (_18643_, _18642_, _18637_);
  or (_18644_, _18643_, _02664_);
  nor (_18645_, _18555_, _05157_);
  and (_18646_, _05157_, _02983_);
  or (_18647_, _18646_, _03387_);
  or (_18648_, _18647_, _18645_);
  and (_18649_, _18648_, _05024_);
  and (_18651_, _18649_, _18644_);
  or (_18652_, _18554_, _02630_);
  nand (_18653_, _02984_, _02630_);
  and (_18654_, _18653_, _02673_);
  and (_18655_, _18654_, _18652_);
  or (_18656_, _18655_, _02598_);
  or (_18657_, _18656_, _18651_);
  and (_18658_, _18657_, _18550_);
  or (_18659_, _18658_, _03144_);
  nand (_18660_, _03144_, _02408_);
  and (_18662_, _18660_, _02000_);
  and (_18663_, _18662_, _18659_);
  nor (_18664_, _02981_, _02000_);
  or (_18665_, _18664_, _18254_);
  or (_18666_, _18665_, _18663_);
  or (_18667_, _05177_, _02086_);
  and (_18668_, _18667_, _18666_);
  or (_18669_, _18668_, _05185_);
  and (_18670_, _05185_, _02682_);
  nor (_18671_, _18670_, _03205_);
  and (_18673_, _18671_, _18669_);
  and (_18674_, _03205_, _02086_);
  or (_18675_, _18674_, _17956_);
  or (_18676_, _18675_, _18673_);
  not (_18677_, _03203_);
  nand (_18678_, _02981_, _17956_);
  and (_18679_, _18678_, _18677_);
  and (_18680_, _18679_, _18676_);
  and (_18681_, _03203_, _02086_);
  or (_18682_, _18681_, _05194_);
  or (_18684_, _18682_, _18680_);
  and (_18685_, _18684_, _18549_);
  or (_18686_, _18685_, _05199_);
  nand (_18687_, _05199_, _02408_);
  and (_18688_, _18687_, _01985_);
  and (_18689_, _18688_, _18686_);
  nor (_18690_, _02682_, _01985_);
  or (_18691_, _18690_, _03140_);
  or (_18692_, _18691_, _18689_);
  nand (_18693_, _03140_, _02408_);
  and (_18695_, _18693_, _18692_);
  or (_18696_, _18695_, _02025_);
  nand (_18697_, _02981_, _02025_);
  and (_18698_, _18697_, _05212_);
  and (_18699_, _18698_, _18696_);
  nand (_18700_, _01959_, _01927_);
  nand (_18701_, _02983_, _02670_);
  nand (_18702_, _18701_, _18700_);
  or (_18703_, _18702_, _18699_);
  or (_18704_, _18700_, _02086_);
  and (_18706_, _18704_, _18703_);
  or (_18707_, _18706_, _18548_);
  nand (_18708_, _18548_, _02408_);
  and (_18709_, _18708_, _03139_);
  and (_18710_, _18709_, _18707_);
  and (_18711_, _02983_, _02024_);
  or (_18712_, _18711_, _05225_);
  or (_18713_, _18712_, _18710_);
  nand (_18714_, _05225_, _02682_);
  and (_18715_, _18714_, _03462_);
  and (_18717_, _18715_, _18713_);
  and (_18718_, _03135_, _02086_);
  or (_18719_, _18718_, _01960_);
  or (_18720_, _18719_, _18717_);
  nand (_18721_, _02981_, _01960_);
  and (_18722_, _18721_, _18720_);
  or (_18723_, _18722_, _05233_);
  and (_18724_, _01966_, _02639_);
  nor (_18725_, _18566_, _05234_);
  nor (_18726_, _18725_, _18724_);
  and (_18727_, _18726_, _18723_);
  and (_18728_, _18724_, _02086_);
  nor (_18729_, _18728_, _18727_);
  nor (_18730_, _18729_, _18547_);
  and (_18731_, _18547_, _02086_);
  and (_18732_, _07487_, _03358_);
  nor (_18733_, _18732_, _02576_);
  or (_18734_, _18733_, _18731_);
  or (_18735_, _18734_, _18730_);
  and (_18736_, _18733_, _02408_);
  and (_18738_, _07710_, _02565_);
  or (_18739_, _18738_, _07322_);
  nor (_18740_, _18739_, _18736_);
  and (_18741_, _18740_, _18735_);
  and (_18742_, _18739_, _02086_);
  or (_18743_, _18742_, _02575_);
  or (_18744_, _18743_, _18741_);
  nand (_18745_, _02984_, _02575_);
  and (_18746_, _18745_, _05244_);
  and (_18747_, _18746_, _18744_);
  and (_18749_, _05243_, _02086_);
  or (_18750_, _18749_, _02573_);
  or (_18751_, _18750_, _18747_);
  not (_18752_, _03134_);
  or (_18753_, _02574_, _02075_);
  and (_18754_, _18753_, _18752_);
  and (_18755_, _18754_, _18751_);
  and (_18756_, _03134_, _02086_);
  or (_18757_, _18756_, _01967_);
  or (_18758_, _18757_, _18755_);
  nand (_18760_, _02981_, _01967_);
  and (_18761_, _18760_, _05291_);
  and (_18762_, _18761_, _18758_);
  or (_18763_, _18566_, _01953_);
  nand (_18764_, _02408_, _01953_);
  and (_18765_, _18764_, _02567_);
  and (_18766_, _18765_, _18763_);
  or (_18767_, _18766_, _05297_);
  or (_18768_, _18767_, _18762_);
  nand (_18769_, _05297_, _02682_);
  and (_18771_, _18769_, _05306_);
  nand (_18772_, _18771_, _18768_);
  nand (_18773_, _05302_, _02086_);
  and (_18774_, _18773_, _18772_);
  nor (_18775_, _18774_, _02656_);
  and (_18776_, _02983_, _02656_);
  or (_18777_, _18776_, _03251_);
  nor (_18778_, _18777_, _18775_);
  and (_18779_, _03251_, _02408_);
  nor (_18780_, _18779_, _18778_);
  nand (_18782_, _18780_, _17855_);
  or (_18783_, _02981_, _17855_);
  and (_18784_, _18783_, _18782_);
  or (_18785_, _18784_, _05315_);
  nor (_18786_, _02408_, _01953_);
  and (_18787_, _18566_, _01953_);
  or (_18788_, _18787_, _18786_);
  and (_18789_, _18788_, _05315_);
  nor (_18790_, _18789_, _05325_);
  nand (_18791_, _18790_, _18785_);
  and (_18793_, _05325_, _02682_);
  nor (_18794_, _18793_, _05329_);
  nand (_18795_, _18794_, _18791_);
  and (_18796_, _05329_, _02086_);
  nor (_18797_, _18796_, _02669_);
  nand (_18798_, _18797_, _18795_);
  and (_18799_, _02984_, _02669_);
  nor (_18800_, _18799_, _03243_);
  nand (_18801_, _18800_, _18798_);
  and (_18802_, _03243_, _02086_);
  nor (_18804_, _18802_, _01965_);
  nand (_18805_, _18804_, _18801_);
  and (_18806_, _02981_, _01965_);
  nor (_18807_, _18806_, _05342_);
  nand (_18808_, _18807_, _18805_);
  nor (_18809_, _18566_, \oc8051_golden_model_1.PSW [7]);
  nor (_18810_, _02086_, _05348_);
  nor (_18811_, _18810_, _05343_);
  not (_18812_, _18811_);
  nor (_18813_, _18812_, _18809_);
  nor (_18815_, _18813_, _01944_);
  nand (_18816_, _18815_, _18808_);
  and (_18817_, _02682_, _01944_);
  nor (_18818_, _18817_, _05355_);
  and (_18819_, _18818_, _18816_);
  and (_18820_, _05355_, _02086_);
  or (_18821_, _18820_, _18819_);
  nand (_18822_, _18821_, _05357_);
  and (_18823_, _02983_, _02654_);
  nor (_18824_, _18823_, _03239_);
  and (_18825_, _18824_, _18822_);
  and (_18826_, _03239_, _02408_);
  or (_18827_, _18826_, _18825_);
  nand (_18828_, _18827_, _17848_);
  and (_18829_, _02981_, _01957_);
  nor (_18830_, _18829_, _05367_);
  nand (_18831_, _18830_, _18828_);
  nor (_18832_, _18566_, _05348_);
  nor (_18833_, _02086_, \oc8051_golden_model_1.PSW [7]);
  nor (_18834_, _18833_, _05368_);
  not (_18837_, _18834_);
  nor (_18838_, _18837_, _18832_);
  nor (_18839_, _18838_, _05391_);
  and (_18840_, _18839_, _18831_);
  or (_18841_, _18840_, _18546_);
  nand (_18842_, _18841_, _05398_);
  and (_18843_, _05393_, _02408_);
  nor (_18844_, _18843_, _05396_);
  nand (_18845_, _18844_, _18842_);
  and (_18846_, _05396_, _02080_);
  nor (_18848_, _18846_, _03109_);
  and (_18849_, _18848_, _18845_);
  or (_18850_, _18849_, _18545_);
  nand (_18851_, _18850_, _05408_);
  and (_18852_, _02981_, _01936_);
  nor (_18853_, _18852_, _02653_);
  nand (_18854_, _18853_, _18851_);
  nor (_18855_, _05702_, _02983_);
  and (_18856_, _18555_, _05702_);
  or (_18857_, _18856_, _03267_);
  nor (_18859_, _18857_, _18855_);
  nor (_18860_, _18859_, _05412_);
  and (_18861_, _18860_, _18854_);
  or (_18862_, _18861_, _18544_);
  nand (_18863_, _18862_, _05728_);
  and (_18864_, _05720_, _02408_);
  nor (_18865_, _18864_, _05724_);
  nand (_18866_, _18865_, _18863_);
  and (_18867_, _05724_, _02080_);
  nor (_18868_, _18867_, _03108_);
  and (_18870_, _18868_, _18866_);
  or (_18871_, _18870_, _18543_);
  nand (_18872_, _18871_, _05748_);
  and (_18873_, _02981_, _01899_);
  nor (_18874_, _18873_, _02647_);
  nand (_18875_, _18874_, _18872_);
  nor (_18876_, _18554_, _05702_);
  and (_18877_, _05702_, _02984_);
  nor (_18878_, _18877_, _18876_);
  and (_18879_, _18878_, _02647_);
  nor (_18881_, _18879_, _05764_);
  nand (_18882_, _18881_, _18875_);
  and (_18883_, _05764_, _02682_);
  nor (_18884_, _18883_, _03123_);
  and (_18885_, _18884_, _18882_);
  or (_18886_, _18885_, _18542_);
  nand (_18887_, _18886_, _05788_);
  and (_18888_, _05780_, _02080_);
  nor (_18889_, _18888_, _06742_);
  nand (_18890_, _18889_, _18887_);
  and (_18892_, _06742_, _02981_);
  nor (_18893_, _18892_, _02650_);
  nand (_18894_, _18893_, _18890_);
  and (_18895_, _18878_, _02650_);
  nor (_18896_, _18895_, _05826_);
  nand (_18897_, _18896_, _18894_);
  nor (_18898_, _05824_, _02080_);
  nor (_18899_, _18898_, _03121_);
  and (_18900_, _18899_, _18897_);
  or (_18901_, _18900_, _18540_);
  nand (_18903_, _18901_, _05848_);
  and (_18904_, _05840_, _02080_);
  nor (_18905_, _18904_, _18101_);
  nand (_18906_, _18905_, _18903_);
  and (_18907_, _18101_, _02981_);
  nor (_18908_, _18907_, _05862_);
  nand (_18909_, _18908_, _18906_);
  and (_18910_, _18909_, _18539_);
  nand (_18911_, _18910_, _27788_);
  or (_18912_, _27788_, \oc8051_golden_model_1.PC [2]);
  and (_18914_, _18912_, _27053_);
  and (_28960_, _18914_, _18911_);
  and (_18915_, _05862_, _02686_);
  not (_18916_, _18915_);
  and (_18917_, _03121_, _02107_);
  and (_18918_, _03123_, _02107_);
  nor (_18919_, _01930_, _02686_);
  and (_18920_, _04118_, _03109_);
  nor (_18921_, _05389_, _02686_);
  and (_18922_, _01944_, _02122_);
  and (_18923_, _05325_, _02122_);
  and (_18924_, _05297_, _02122_);
  and (_18925_, _02577_, _02108_);
  and (_18926_, _03140_, _02108_);
  and (_18927_, _05194_, _02122_);
  nor (_18928_, _05177_, _02107_);
  and (_18929_, _02598_, _02122_);
  and (_18930_, _04494_, _02947_);
  or (_18931_, _02950_, _02949_);
  and (_18932_, _18931_, _03058_);
  nor (_18934_, _18931_, _03058_);
  nor (_18935_, _18934_, _18932_);
  not (_18936_, _18935_);
  nor (_18937_, _18936_, _04494_);
  or (_18938_, _18937_, _18930_);
  nor (_18939_, _18938_, _04499_);
  or (_18940_, _18935_, _04985_);
  or (_18941_, _04987_, _02947_);
  and (_18942_, _18941_, _18940_);
  or (_18943_, _18942_, _02662_);
  and (_18945_, _04540_, _02107_);
  or (_18946_, _02407_, _02406_);
  and (_18947_, _18946_, _02513_);
  nor (_18948_, _18946_, _02513_);
  nor (_18949_, _18948_, _18947_);
  and (_18950_, _18949_, _04537_);
  nor (_18951_, _18950_, _18945_);
  nand (_18952_, _18951_, _03406_);
  nor (_18953_, _04512_, \oc8051_golden_model_1.PC [3]);
  nor (_18954_, _18953_, _04505_);
  not (_18956_, _18954_);
  and (_18957_, _04505_, _02107_);
  nor (_18958_, _18957_, _04520_);
  and (_18959_, _18958_, _18956_);
  not (_18960_, _18959_);
  nor (_18961_, _04521_, _02686_);
  nor (_18962_, _18961_, _04504_);
  and (_18963_, _18962_, _18960_);
  nor (_18964_, _02945_, _01988_);
  or (_18965_, _18964_, _04510_);
  nor (_18967_, _18965_, _18963_);
  and (_18968_, _04510_, _02122_);
  nor (_18969_, _18968_, _03154_);
  not (_18970_, _18969_);
  nor (_18971_, _18970_, _18967_);
  and (_18972_, _03154_, _02107_);
  or (_18973_, _18972_, _18971_);
  and (_18974_, _18973_, _18144_);
  and (_18975_, _04502_, _02686_);
  or (_18976_, _18975_, _18974_);
  and (_18978_, _18976_, _01998_);
  nor (_18979_, _02945_, _01998_);
  nor (_18980_, _18979_, _03406_);
  not (_18981_, _18980_);
  nor (_18982_, _18981_, _18978_);
  nor (_18983_, _18982_, _04545_);
  and (_18984_, _18983_, _18952_);
  and (_18985_, _04545_, _02686_);
  or (_18986_, _18985_, _02661_);
  or (_18987_, _18986_, _18984_);
  nand (_18989_, _18987_, _18943_);
  nand (_18990_, _18989_, _18134_);
  and (_18991_, _04992_, _02122_);
  nor (_18992_, _18991_, _03150_);
  nand (_18993_, _18992_, _18990_);
  and (_18994_, _03150_, _02107_);
  nor (_18995_, _18994_, _07558_);
  nand (_18996_, _18995_, _18993_);
  and (_18997_, _02945_, _07558_);
  nor (_18998_, _18997_, _03162_);
  nand (_19000_, _18998_, _18996_);
  and (_19001_, _03162_, _02107_);
  nor (_19002_, _19001_, _05000_);
  nand (_19003_, _19002_, _19000_);
  and (_19004_, _05000_, _02122_);
  nor (_19005_, _19004_, _03168_);
  nand (_19006_, _19005_, _19003_);
  and (_19007_, _03168_, _02107_);
  nor (_19008_, _19007_, _05009_);
  nand (_19009_, _19008_, _19006_);
  and (_19011_, _05009_, _02122_);
  nor (_19012_, _19011_, _03176_);
  nand (_19013_, _19012_, _19009_);
  and (_19014_, _03176_, _02107_);
  nor (_19015_, _19014_, _17919_);
  nand (_19016_, _19015_, _19013_);
  and (_19017_, _02945_, _17919_);
  nor (_19018_, _19017_, _03187_);
  nand (_19019_, _19018_, _19016_);
  and (_19020_, _03187_, _02107_);
  nor (_19022_, _19020_, _04498_);
  and (_19023_, _19022_, _19019_);
  nor (_19024_, _19023_, _18939_);
  or (_19025_, _19024_, _02675_);
  and (_19026_, _18935_, _04277_);
  and (_19027_, _04275_, _02947_);
  or (_19028_, _19027_, _03107_);
  or (_19029_, _19028_, _19026_);
  nand (_19030_, _19029_, _19025_);
  or (_19031_, _19030_, _02664_);
  nor (_19033_, _18936_, _05157_);
  and (_19034_, _05157_, _02947_);
  nor (_19035_, _19034_, _19033_);
  or (_19036_, _19035_, _03387_);
  and (_19037_, _19036_, _19031_);
  or (_19038_, _19037_, _02673_);
  nor (_19039_, _18935_, _02630_);
  and (_19040_, _02948_, _02630_);
  or (_19041_, _19040_, _05024_);
  or (_19042_, _19041_, _19039_);
  and (_19044_, _19042_, _02599_);
  and (_19045_, _19044_, _19038_);
  or (_19046_, _19045_, _18929_);
  nand (_19047_, _19046_, _05168_);
  and (_19048_, _03144_, _02108_);
  nor (_19049_, _19048_, _06664_);
  nand (_19050_, _19049_, _19047_);
  nor (_19051_, _02945_, _02000_);
  nor (_19052_, _19051_, _18254_);
  and (_19053_, _19052_, _19050_);
  or (_19055_, _19053_, _18928_);
  nand (_19056_, _19055_, _05186_);
  and (_19057_, _05185_, _02122_);
  nor (_19058_, _19057_, _03205_);
  nand (_19059_, _19058_, _19056_);
  and (_19060_, _03205_, _02107_);
  nor (_19061_, _19060_, _17956_);
  nand (_19062_, _19061_, _19059_);
  and (_19063_, _02945_, _17956_);
  nor (_19064_, _19063_, _03203_);
  nand (_19066_, _19064_, _19062_);
  and (_19067_, _03203_, _02107_);
  nor (_19068_, _19067_, _05194_);
  and (_19069_, _19068_, _19066_);
  or (_19070_, _19069_, _18927_);
  nand (_19071_, _19070_, _05203_);
  and (_19072_, _05199_, _02108_);
  nor (_19073_, _19072_, _02047_);
  nand (_19074_, _19073_, _19071_);
  nor (_19075_, _01985_, _02122_);
  nor (_19077_, _19075_, _03140_);
  and (_19078_, _19077_, _19074_);
  or (_19079_, _19078_, _18926_);
  nand (_19080_, _19079_, _07791_);
  and (_19081_, _02945_, _02025_);
  nor (_19082_, _19081_, _02670_);
  nand (_19083_, _19082_, _19080_);
  and (_19084_, _02947_, _02670_);
  nor (_19085_, _19084_, _05217_);
  nand (_19086_, _19085_, _19083_);
  and (_19088_, _05217_, _02108_);
  nor (_19089_, _19088_, _02024_);
  nand (_19090_, _19089_, _19086_);
  and (_19091_, _02947_, _02024_);
  nor (_19092_, _19091_, _05225_);
  nand (_19093_, _19092_, _19090_);
  and (_19094_, _05225_, _02122_);
  nor (_19095_, _19094_, _03135_);
  nand (_19096_, _19095_, _19093_);
  and (_19097_, _03135_, _02107_);
  nor (_19099_, _19097_, _01960_);
  nand (_19100_, _19099_, _19096_);
  and (_19101_, _02945_, _01960_);
  nor (_19102_, _19101_, _05233_);
  nand (_19103_, _19102_, _19100_);
  and (_19104_, _18949_, _05233_);
  nor (_19105_, _19104_, _02577_);
  and (_19106_, _19105_, _19103_);
  or (_19107_, _19106_, _18925_);
  nand (_19108_, _19107_, _05245_);
  and (_19109_, _02948_, _02575_);
  nor (_19110_, _19109_, _05243_);
  nand (_19111_, _19110_, _19108_);
  and (_19112_, _05243_, _02107_);
  nor (_19113_, _19112_, _02573_);
  nand (_19114_, _19113_, _19111_);
  nor (_19115_, _02574_, _02118_);
  nor (_19116_, _19115_, _03134_);
  and (_19117_, _19116_, _19114_);
  and (_19118_, _03134_, _02107_);
  or (_19120_, _19118_, _01967_);
  or (_19121_, _19120_, _19117_);
  and (_19122_, _02945_, _01967_);
  nor (_19123_, _19122_, _02567_);
  nand (_19124_, _19123_, _19121_);
  and (_19125_, _02107_, _01953_);
  and (_19126_, _18949_, _02568_);
  or (_19127_, _19126_, _19125_);
  and (_19128_, _19127_, _02567_);
  nor (_19129_, _19128_, _05297_);
  and (_19131_, _19129_, _19124_);
  or (_19132_, _19131_, _18924_);
  nand (_19133_, _19132_, _05306_);
  and (_19134_, _05302_, _02108_);
  nor (_19135_, _19134_, _02656_);
  and (_19136_, _19135_, _19133_);
  and (_19137_, _02947_, _02656_);
  or (_19138_, _19137_, _03251_);
  nor (_19139_, _19138_, _19136_);
  and (_19140_, _03251_, _02108_);
  or (_19142_, _19140_, _19139_);
  nand (_19143_, _19142_, _17855_);
  and (_19144_, _02945_, _01974_);
  nor (_19145_, _19144_, _05315_);
  nand (_19146_, _19145_, _19143_);
  and (_19147_, _02107_, _02568_);
  and (_19148_, _18949_, _01953_);
  or (_19149_, _19148_, _19147_);
  and (_19150_, _19149_, _05315_);
  nor (_19151_, _19150_, _05325_);
  and (_19153_, _19151_, _19146_);
  or (_19154_, _19153_, _18923_);
  nand (_19155_, _19154_, _05333_);
  and (_19156_, _05329_, _02108_);
  nor (_19157_, _19156_, _02669_);
  and (_19158_, _19157_, _19155_);
  and (_19159_, _02947_, _02669_);
  or (_19160_, _19159_, _03243_);
  nor (_19161_, _19160_, _19158_);
  and (_19162_, _03243_, _02108_);
  or (_19164_, _19162_, _19161_);
  nand (_19165_, _19164_, _17852_);
  and (_19166_, _02945_, _01965_);
  nor (_19167_, _19166_, _05342_);
  nand (_19168_, _19167_, _19165_);
  nor (_19169_, _18949_, \oc8051_golden_model_1.PSW [7]);
  nor (_19170_, _02107_, _05348_);
  nor (_19171_, _19170_, _05343_);
  not (_19172_, _19171_);
  nor (_19173_, _19172_, _19169_);
  nor (_19175_, _19173_, _01944_);
  and (_19176_, _19175_, _19168_);
  or (_19177_, _19176_, _18922_);
  nand (_19178_, _19177_, _05358_);
  and (_19179_, _05355_, _02108_);
  nor (_19180_, _19179_, _02654_);
  and (_19181_, _19180_, _19178_);
  and (_19182_, _02947_, _02654_);
  or (_19183_, _19182_, _03239_);
  nor (_19184_, _19183_, _19181_);
  and (_19186_, _03239_, _02108_);
  or (_19187_, _19186_, _19184_);
  nand (_19188_, _19187_, _17848_);
  and (_19189_, _02945_, _01957_);
  nor (_19190_, _19189_, _05367_);
  nand (_19191_, _19190_, _19188_);
  nor (_19192_, _18949_, _05348_);
  nor (_19193_, _02107_, \oc8051_golden_model_1.PSW [7]);
  nor (_19194_, _19193_, _05368_);
  not (_19195_, _19194_);
  nor (_19197_, _19195_, _19192_);
  nor (_19198_, _19197_, _05391_);
  and (_19199_, _19198_, _19191_);
  or (_19200_, _19199_, _18921_);
  nand (_19201_, _19200_, _05398_);
  and (_19202_, _05393_, _02108_);
  nor (_19203_, _19202_, _05396_);
  nand (_19204_, _19203_, _19201_);
  and (_19205_, _05396_, _02686_);
  nor (_19206_, _19205_, _03109_);
  and (_19208_, _19206_, _19204_);
  or (_19209_, _19208_, _18920_);
  nand (_19210_, _19209_, _05408_);
  and (_19211_, _02945_, _01936_);
  nor (_19212_, _19211_, _02653_);
  nand (_19213_, _19212_, _19210_);
  and (_19214_, _18936_, _05702_);
  nor (_19215_, _05702_, _02947_);
  or (_19216_, _19215_, _03267_);
  nor (_19217_, _19216_, _19214_);
  nor (_19219_, _19217_, _05412_);
  and (_19220_, _19219_, _19213_);
  or (_19221_, _19220_, _18919_);
  nand (_19222_, _19221_, _05728_);
  and (_19223_, _05720_, _02108_);
  nor (_19224_, _19223_, _05724_);
  nand (_19225_, _19224_, _19222_);
  and (_19226_, _05724_, _02686_);
  nor (_19227_, _19226_, _03108_);
  and (_19228_, _19227_, _19225_);
  and (_19230_, _04118_, _03108_);
  or (_19231_, _19230_, _19228_);
  nand (_19232_, _19231_, _05748_);
  and (_19233_, _02945_, _01899_);
  nor (_19234_, _19233_, _02647_);
  nand (_19235_, _19234_, _19232_);
  and (_19236_, _05702_, _02948_);
  nor (_19237_, _18935_, _05702_);
  nor (_19238_, _19237_, _19236_);
  and (_19239_, _19238_, _02647_);
  nor (_19241_, _19239_, _05764_);
  nand (_19242_, _19241_, _19235_);
  and (_19243_, _05764_, _02122_);
  nor (_19244_, _19243_, _03123_);
  and (_19245_, _19244_, _19242_);
  or (_19246_, _19245_, _18918_);
  nand (_19247_, _19246_, _05788_);
  and (_19248_, _05780_, _02686_);
  nor (_19249_, _19248_, _06742_);
  nand (_19250_, _19249_, _19247_);
  and (_19252_, _06742_, _02945_);
  nor (_19253_, _19252_, _02650_);
  nand (_19254_, _19253_, _19250_);
  and (_19255_, _19238_, _02650_);
  nor (_19256_, _19255_, _05826_);
  nand (_19257_, _19256_, _19254_);
  nor (_19258_, _05824_, _02686_);
  nor (_19259_, _19258_, _03121_);
  and (_19260_, _19259_, _19257_);
  or (_19261_, _19260_, _18917_);
  nand (_19263_, _19261_, _05848_);
  and (_19264_, _05840_, _02686_);
  nor (_19265_, _19264_, _18101_);
  nand (_19266_, _19265_, _19263_);
  and (_19267_, _18101_, _02945_);
  nor (_19268_, _19267_, _05862_);
  nand (_19269_, _19268_, _19266_);
  and (_19270_, _19269_, _18916_);
  nand (_19271_, _19270_, _27788_);
  or (_19272_, _27788_, \oc8051_golden_model_1.PC [3]);
  and (_19274_, _19272_, _27053_);
  and (_28961_, _19274_, _19271_);
  not (_19275_, \oc8051_golden_model_1.PC [4]);
  nor (_19276_, _01634_, _19275_);
  and (_19277_, _01634_, _19275_);
  nor (_19278_, _19277_, _19276_);
  and (_19279_, _19278_, _05862_);
  not (_19280_, _19279_);
  and (_19281_, _06742_, _02910_);
  and (_19282_, _02372_, _05348_);
  and (_19283_, _02518_, _02515_);
  nor (_19284_, _19283_, _02519_);
  and (_19285_, _19284_, \oc8051_golden_model_1.PSW [7]);
  or (_19286_, _19285_, _19282_);
  and (_19287_, _19286_, _05367_);
  and (_19288_, _02372_, _01953_);
  and (_19289_, _19284_, _02568_);
  or (_19290_, _19289_, _19288_);
  and (_19291_, _19290_, _02567_);
  and (_19292_, _02577_, _02373_);
  not (_19294_, _19278_);
  and (_19295_, _19294_, _05225_);
  and (_19296_, _02910_, _17956_);
  or (_19297_, _19296_, _03203_);
  nor (_19298_, _05177_, _02372_);
  and (_19299_, _03063_, _03060_);
  nor (_19300_, _19299_, _03064_);
  not (_19301_, _19300_);
  nor (_19302_, _19301_, _05157_);
  and (_19303_, _05157_, _02912_);
  nor (_19305_, _19303_, _19302_);
  or (_19306_, _19305_, _03387_);
  or (_19307_, _04987_, _02913_);
  or (_19308_, _19301_, _04985_);
  and (_19309_, _19308_, _02661_);
  and (_19310_, _19309_, _19307_);
  and (_19311_, _04540_, _02372_);
  and (_19312_, _19284_, _04537_);
  nor (_19313_, _19312_, _19311_);
  nand (_19314_, _19313_, _03406_);
  and (_19316_, _02910_, _04504_);
  and (_19317_, _04505_, _02373_);
  nor (_19318_, _19317_, _04520_);
  nor (_19319_, _04512_, _19275_);
  or (_19320_, _19319_, _04505_);
  nand (_19321_, _19320_, _19318_);
  or (_19322_, _19294_, _04521_);
  and (_19323_, _19322_, _01988_);
  and (_19324_, _19323_, _19321_);
  nor (_19325_, _19324_, _04510_);
  not (_19327_, _19325_);
  nor (_19328_, _19327_, _19316_);
  and (_19329_, _19278_, _04510_);
  or (_19330_, _19329_, _03154_);
  or (_19331_, _19330_, _19328_);
  nand (_19332_, _03154_, _02373_);
  and (_19333_, _19332_, _19331_);
  and (_19334_, _19333_, _18144_);
  and (_19335_, _19278_, _04502_);
  or (_19336_, _19335_, _19334_);
  and (_19339_, _19336_, _01998_);
  nor (_19340_, _02910_, _01998_);
  nor (_19341_, _19340_, _03406_);
  not (_19342_, _19341_);
  nor (_19343_, _19342_, _19339_);
  nor (_19344_, _19343_, _04545_);
  nand (_19345_, _19344_, _19314_);
  and (_19346_, _19345_, _02662_);
  or (_19347_, _19346_, _04992_);
  or (_19348_, _19347_, _19310_);
  or (_19350_, _19294_, _04996_);
  and (_19351_, _19350_, _03390_);
  nand (_19352_, _19351_, _19348_);
  and (_19353_, _03150_, _02373_);
  nor (_19354_, _19353_, _07558_);
  and (_19355_, _19354_, _19352_);
  nor (_19356_, _02910_, _01995_);
  or (_19357_, _19356_, _03162_);
  or (_19358_, _19357_, _19355_);
  and (_19359_, _03162_, _02373_);
  nor (_19362_, _19359_, _05000_);
  nand (_19363_, _19362_, _19358_);
  and (_19364_, _19278_, _05000_);
  nor (_19365_, _19364_, _03168_);
  nand (_19366_, _19365_, _19363_);
  and (_19367_, _03168_, _02373_);
  nor (_19368_, _19367_, _05009_);
  and (_19369_, _19368_, _19366_);
  and (_19370_, _19278_, _05009_);
  or (_19371_, _19370_, _03176_);
  or (_19373_, _19371_, _19369_);
  and (_19374_, _03176_, _02373_);
  nor (_19375_, _19374_, _17919_);
  and (_19376_, _19375_, _19373_);
  nor (_19377_, _02910_, _01990_);
  or (_19378_, _19377_, _19376_);
  nand (_19379_, _19378_, _03430_);
  and (_19380_, _03187_, _02372_);
  nor (_19381_, _19380_, _04498_);
  and (_19382_, _19381_, _19379_);
  and (_19385_, _04494_, _02912_);
  nor (_19386_, _19301_, _04494_);
  or (_19387_, _19386_, _19385_);
  nor (_19388_, _19387_, _04499_);
  or (_19389_, _19388_, _19382_);
  and (_19390_, _19389_, _03107_);
  and (_19391_, _04275_, _02912_);
  and (_19392_, _19300_, _04277_);
  or (_19393_, _19392_, _03107_);
  nor (_19394_, _19393_, _19391_);
  or (_19396_, _19394_, _19390_);
  or (_19397_, _19396_, _02664_);
  and (_19398_, _19397_, _19306_);
  or (_19399_, _19398_, _02673_);
  nand (_19400_, _02912_, _02630_);
  not (_19401_, _02630_);
  nand (_19402_, _19300_, _19401_);
  and (_19403_, _19402_, _19400_);
  or (_19404_, _19403_, _05024_);
  and (_19405_, _19404_, _19399_);
  or (_19408_, _19405_, _02598_);
  nand (_19409_, _19278_, _02598_);
  and (_19410_, _19409_, _19408_);
  nand (_19411_, _19410_, _05168_);
  and (_19412_, _03144_, _02373_);
  nor (_19413_, _19412_, _06664_);
  nand (_19414_, _19413_, _19411_);
  nor (_19415_, _02910_, _02000_);
  nor (_19416_, _19415_, _18254_);
  and (_19417_, _19416_, _19414_);
  or (_19419_, _19417_, _19298_);
  nand (_19420_, _19419_, _05186_);
  and (_19421_, _19294_, _05185_);
  nor (_19422_, _19421_, _03205_);
  nand (_19423_, _19422_, _19420_);
  and (_19424_, _03205_, _02372_);
  nor (_19425_, _19424_, _17956_);
  and (_19426_, _19425_, _19423_);
  nor (_19427_, _19426_, _19297_);
  and (_19428_, _03203_, _02372_);
  or (_19430_, _19428_, _19427_);
  nand (_19431_, _19430_, _05195_);
  and (_19432_, _19278_, _05194_);
  nor (_19433_, _19432_, _05199_);
  nand (_19434_, _19433_, _19431_);
  and (_19435_, _05199_, _02373_);
  nor (_19436_, _19435_, _02047_);
  and (_19437_, _19436_, _19434_);
  nor (_19438_, _19294_, _01985_);
  or (_19439_, _19438_, _03140_);
  nor (_19441_, _19439_, _19437_);
  and (_19442_, _03140_, _02373_);
  or (_19443_, _19442_, _19441_);
  nand (_19444_, _19443_, _07791_);
  and (_19445_, _02910_, _02025_);
  nor (_19446_, _19445_, _02670_);
  nand (_19447_, _19446_, _19444_);
  and (_19448_, _02912_, _02670_);
  nor (_19449_, _19448_, _05217_);
  nand (_19450_, _19449_, _19447_);
  and (_19452_, _05217_, _02373_);
  nor (_19453_, _19452_, _02024_);
  nand (_19454_, _19453_, _19450_);
  and (_19455_, _02912_, _02024_);
  nor (_19456_, _19455_, _05225_);
  and (_19457_, _19456_, _19454_);
  or (_19458_, _19457_, _19295_);
  nand (_19459_, _19458_, _03462_);
  and (_19460_, _03135_, _02373_);
  nor (_19461_, _19460_, _01960_);
  and (_19462_, _19461_, _19459_);
  nor (_19463_, _02910_, _17983_);
  or (_19464_, _19463_, _19462_);
  nand (_19465_, _19464_, _05234_);
  and (_19466_, _19284_, _05233_);
  nor (_19467_, _19466_, _02577_);
  and (_19468_, _19467_, _19465_);
  or (_19469_, _19468_, _19292_);
  nand (_19470_, _19469_, _05245_);
  and (_19471_, _02913_, _02575_);
  nor (_19473_, _19471_, _05243_);
  nand (_19474_, _19473_, _19470_);
  and (_19475_, _05243_, _02372_);
  nor (_19476_, _19475_, _02573_);
  nand (_19477_, _19476_, _19474_);
  and (_19478_, _05269_, _05266_);
  nor (_19479_, _19478_, _05270_);
  nor (_19480_, _19479_, _02574_);
  nor (_19481_, _19480_, _03134_);
  nand (_19482_, _19481_, _19477_);
  and (_19484_, _03134_, _02372_);
  nor (_19485_, _19484_, _01967_);
  nand (_19486_, _19485_, _19482_);
  and (_19487_, _02910_, _01967_);
  nor (_19488_, _19487_, _02567_);
  and (_19489_, _19488_, _19486_);
  or (_19490_, _19489_, _19291_);
  nand (_19491_, _19490_, _05298_);
  and (_19492_, _19278_, _05297_);
  nor (_19493_, _19492_, _05302_);
  nand (_19495_, _19493_, _19491_);
  and (_19496_, _05302_, _02373_);
  nor (_19497_, _19496_, _02656_);
  nand (_19498_, _19497_, _19495_);
  and (_19499_, _02912_, _02656_);
  nor (_19500_, _19499_, _03251_);
  and (_19501_, _19500_, _19498_);
  and (_19502_, _03251_, _02373_);
  or (_19503_, _19502_, _19501_);
  nand (_19504_, _19503_, _17855_);
  and (_19506_, _02910_, _01974_);
  nor (_19507_, _19506_, _05315_);
  nand (_19508_, _19507_, _19504_);
  nand (_19509_, _02372_, _02568_);
  nand (_19510_, _19284_, _01953_);
  and (_19511_, _19510_, _19509_);
  or (_19512_, _19511_, _05316_);
  nand (_19513_, _19512_, _19508_);
  nand (_19514_, _19513_, _05326_);
  and (_19515_, _19278_, _05325_);
  nor (_19517_, _19515_, _05329_);
  nand (_19518_, _19517_, _19514_);
  and (_19519_, _05329_, _02373_);
  nor (_19520_, _19519_, _02669_);
  nand (_19521_, _19520_, _19518_);
  and (_19522_, _02912_, _02669_);
  nor (_19523_, _19522_, _03243_);
  and (_19524_, _19523_, _19521_);
  and (_19525_, _03243_, _02373_);
  or (_19526_, _19525_, _19524_);
  nand (_19528_, _19526_, _17852_);
  and (_19529_, _02910_, _01965_);
  nor (_19530_, _19529_, _05342_);
  nand (_19531_, _19530_, _19528_);
  nand (_19532_, _02372_, \oc8051_golden_model_1.PSW [7]);
  nand (_19533_, _19284_, _05348_);
  and (_19534_, _19533_, _19532_);
  or (_19535_, _19534_, _05343_);
  nand (_19536_, _19535_, _19531_);
  nand (_19537_, _19536_, _01945_);
  and (_19539_, _19278_, _01944_);
  nor (_19540_, _19539_, _05355_);
  nand (_19541_, _19540_, _19537_);
  and (_19542_, _05355_, _02373_);
  nor (_19543_, _19542_, _02654_);
  nand (_19544_, _19543_, _19541_);
  and (_19545_, _02912_, _02654_);
  nor (_19546_, _19545_, _03239_);
  and (_19547_, _19546_, _19544_);
  and (_19548_, _03239_, _02373_);
  or (_19550_, _19548_, _19547_);
  nand (_19551_, _19550_, _17848_);
  and (_19552_, _02910_, _01957_);
  nor (_19553_, _19552_, _05367_);
  and (_19554_, _19553_, _19551_);
  or (_19555_, _19554_, _19287_);
  nand (_19556_, _19555_, _05389_);
  nor (_19557_, _19294_, _05389_);
  nor (_19558_, _19557_, _05393_);
  nand (_19559_, _19558_, _19556_);
  and (_19561_, _05393_, _02373_);
  nor (_19562_, _19561_, _05396_);
  nand (_19563_, _19562_, _19559_);
  and (_19564_, _19278_, _05396_);
  nor (_19565_, _19564_, _03109_);
  and (_19566_, _19565_, _19563_);
  and (_19567_, _04014_, _03109_);
  or (_19568_, _19567_, _19566_);
  nand (_19569_, _19568_, _05408_);
  and (_19570_, _02910_, _01936_);
  nor (_19572_, _19570_, _02653_);
  and (_19573_, _19572_, _19569_);
  nor (_19574_, _05702_, _02913_);
  and (_19575_, _19300_, _05702_);
  nor (_19576_, _19575_, _19574_);
  nor (_19577_, _19576_, _03267_);
  or (_19578_, _19577_, _19573_);
  nand (_19579_, _19578_, _01930_);
  nor (_19580_, _19294_, _01930_);
  nor (_19581_, _19580_, _05720_);
  nand (_19583_, _19581_, _19579_);
  and (_19584_, _05720_, _02373_);
  nor (_19585_, _19584_, _05724_);
  nand (_19586_, _19585_, _19583_);
  and (_19587_, _19278_, _05724_);
  nor (_19588_, _19587_, _03108_);
  nand (_19589_, _19588_, _19586_);
  and (_19590_, _04014_, _03108_);
  nor (_19591_, _19590_, _01899_);
  nand (_19592_, _19591_, _19589_);
  nor (_19594_, _02910_, _05748_);
  nor (_19595_, _19594_, _02647_);
  nand (_19596_, _19595_, _19592_);
  and (_19597_, _05702_, _02913_);
  nor (_19598_, _19300_, _05702_);
  nor (_19599_, _19598_, _19597_);
  nor (_19600_, _19599_, _03125_);
  nor (_19601_, _19600_, _05764_);
  nand (_19602_, _19601_, _19596_);
  and (_19603_, _19278_, _05764_);
  nor (_19605_, _19603_, _03123_);
  nand (_19606_, _19605_, _19602_);
  and (_19607_, _03123_, _02373_);
  nor (_19608_, _19607_, _05780_);
  nand (_19609_, _19608_, _19606_);
  and (_19610_, _19278_, _05780_);
  nor (_19611_, _19610_, _06742_);
  and (_19612_, _19611_, _19609_);
  or (_19613_, _19612_, _19281_);
  nand (_19614_, _19613_, _03122_);
  nor (_19616_, _19599_, _03122_);
  nor (_19617_, _19616_, _05826_);
  nand (_19618_, _19617_, _19614_);
  nor (_19619_, _19294_, _05824_);
  nor (_19620_, _19619_, _03121_);
  nand (_19621_, _19620_, _19618_);
  and (_19622_, _03121_, _02373_);
  nor (_19623_, _19622_, _05840_);
  nand (_19624_, _19623_, _19621_);
  and (_19625_, _19278_, _05840_);
  nor (_19627_, _19625_, _18101_);
  nand (_19628_, _19627_, _19624_);
  and (_19629_, _18101_, _02910_);
  nor (_19630_, _19629_, _05862_);
  nand (_19631_, _19630_, _19628_);
  and (_19632_, _19631_, _19280_);
  nand (_19633_, _19632_, _27788_);
  or (_19634_, _27788_, \oc8051_golden_model_1.PC [4]);
  and (_19635_, _19634_, _27053_);
  and (_28964_, _19635_, _19633_);
  nor (_19636_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_19637_, _02336_, _01647_);
  nor (_19638_, _19637_, _19636_);
  and (_19639_, _19638_, _05862_);
  not (_19640_, _19639_);
  and (_19641_, _03121_, _02336_);
  and (_19642_, _03123_, _02336_);
  nor (_19643_, _19638_, _01930_);
  nor (_19644_, _19638_, _05389_);
  not (_19645_, _19638_);
  and (_19647_, _19645_, _01944_);
  and (_19648_, _19645_, _05325_);
  and (_19649_, _19645_, _05297_);
  and (_19650_, _02577_, _02337_);
  and (_19651_, _03140_, _02337_);
  and (_19652_, _19645_, _05194_);
  nor (_19653_, _05177_, _02336_);
  or (_19654_, _02879_, _02878_);
  not (_19655_, _19654_);
  nor (_19656_, _19655_, _03065_);
  and (_19658_, _19655_, _03065_);
  nor (_19659_, _19658_, _19656_);
  nor (_19660_, _19659_, _05157_);
  and (_19661_, _05157_, _02876_);
  nor (_19662_, _19661_, _19660_);
  or (_19663_, _19662_, _03387_);
  and (_19664_, _04494_, _02876_);
  nor (_19665_, _19659_, _04494_);
  or (_19666_, _19665_, _19664_);
  nor (_19667_, _19666_, _04499_);
  and (_19669_, _19659_, _04987_);
  and (_19670_, _04985_, _02877_);
  nor (_19671_, _19670_, _19669_);
  or (_19672_, _19671_, _02662_);
  and (_19673_, _04540_, _02336_);
  or (_19674_, _02338_, _02339_);
  and (_19675_, _19674_, _02520_);
  nor (_19676_, _19674_, _02520_);
  nor (_19677_, _19676_, _19675_);
  and (_19678_, _19677_, _04537_);
  or (_19680_, _19678_, _19673_);
  nor (_19681_, _19680_, _04539_);
  nor (_19682_, _02873_, _01988_);
  and (_19683_, _04505_, _02337_);
  nor (_19684_, _19683_, _04520_);
  not (_19685_, _04512_);
  and (_19686_, _19685_, \oc8051_golden_model_1.PC [5]);
  or (_19687_, _19686_, _04505_);
  and (_19688_, _19687_, _19684_);
  nor (_19689_, _19645_, _04521_);
  or (_19691_, _19689_, _04510_);
  or (_19692_, _19691_, _19688_);
  and (_19693_, _19692_, _01988_);
  nor (_19694_, _19693_, _19682_);
  and (_19695_, _19645_, _04510_);
  nor (_19696_, _19695_, _03154_);
  not (_19697_, _19696_);
  nor (_19698_, _19697_, _19694_);
  and (_19699_, _03154_, _02336_);
  or (_19700_, _19699_, _19698_);
  and (_19702_, _19700_, _18144_);
  and (_19703_, _19638_, _04502_);
  or (_19704_, _19703_, _19702_);
  and (_19705_, _19704_, _01998_);
  nor (_19706_, _02873_, _01998_);
  nor (_19707_, _19706_, _03406_);
  not (_19708_, _19707_);
  nor (_19709_, _19708_, _19705_);
  or (_19710_, _19709_, _04545_);
  nor (_19711_, _19710_, _19681_);
  and (_19713_, _19638_, _04545_);
  or (_19714_, _19713_, _02661_);
  or (_19715_, _19714_, _19711_);
  and (_19716_, _19715_, _19672_);
  nor (_19717_, _19716_, _04992_);
  and (_19718_, _19645_, _04992_);
  nor (_19719_, _19718_, _03150_);
  not (_19720_, _19719_);
  or (_19721_, _19720_, _19717_);
  and (_19722_, _03150_, _02336_);
  nor (_19724_, _19722_, _07558_);
  nand (_19725_, _19724_, _19721_);
  and (_19726_, _02873_, _07558_);
  nor (_19727_, _19726_, _03162_);
  nand (_19728_, _19727_, _19725_);
  and (_19729_, _03162_, _02336_);
  nor (_19730_, _19729_, _05000_);
  nand (_19731_, _19730_, _19728_);
  and (_19732_, _19645_, _05000_);
  nor (_19733_, _19732_, _03168_);
  nand (_19735_, _19733_, _19731_);
  and (_19736_, _03168_, _02336_);
  nor (_19737_, _19736_, _05009_);
  nand (_19738_, _19737_, _19735_);
  and (_19739_, _19645_, _05009_);
  nor (_19740_, _19739_, _03176_);
  nand (_19741_, _19740_, _19738_);
  and (_19742_, _03176_, _02336_);
  nor (_19743_, _19742_, _17919_);
  nand (_19744_, _19743_, _19741_);
  and (_19746_, _02873_, _17919_);
  nor (_19747_, _19746_, _03187_);
  nand (_19748_, _19747_, _19744_);
  and (_19749_, _03187_, _02336_);
  nor (_19750_, _19749_, _04498_);
  and (_19751_, _19750_, _19748_);
  or (_19752_, _19751_, _19667_);
  and (_19753_, _19752_, _03107_);
  and (_19754_, _04275_, _02876_);
  not (_19755_, _19659_);
  and (_19757_, _19755_, _04277_);
  or (_19758_, _19757_, _03107_);
  nor (_19759_, _19758_, _19754_);
  or (_19760_, _19759_, _19753_);
  or (_19761_, _19760_, _02664_);
  and (_19762_, _19761_, _19663_);
  or (_19763_, _19762_, _02673_);
  nand (_19764_, _02876_, _02630_);
  or (_19765_, _19659_, _02630_);
  and (_19766_, _19765_, _19764_);
  or (_19768_, _19766_, _05024_);
  and (_19769_, _19768_, _19763_);
  or (_19770_, _19769_, _02598_);
  nand (_19771_, _19638_, _02598_);
  and (_19772_, _19771_, _19770_);
  nand (_19773_, _19772_, _05168_);
  and (_19774_, _03144_, _02337_);
  nor (_19775_, _19774_, _06664_);
  nand (_19776_, _19775_, _19773_);
  nor (_19777_, _02873_, _02000_);
  nor (_19779_, _19777_, _18254_);
  and (_19780_, _19779_, _19776_);
  or (_19781_, _19780_, _19653_);
  nand (_19782_, _19781_, _05186_);
  and (_19783_, _19645_, _05185_);
  nor (_19784_, _19783_, _03205_);
  nand (_19785_, _19784_, _19782_);
  and (_19786_, _03205_, _02336_);
  nor (_19787_, _19786_, _17956_);
  nand (_19788_, _19787_, _19785_);
  and (_19790_, _02873_, _17956_);
  nor (_19791_, _19790_, _03203_);
  nand (_19792_, _19791_, _19788_);
  and (_19793_, _03203_, _02336_);
  nor (_19794_, _19793_, _05194_);
  and (_19795_, _19794_, _19792_);
  or (_19796_, _19795_, _19652_);
  nand (_19797_, _19796_, _05203_);
  and (_19798_, _05199_, _02337_);
  nor (_19799_, _19798_, _02047_);
  nand (_19801_, _19799_, _19797_);
  nor (_19802_, _19645_, _01985_);
  nor (_19803_, _19802_, _03140_);
  and (_19804_, _19803_, _19801_);
  or (_19805_, _19804_, _19651_);
  nand (_19806_, _19805_, _07791_);
  and (_19807_, _02873_, _02025_);
  nor (_19808_, _19807_, _02670_);
  nand (_19809_, _19808_, _19806_);
  and (_19810_, _02876_, _02670_);
  nor (_19811_, _19810_, _05217_);
  nand (_19812_, _19811_, _19809_);
  and (_19813_, _05217_, _02337_);
  nor (_19814_, _19813_, _02024_);
  nand (_19815_, _19814_, _19812_);
  and (_19816_, _02876_, _02024_);
  nor (_19817_, _19816_, _05225_);
  nand (_19818_, _19817_, _19815_);
  and (_19819_, _19645_, _05225_);
  nor (_19820_, _19819_, _03135_);
  nand (_19822_, _19820_, _19818_);
  and (_19823_, _03135_, _02336_);
  nor (_19824_, _19823_, _01960_);
  nand (_19825_, _19824_, _19822_);
  and (_19826_, _02873_, _01960_);
  nor (_19827_, _19826_, _05233_);
  nand (_19828_, _19827_, _19825_);
  and (_19829_, _19677_, _05233_);
  nor (_19830_, _19829_, _02577_);
  and (_19831_, _19830_, _19828_);
  or (_19833_, _19831_, _19650_);
  nand (_19834_, _19833_, _05245_);
  and (_19835_, _02877_, _02575_);
  nor (_19836_, _19835_, _05243_);
  nand (_19837_, _19836_, _19834_);
  and (_19838_, _05243_, _02336_);
  nor (_19839_, _19838_, _02573_);
  nand (_19840_, _19839_, _19837_);
  and (_19841_, _05271_, _05264_);
  nor (_19842_, _19841_, _05272_);
  nor (_19844_, _19842_, _02574_);
  nor (_19845_, _19844_, _03134_);
  nand (_19846_, _19845_, _19840_);
  and (_19847_, _03134_, _02336_);
  nor (_19848_, _19847_, _01967_);
  nand (_19849_, _19848_, _19846_);
  and (_19850_, _02873_, _01967_);
  nor (_19851_, _19850_, _02567_);
  nand (_19852_, _19851_, _19849_);
  and (_19853_, _02336_, _01953_);
  and (_19855_, _19677_, _02568_);
  or (_19856_, _19855_, _19853_);
  and (_19857_, _19856_, _02567_);
  nor (_19858_, _19857_, _05297_);
  and (_19859_, _19858_, _19852_);
  or (_19860_, _19859_, _19649_);
  nand (_19861_, _19860_, _05306_);
  and (_19862_, _05302_, _02337_);
  nor (_19863_, _19862_, _02656_);
  nand (_19864_, _19863_, _19861_);
  and (_19866_, _02876_, _02656_);
  nor (_19867_, _19866_, _03251_);
  and (_19868_, _19867_, _19864_);
  and (_19869_, _03251_, _02337_);
  or (_19870_, _19869_, _19868_);
  nand (_19871_, _19870_, _17855_);
  and (_19872_, _02873_, _01974_);
  nor (_19873_, _19872_, _05315_);
  nand (_19874_, _19873_, _19871_);
  and (_19875_, _02336_, _02568_);
  and (_19877_, _19677_, _01953_);
  or (_19878_, _19877_, _19875_);
  and (_19879_, _19878_, _05315_);
  nor (_19880_, _19879_, _05325_);
  and (_19881_, _19880_, _19874_);
  or (_19882_, _19881_, _19648_);
  nand (_19883_, _19882_, _05333_);
  and (_19884_, _05329_, _02337_);
  nor (_19885_, _19884_, _02669_);
  nand (_19886_, _19885_, _19883_);
  and (_19888_, _02876_, _02669_);
  nor (_19889_, _19888_, _03243_);
  and (_19890_, _19889_, _19886_);
  and (_19891_, _03243_, _02337_);
  or (_19892_, _19891_, _19890_);
  nand (_19893_, _19892_, _17852_);
  and (_19894_, _02873_, _01965_);
  nor (_19895_, _19894_, _05342_);
  nand (_19896_, _19895_, _19893_);
  nor (_19897_, _19677_, \oc8051_golden_model_1.PSW [7]);
  nor (_19899_, _02336_, _05348_);
  nor (_19900_, _19899_, _05343_);
  not (_19901_, _19900_);
  nor (_19902_, _19901_, _19897_);
  nor (_19903_, _19902_, _01944_);
  and (_19904_, _19903_, _19896_);
  or (_19905_, _19904_, _19647_);
  nand (_19906_, _19905_, _05358_);
  and (_19907_, _05355_, _02337_);
  nor (_19908_, _19907_, _02654_);
  nand (_19910_, _19908_, _19906_);
  and (_19911_, _02876_, _02654_);
  nor (_19912_, _19911_, _03239_);
  and (_19913_, _19912_, _19910_);
  and (_19914_, _03239_, _02337_);
  or (_19915_, _19914_, _19913_);
  nand (_19916_, _19915_, _17848_);
  and (_19917_, _02873_, _01957_);
  nor (_19918_, _19917_, _05367_);
  nand (_19919_, _19918_, _19916_);
  nor (_19921_, _19677_, _05348_);
  nor (_19922_, _02336_, \oc8051_golden_model_1.PSW [7]);
  nor (_19923_, _19922_, _05368_);
  not (_19924_, _19923_);
  nor (_19925_, _19924_, _19921_);
  nor (_19926_, _19925_, _05391_);
  and (_19927_, _19926_, _19919_);
  or (_19928_, _19927_, _19644_);
  nand (_19929_, _19928_, _05398_);
  and (_19930_, _05393_, _02337_);
  nor (_19932_, _19930_, _05396_);
  nand (_19933_, _19932_, _19929_);
  and (_19934_, _19638_, _05396_);
  nor (_19935_, _19934_, _03109_);
  and (_19936_, _19935_, _19933_);
  and (_19937_, _03906_, _03109_);
  or (_19938_, _19937_, _19936_);
  nand (_19939_, _19938_, _05408_);
  and (_19940_, _02873_, _01936_);
  nor (_19941_, _19940_, _02653_);
  nand (_19943_, _19941_, _19939_);
  and (_19944_, _19659_, _05702_);
  nor (_19945_, _05702_, _02876_);
  or (_19946_, _19945_, _03267_);
  nor (_19947_, _19946_, _19944_);
  nor (_19948_, _19947_, _05412_);
  and (_19949_, _19948_, _19943_);
  or (_19950_, _19949_, _19643_);
  nand (_19951_, _19950_, _05728_);
  and (_19952_, _05720_, _02337_);
  nor (_19954_, _19952_, _05724_);
  nand (_19955_, _19954_, _19951_);
  and (_19956_, _19638_, _05724_);
  nor (_19957_, _19956_, _03108_);
  and (_19958_, _19957_, _19955_);
  and (_19959_, _03906_, _03108_);
  or (_19960_, _19959_, _19958_);
  nand (_19961_, _19960_, _05748_);
  and (_19962_, _02873_, _01899_);
  nor (_19963_, _19962_, _02647_);
  nand (_19965_, _19963_, _19961_);
  and (_19966_, _05702_, _02877_);
  nor (_19967_, _19755_, _05702_);
  nor (_19968_, _19967_, _19966_);
  and (_19969_, _19968_, _02647_);
  nor (_19970_, _19969_, _05764_);
  nand (_19971_, _19970_, _19965_);
  and (_19972_, _19645_, _05764_);
  nor (_19973_, _19972_, _03123_);
  and (_19974_, _19973_, _19971_);
  or (_19976_, _19974_, _19642_);
  nand (_19977_, _19976_, _05788_);
  and (_19978_, _19638_, _05780_);
  nor (_19979_, _19978_, _06742_);
  nand (_19980_, _19979_, _19977_);
  and (_19981_, _06742_, _02873_);
  nor (_19982_, _19981_, _02650_);
  nand (_19983_, _19982_, _19980_);
  and (_19984_, _19968_, _02650_);
  nor (_19985_, _19984_, _05826_);
  nand (_19987_, _19985_, _19983_);
  nor (_19988_, _19638_, _05824_);
  nor (_19989_, _19988_, _03121_);
  and (_19990_, _19989_, _19987_);
  or (_19991_, _19990_, _19641_);
  nand (_19992_, _19991_, _05848_);
  and (_19993_, _19638_, _05840_);
  nor (_19994_, _19993_, _18101_);
  nand (_19995_, _19994_, _19992_);
  and (_19996_, _18101_, _02873_);
  nor (_19998_, _19996_, _05862_);
  nand (_19999_, _19998_, _19995_);
  and (_20000_, _19999_, _19640_);
  nand (_20001_, _20000_, _27788_);
  or (_20002_, _27788_, \oc8051_golden_model_1.PC [5]);
  and (_20003_, _20002_, _27053_);
  and (_28965_, _20003_, _20001_);
  nor (_20004_, _01902_, \oc8051_golden_model_1.PC [6]);
  nor (_20005_, _20004_, _01903_);
  and (_20006_, _20005_, _05862_);
  and (_20008_, _06742_, _02834_);
  and (_20009_, _05157_, _02837_);
  and (_20010_, _03067_, _02842_);
  nor (_20011_, _20010_, _03068_);
  not (_20012_, _20011_);
  nor (_20013_, _20012_, _05157_);
  nor (_20014_, _20013_, _20009_);
  or (_20015_, _20014_, _03387_);
  or (_20016_, _04987_, _02838_);
  or (_20017_, _20012_, _04985_);
  and (_20019_, _20017_, _02661_);
  and (_20020_, _20019_, _20016_);
  and (_20021_, _04540_, _02298_);
  nor (_20022_, _02522_, _02302_);
  nor (_20023_, _20022_, _02523_);
  and (_20024_, _20023_, _04537_);
  nor (_20025_, _20024_, _20021_);
  nand (_20026_, _20025_, _03406_);
  and (_20027_, _03154_, _02299_);
  and (_20028_, _02834_, _04504_);
  nor (_20030_, _04512_, \oc8051_golden_model_1.PC [6]);
  or (_20031_, _20030_, _04505_);
  and (_20032_, _04505_, _02298_);
  nor (_20033_, _20032_, _04520_);
  and (_20034_, _20033_, _20031_);
  nor (_20035_, _20005_, _04521_);
  or (_20036_, _20035_, _04510_);
  or (_20037_, _20036_, _20034_);
  and (_20038_, _20037_, _01988_);
  nor (_20039_, _20038_, _20028_);
  and (_20041_, _20005_, _04510_);
  nor (_20042_, _20041_, _03154_);
  not (_20043_, _20042_);
  nor (_20044_, _20043_, _20039_);
  nor (_20045_, _20044_, _20027_);
  and (_20046_, _20045_, _18144_);
  and (_20047_, _20005_, _04502_);
  or (_20048_, _20047_, _20046_);
  and (_20049_, _20048_, _01998_);
  nor (_20050_, _02834_, _01998_);
  nor (_20052_, _20050_, _03406_);
  not (_20053_, _20052_);
  nor (_20054_, _20053_, _20049_);
  nor (_20055_, _20054_, _04545_);
  nand (_20056_, _20055_, _20026_);
  and (_20057_, _20056_, _02662_);
  or (_20058_, _20057_, _04992_);
  or (_20059_, _20058_, _20020_);
  not (_20060_, _20005_);
  or (_20061_, _20060_, _04996_);
  and (_20063_, _20061_, _03390_);
  nand (_20064_, _20063_, _20059_);
  and (_20065_, _03150_, _02299_);
  nor (_20066_, _20065_, _07558_);
  and (_20067_, _20066_, _20064_);
  nor (_20068_, _02834_, _01995_);
  or (_20069_, _20068_, _03162_);
  or (_20070_, _20069_, _20067_);
  and (_20071_, _03162_, _02299_);
  nor (_20072_, _20071_, _05000_);
  nand (_20074_, _20072_, _20070_);
  and (_20075_, _20005_, _05000_);
  nor (_20076_, _20075_, _03168_);
  nand (_20077_, _20076_, _20074_);
  and (_20078_, _03168_, _02299_);
  nor (_20079_, _20078_, _05009_);
  and (_20080_, _20079_, _20077_);
  and (_20081_, _20005_, _05009_);
  or (_20082_, _20081_, _03176_);
  or (_20083_, _20082_, _20080_);
  and (_20085_, _03176_, _02299_);
  nor (_20086_, _20085_, _17919_);
  and (_20087_, _20086_, _20083_);
  nor (_20088_, _02834_, _01990_);
  or (_20089_, _20088_, _20087_);
  nand (_20090_, _20089_, _03430_);
  and (_20091_, _03187_, _02298_);
  nor (_20092_, _20091_, _04498_);
  and (_20093_, _20092_, _20090_);
  and (_20094_, _04494_, _02837_);
  nor (_20096_, _20012_, _04494_);
  or (_20097_, _20096_, _20094_);
  nor (_20098_, _20097_, _04499_);
  or (_20099_, _20098_, _20093_);
  and (_20100_, _20099_, _03107_);
  and (_20101_, _04275_, _02837_);
  and (_20102_, _20011_, _04277_);
  or (_20103_, _20102_, _03107_);
  nor (_20104_, _20103_, _20101_);
  or (_20105_, _20104_, _20100_);
  or (_20107_, _20105_, _02664_);
  and (_20108_, _20107_, _20015_);
  or (_20109_, _20108_, _02673_);
  nand (_20110_, _02837_, _02630_);
  nand (_20111_, _20011_, _19401_);
  and (_20112_, _20111_, _20110_);
  or (_20113_, _20112_, _05024_);
  and (_20114_, _20113_, _20109_);
  or (_20115_, _20114_, _02598_);
  nand (_20116_, _20005_, _02598_);
  and (_20118_, _20116_, _20115_);
  nand (_20119_, _20118_, _05168_);
  and (_20120_, _03144_, _02299_);
  nor (_20121_, _20120_, _06664_);
  nand (_20122_, _20121_, _20119_);
  nor (_20123_, _02834_, _02000_);
  nor (_20124_, _20123_, _18254_);
  and (_20125_, _20124_, _20122_);
  nor (_20126_, _05177_, _02298_);
  or (_20127_, _20126_, _20125_);
  nand (_20129_, _20127_, _05186_);
  and (_20130_, _20060_, _05185_);
  nor (_20131_, _20130_, _03205_);
  nand (_20132_, _20131_, _20129_);
  and (_20133_, _03205_, _02298_);
  nor (_20134_, _20133_, _17956_);
  nand (_20135_, _20134_, _20132_);
  and (_20136_, _02834_, _17956_);
  nor (_20137_, _20136_, _03203_);
  nand (_20138_, _20137_, _20135_);
  and (_20140_, _03203_, _02298_);
  nor (_20141_, _20140_, _05194_);
  nand (_20142_, _20141_, _20138_);
  and (_20143_, _20060_, _05194_);
  nor (_20144_, _20143_, _05199_);
  and (_20145_, _20144_, _20142_);
  and (_20146_, _05199_, _02298_);
  or (_20147_, _20146_, _20145_);
  and (_20148_, _20147_, _01985_);
  nor (_20149_, _20060_, _01985_);
  or (_20151_, _20149_, _03140_);
  or (_20152_, _20151_, _20148_);
  and (_20153_, _03140_, _02299_);
  nor (_20154_, _20153_, _02025_);
  nand (_20155_, _20154_, _20152_);
  nor (_20156_, _02834_, _07791_);
  nor (_20157_, _20156_, _02670_);
  nand (_20158_, _20157_, _20155_);
  and (_20159_, _02838_, _02670_);
  nor (_20160_, _20159_, _05217_);
  nand (_20162_, _20160_, _20158_);
  and (_20163_, _05217_, _02298_);
  nor (_20164_, _20163_, _02024_);
  nand (_20165_, _20164_, _20162_);
  and (_20166_, _02838_, _02024_);
  nor (_20167_, _20166_, _05225_);
  nand (_20168_, _20167_, _20165_);
  and (_20169_, _20005_, _05225_);
  nor (_20170_, _20169_, _03135_);
  nand (_20171_, _20170_, _20168_);
  and (_20173_, _03135_, _02299_);
  nor (_20174_, _20173_, _01960_);
  nand (_20175_, _20174_, _20171_);
  nor (_20176_, _02834_, _17983_);
  nor (_20177_, _20176_, _05233_);
  and (_20178_, _20177_, _20175_);
  nor (_20179_, _20023_, _05234_);
  or (_20180_, _20179_, _20178_);
  or (_20181_, _20180_, _02577_);
  nand (_20182_, _02577_, _02298_);
  and (_20184_, _20182_, _05245_);
  nand (_20185_, _20184_, _20181_);
  and (_20186_, _02838_, _02575_);
  nor (_20187_, _20186_, _05243_);
  nand (_20188_, _20187_, _20185_);
  and (_20189_, _05243_, _02298_);
  nor (_20190_, _20189_, _02573_);
  nand (_20191_, _20190_, _20188_);
  and (_20192_, _05273_, _05260_);
  nor (_20193_, _20192_, _05274_);
  nor (_20195_, _20193_, _02574_);
  nor (_20196_, _20195_, _03134_);
  nand (_20197_, _20196_, _20191_);
  and (_20198_, _03134_, _02298_);
  nor (_20199_, _20198_, _01967_);
  nand (_20200_, _20199_, _20197_);
  and (_20201_, _02834_, _01967_);
  nor (_20202_, _20201_, _02567_);
  nand (_20203_, _20202_, _20200_);
  and (_20204_, _02298_, _01953_);
  and (_20206_, _20023_, _02568_);
  or (_20207_, _20206_, _20204_);
  and (_20208_, _20207_, _02567_);
  nor (_20209_, _20208_, _05297_);
  nand (_20210_, _20209_, _20203_);
  and (_20211_, _20060_, _05297_);
  nor (_20212_, _20211_, _05302_);
  nand (_20213_, _20212_, _20210_);
  and (_20214_, _05302_, _02298_);
  nor (_20215_, _20214_, _02656_);
  and (_20217_, _20215_, _20213_);
  and (_20218_, _02838_, _02656_);
  or (_20219_, _20218_, _20217_);
  nand (_20220_, _20219_, _03252_);
  and (_20221_, _03251_, _02299_);
  nor (_20222_, _20221_, _01974_);
  and (_20223_, _20222_, _20220_);
  nor (_20224_, _02834_, _17855_);
  or (_20225_, _20224_, _20223_);
  nand (_20226_, _20225_, _05316_);
  and (_20228_, _02298_, _02568_);
  and (_20229_, _20023_, _01953_);
  or (_20230_, _20229_, _20228_);
  and (_20231_, _20230_, _05315_);
  nor (_20232_, _20231_, _05325_);
  nand (_20233_, _20232_, _20226_);
  and (_20234_, _20060_, _05325_);
  nor (_20235_, _20234_, _05329_);
  nand (_20236_, _20235_, _20233_);
  and (_20237_, _05329_, _02298_);
  nor (_20239_, _20237_, _02669_);
  and (_20240_, _20239_, _20236_);
  and (_20241_, _02838_, _02669_);
  or (_20242_, _20241_, _20240_);
  nand (_20243_, _20242_, _03244_);
  and (_20244_, _03243_, _02299_);
  nor (_20245_, _20244_, _01965_);
  and (_20246_, _20245_, _20243_);
  nor (_20247_, _02834_, _17852_);
  or (_20248_, _20247_, _20246_);
  nand (_20250_, _20248_, _05343_);
  nor (_20251_, _20023_, \oc8051_golden_model_1.PSW [7]);
  nor (_20252_, _02298_, _05348_);
  nor (_20253_, _20252_, _05343_);
  not (_20254_, _20253_);
  nor (_20255_, _20254_, _20251_);
  nor (_20256_, _20255_, _01944_);
  nand (_20257_, _20256_, _20250_);
  and (_20258_, _20060_, _01944_);
  nor (_20259_, _20258_, _05355_);
  nand (_20261_, _20259_, _20257_);
  and (_20262_, _05355_, _02298_);
  nor (_20263_, _20262_, _02654_);
  and (_20264_, _20263_, _20261_);
  and (_20265_, _02838_, _02654_);
  or (_20266_, _20265_, _20264_);
  nand (_20267_, _20266_, _05883_);
  and (_20268_, _03239_, _02299_);
  nor (_20269_, _20268_, _01957_);
  and (_20270_, _20269_, _20267_);
  nor (_20272_, _02834_, _17848_);
  or (_20273_, _20272_, _20270_);
  nand (_20274_, _20273_, _05368_);
  nor (_20275_, _20023_, _05348_);
  nor (_20276_, _02298_, \oc8051_golden_model_1.PSW [7]);
  nor (_20277_, _20276_, _05368_);
  not (_20278_, _20277_);
  nor (_20279_, _20278_, _20275_);
  nor (_20280_, _20279_, _05391_);
  nand (_20281_, _20280_, _20274_);
  nor (_20283_, _20005_, _05389_);
  nor (_20284_, _20283_, _05393_);
  and (_20285_, _20284_, _20281_);
  and (_20286_, _05393_, _02298_);
  or (_20287_, _20286_, _20285_);
  and (_20288_, _20287_, _05397_);
  and (_20289_, _20005_, _05396_);
  or (_20290_, _20289_, _20288_);
  nand (_20291_, _20290_, _06612_);
  and (_20292_, _03960_, _03109_);
  nor (_20294_, _20292_, _01936_);
  nand (_20295_, _20294_, _20291_);
  and (_20296_, _02834_, _01936_);
  nor (_20297_, _20296_, _02653_);
  nand (_20298_, _20297_, _20295_);
  and (_20299_, _20012_, _05702_);
  nor (_20300_, _05702_, _02837_);
  or (_20301_, _20300_, _03267_);
  nor (_20302_, _20301_, _20299_);
  nor (_20303_, _20302_, _05412_);
  nand (_20305_, _20303_, _20298_);
  nor (_20306_, _20005_, _01930_);
  nor (_20307_, _20306_, _05720_);
  and (_20308_, _20307_, _20305_);
  and (_20309_, _05720_, _02298_);
  or (_20310_, _20309_, _20308_);
  nand (_20311_, _20310_, _05726_);
  and (_20312_, _20005_, _05724_);
  nor (_20313_, _20312_, _03108_);
  nand (_20314_, _20313_, _20311_);
  and (_20316_, _03958_, _03108_);
  nor (_20317_, _20316_, _01899_);
  nand (_20318_, _20317_, _20314_);
  nor (_20319_, _02834_, _05748_);
  nor (_20320_, _20319_, _02647_);
  and (_20321_, _20320_, _20318_);
  nor (_20322_, _20011_, _05702_);
  and (_20323_, _05702_, _02838_);
  nor (_20324_, _20323_, _20322_);
  nor (_20325_, _20324_, _03125_);
  or (_20327_, _20325_, _20321_);
  and (_20328_, _20327_, _05770_);
  and (_20329_, _20060_, _05764_);
  or (_20330_, _20329_, _20328_);
  nand (_20331_, _20330_, _03124_);
  and (_20332_, _03123_, _02299_);
  nor (_20333_, _20332_, _05780_);
  nand (_20334_, _20333_, _20331_);
  and (_20335_, _20005_, _05780_);
  nor (_20336_, _20335_, _06742_);
  and (_20338_, _20336_, _20334_);
  or (_20339_, _20338_, _20008_);
  nand (_20340_, _20339_, _03122_);
  nor (_20341_, _20324_, _03122_);
  nor (_20342_, _20341_, _05826_);
  nand (_20343_, _20342_, _20340_);
  nor (_20344_, _20060_, _05824_);
  nor (_20345_, _20344_, _03121_);
  nand (_20346_, _20345_, _20343_);
  and (_20347_, _03121_, _02299_);
  nor (_20349_, _20347_, _05840_);
  nand (_20350_, _20349_, _20346_);
  and (_20351_, _20005_, _05840_);
  nor (_20352_, _20351_, _18101_);
  nand (_20353_, _20352_, _20350_);
  and (_20354_, _18101_, _02834_);
  nor (_20355_, _20354_, _05862_);
  and (_20356_, _20355_, _20353_);
  or (_20357_, _20356_, _20006_);
  or (_20358_, _20357_, _27789_);
  or (_20360_, _27788_, \oc8051_golden_model_1.PC [6]);
  and (_20361_, _20360_, _27053_);
  and (_28966_, _20361_, _20358_);
  and (_20362_, _03121_, _02259_);
  and (_20363_, _02256_, _01900_);
  and (_20364_, _20363_, \oc8051_golden_model_1.PC [7]);
  nor (_20365_, _20363_, \oc8051_golden_model_1.PC [7]);
  nor (_20366_, _20365_, _20364_);
  nor (_20367_, _20366_, _01930_);
  nor (_20368_, _20366_, _05389_);
  not (_20370_, _20366_);
  and (_20371_, _20370_, _01944_);
  and (_20372_, _20370_, _05325_);
  and (_20373_, _20370_, _05297_);
  and (_20374_, _02577_, _02260_);
  and (_20375_, _03140_, _02260_);
  and (_20376_, _20370_, _05194_);
  nor (_20377_, _05177_, _02259_);
  and (_20378_, _20370_, _02598_);
  and (_20379_, _04494_, _02800_);
  or (_20381_, _02802_, _02803_);
  not (_20382_, _20381_);
  nor (_20383_, _20382_, _03069_);
  and (_20384_, _20382_, _03069_);
  nor (_20385_, _20384_, _20383_);
  nor (_20386_, _20385_, _04494_);
  or (_20387_, _20386_, _20379_);
  nor (_20388_, _20387_, _04499_);
  and (_20389_, _20385_, _04987_);
  and (_20390_, _04985_, _02801_);
  nor (_20392_, _20390_, _20389_);
  or (_20393_, _20392_, _02662_);
  and (_20394_, _04540_, _02259_);
  and (_20395_, _02524_, _02264_);
  nor (_20396_, _20395_, _02525_);
  and (_20397_, _20396_, _04537_);
  or (_20398_, _20397_, _20394_);
  nor (_20399_, _20398_, _04539_);
  and (_20400_, _20370_, _04510_);
  nor (_20401_, _02752_, _01988_);
  and (_20403_, _04505_, _02260_);
  nor (_20404_, _20403_, _04520_);
  and (_20405_, _19685_, \oc8051_golden_model_1.PC [7]);
  or (_20406_, _20405_, _04505_);
  and (_20407_, _20406_, _20404_);
  nor (_20408_, _20370_, _04521_);
  or (_20409_, _20408_, _04510_);
  or (_20410_, _20409_, _20407_);
  and (_20411_, _20410_, _01988_);
  nor (_20412_, _20411_, _20401_);
  or (_20414_, _20412_, _03154_);
  nor (_20415_, _20414_, _20400_);
  and (_20416_, _03154_, _02259_);
  or (_20417_, _20416_, _20415_);
  and (_20418_, _20417_, _18144_);
  and (_20419_, _20366_, _04502_);
  or (_20420_, _20419_, _20418_);
  and (_20421_, _20420_, _01998_);
  nor (_20422_, _02752_, _01998_);
  nor (_20423_, _20422_, _03406_);
  not (_20425_, _20423_);
  nor (_20426_, _20425_, _20421_);
  or (_20427_, _20426_, _04545_);
  nor (_20428_, _20427_, _20399_);
  and (_20429_, _20366_, _04545_);
  or (_20430_, _20429_, _02661_);
  or (_20431_, _20430_, _20428_);
  and (_20432_, _20431_, _20393_);
  nor (_20433_, _20432_, _04992_);
  and (_20434_, _20370_, _04992_);
  nor (_20436_, _20434_, _03150_);
  not (_20437_, _20436_);
  or (_20438_, _20437_, _20433_);
  and (_20439_, _03150_, _02259_);
  nor (_20440_, _20439_, _07558_);
  nand (_20441_, _20440_, _20438_);
  and (_20442_, _02752_, _07558_);
  nor (_20443_, _20442_, _03162_);
  nand (_20444_, _20443_, _20441_);
  and (_20445_, _03162_, _02259_);
  nor (_20447_, _20445_, _05000_);
  nand (_20448_, _20447_, _20444_);
  and (_20449_, _20370_, _05000_);
  nor (_20450_, _20449_, _03168_);
  nand (_20451_, _20450_, _20448_);
  and (_20452_, _03168_, _02259_);
  nor (_20453_, _20452_, _05009_);
  nand (_20454_, _20453_, _20451_);
  and (_20455_, _20370_, _05009_);
  nor (_20456_, _20455_, _03176_);
  nand (_20458_, _20456_, _20454_);
  and (_20459_, _03176_, _02259_);
  nor (_20460_, _20459_, _17919_);
  nand (_20461_, _20460_, _20458_);
  and (_20462_, _02752_, _17919_);
  nor (_20463_, _20462_, _03187_);
  nand (_20464_, _20463_, _20461_);
  and (_20465_, _03187_, _02259_);
  nor (_20466_, _20465_, _04498_);
  and (_20467_, _20466_, _20464_);
  nor (_20469_, _20467_, _20388_);
  or (_20470_, _20469_, _02675_);
  not (_20471_, _20385_);
  and (_20472_, _20471_, _04277_);
  and (_20473_, _04275_, _02800_);
  or (_20474_, _20473_, _03107_);
  or (_20475_, _20474_, _20472_);
  nand (_20476_, _20475_, _20470_);
  or (_20477_, _20476_, _02664_);
  nor (_20478_, _20385_, _05157_);
  and (_20480_, _05157_, _02800_);
  nor (_20481_, _20480_, _20478_);
  or (_20482_, _20481_, _03387_);
  and (_20483_, _20482_, _20477_);
  or (_20484_, _20483_, _02673_);
  and (_20485_, _02800_, _02630_);
  nor (_20486_, _20385_, _02630_);
  or (_20487_, _20486_, _20485_);
  and (_20488_, _20487_, _02673_);
  nor (_20489_, _20488_, _02598_);
  and (_20491_, _20489_, _20484_);
  or (_20492_, _20491_, _20378_);
  nand (_20493_, _20492_, _05168_);
  and (_20494_, _03144_, _02260_);
  nor (_20495_, _20494_, _06664_);
  nand (_20496_, _20495_, _20493_);
  nor (_20497_, _02752_, _02000_);
  nor (_20498_, _20497_, _18254_);
  and (_20499_, _20498_, _20496_);
  or (_20500_, _20499_, _20377_);
  nand (_20502_, _20500_, _05186_);
  and (_20503_, _20370_, _05185_);
  nor (_20504_, _20503_, _03205_);
  nand (_20505_, _20504_, _20502_);
  and (_20506_, _03205_, _02259_);
  nor (_20507_, _20506_, _17956_);
  nand (_20508_, _20507_, _20505_);
  and (_20509_, _02752_, _17956_);
  nor (_20510_, _20509_, _03203_);
  nand (_20511_, _20510_, _20508_);
  and (_20513_, _03203_, _02259_);
  nor (_20514_, _20513_, _05194_);
  and (_20515_, _20514_, _20511_);
  or (_20516_, _20515_, _20376_);
  nand (_20517_, _20516_, _05203_);
  and (_20518_, _05199_, _02260_);
  nor (_20519_, _20518_, _02047_);
  nand (_20520_, _20519_, _20517_);
  nor (_20521_, _20370_, _01985_);
  nor (_20522_, _20521_, _03140_);
  and (_20524_, _20522_, _20520_);
  or (_20525_, _20524_, _20375_);
  nand (_20526_, _20525_, _07791_);
  and (_20527_, _02752_, _02025_);
  nor (_20528_, _20527_, _02670_);
  nand (_20529_, _20528_, _20526_);
  and (_20530_, _02800_, _02670_);
  nor (_20531_, _20530_, _05217_);
  nand (_20532_, _20531_, _20529_);
  and (_20533_, _05217_, _02260_);
  nor (_20535_, _20533_, _02024_);
  nand (_20536_, _20535_, _20532_);
  and (_20537_, _02800_, _02024_);
  nor (_20538_, _20537_, _05225_);
  nand (_20539_, _20538_, _20536_);
  and (_20540_, _20370_, _05225_);
  nor (_20541_, _20540_, _03135_);
  nand (_20542_, _20541_, _20539_);
  and (_20543_, _03135_, _02259_);
  nor (_20544_, _20543_, _01960_);
  nand (_20546_, _20544_, _20542_);
  and (_20547_, _02752_, _01960_);
  nor (_20548_, _20547_, _05233_);
  nand (_20549_, _20548_, _20546_);
  and (_20550_, _20396_, _05233_);
  nor (_20551_, _20550_, _02577_);
  and (_20552_, _20551_, _20549_);
  or (_20553_, _20552_, _20374_);
  nand (_20554_, _20553_, _05245_);
  and (_20555_, _02801_, _02575_);
  nor (_20557_, _20555_, _05243_);
  and (_20558_, _20557_, _20554_);
  and (_20559_, _05243_, _02259_);
  or (_20560_, _20559_, _20558_);
  nand (_20561_, _20560_, _02574_);
  or (_20562_, _05256_, _05255_);
  nor (_20563_, _20562_, _05275_);
  and (_20564_, _20562_, _05275_);
  or (_20565_, _20564_, _02574_);
  or (_20566_, _20565_, _20563_);
  and (_20568_, _20566_, _18752_);
  and (_20569_, _20568_, _20561_);
  and (_20570_, _03134_, _02260_);
  or (_20571_, _20570_, _20569_);
  nand (_20572_, _20571_, _13603_);
  and (_20573_, _02752_, _01967_);
  nor (_20574_, _20573_, _02567_);
  nand (_20575_, _20574_, _20572_);
  and (_20576_, _02259_, _01953_);
  and (_20577_, _20396_, _02568_);
  or (_20579_, _20577_, _20576_);
  and (_20580_, _20579_, _02567_);
  nor (_20581_, _20580_, _05297_);
  and (_20582_, _20581_, _20575_);
  or (_20583_, _20582_, _20373_);
  nand (_20584_, _20583_, _05306_);
  and (_20585_, _05302_, _02260_);
  nor (_20586_, _20585_, _02656_);
  nand (_20587_, _20586_, _20584_);
  and (_20588_, _02800_, _02656_);
  nor (_20590_, _20588_, _03251_);
  and (_20591_, _20590_, _20587_);
  and (_20592_, _03251_, _02260_);
  or (_20593_, _20592_, _20591_);
  nand (_20594_, _20593_, _17855_);
  and (_20595_, _02752_, _01974_);
  nor (_20596_, _20595_, _05315_);
  nand (_20597_, _20596_, _20594_);
  and (_20598_, _02259_, _02568_);
  and (_20599_, _20396_, _01953_);
  or (_20601_, _20599_, _20598_);
  and (_20602_, _20601_, _05315_);
  nor (_20603_, _20602_, _05325_);
  and (_20604_, _20603_, _20597_);
  or (_20605_, _20604_, _20372_);
  nand (_20606_, _20605_, _05333_);
  and (_20607_, _05329_, _02260_);
  nor (_20608_, _20607_, _02669_);
  nand (_20609_, _20608_, _20606_);
  and (_20610_, _02800_, _02669_);
  nor (_20612_, _20610_, _03243_);
  and (_20613_, _20612_, _20609_);
  and (_20614_, _03243_, _02260_);
  or (_20615_, _20614_, _20613_);
  nand (_20616_, _20615_, _17852_);
  and (_20617_, _02752_, _01965_);
  nor (_20618_, _20617_, _05342_);
  nand (_20619_, _20618_, _20616_);
  nor (_20620_, _20396_, \oc8051_golden_model_1.PSW [7]);
  nor (_20621_, _02259_, _05348_);
  nor (_20623_, _20621_, _05343_);
  not (_20624_, _20623_);
  nor (_20625_, _20624_, _20620_);
  nor (_20626_, _20625_, _01944_);
  and (_20627_, _20626_, _20619_);
  or (_20628_, _20627_, _20371_);
  nand (_20629_, _20628_, _05358_);
  and (_20630_, _05355_, _02260_);
  nor (_20631_, _20630_, _02654_);
  nand (_20632_, _20631_, _20629_);
  and (_20634_, _02800_, _02654_);
  nor (_20635_, _20634_, _03239_);
  and (_20636_, _20635_, _20632_);
  and (_20637_, _03239_, _02260_);
  or (_20638_, _20637_, _20636_);
  nand (_20639_, _20638_, _17848_);
  and (_20640_, _02752_, _01957_);
  nor (_20641_, _20640_, _05367_);
  nand (_20642_, _20641_, _20639_);
  and (_20643_, _02259_, _05348_);
  and (_20645_, _20396_, \oc8051_golden_model_1.PSW [7]);
  or (_20646_, _20645_, _20643_);
  and (_20647_, _20646_, _05367_);
  nor (_20648_, _20647_, _05391_);
  and (_20649_, _20648_, _20642_);
  or (_20650_, _20649_, _20368_);
  nand (_20651_, _20650_, _05398_);
  and (_20652_, _05393_, _02260_);
  nor (_20653_, _20652_, _05396_);
  nand (_20654_, _20653_, _20651_);
  and (_20656_, _20366_, _05396_);
  nor (_20657_, _20656_, _03109_);
  and (_20658_, _20657_, _20654_);
  and (_20659_, _04069_, _03109_);
  or (_20660_, _20659_, _20658_);
  nand (_20661_, _20660_, _05408_);
  and (_20662_, _02752_, _01936_);
  nor (_20663_, _20662_, _02653_);
  nand (_20664_, _20663_, _20661_);
  and (_20665_, _20385_, _05702_);
  nor (_20667_, _05702_, _02800_);
  or (_20668_, _20667_, _03267_);
  or (_20669_, _20668_, _20665_);
  and (_20670_, _20669_, _01930_);
  and (_20671_, _20670_, _20664_);
  or (_20672_, _20671_, _20367_);
  nand (_20673_, _20672_, _05728_);
  and (_20674_, _05720_, _02260_);
  nor (_20675_, _20674_, _05724_);
  nand (_20676_, _20675_, _20673_);
  and (_20678_, _20366_, _05724_);
  nor (_20679_, _20678_, _03108_);
  and (_20680_, _20679_, _20676_);
  and (_20681_, _04069_, _03108_);
  or (_20682_, _20681_, _20680_);
  nand (_20683_, _20682_, _05748_);
  and (_20684_, _02752_, _01899_);
  nor (_20685_, _20684_, _02647_);
  nand (_20686_, _20685_, _20683_);
  and (_20687_, _05702_, _02801_);
  nor (_20689_, _20471_, _05702_);
  nor (_20690_, _20689_, _20687_);
  and (_20691_, _20690_, _02647_);
  nor (_20692_, _20691_, _05764_);
  nand (_20693_, _20692_, _20686_);
  and (_20694_, _20370_, _05764_);
  nor (_20695_, _20694_, _03123_);
  nand (_20696_, _20695_, _20693_);
  and (_20697_, _03123_, _02259_);
  nor (_20698_, _20697_, _05780_);
  and (_20700_, _20698_, _20696_);
  and (_20701_, _20370_, _05780_);
  or (_20702_, _20701_, _20700_);
  nand (_20703_, _20702_, _06741_);
  and (_20704_, _06742_, _02752_);
  nor (_20705_, _20704_, _02650_);
  nand (_20706_, _20705_, _20703_);
  and (_20707_, _20690_, _02650_);
  nor (_20708_, _20707_, _05826_);
  nand (_20709_, _20708_, _20706_);
  nor (_20711_, _20366_, _05824_);
  nor (_20712_, _20711_, _03121_);
  and (_20713_, _20712_, _20709_);
  or (_20714_, _20713_, _20362_);
  nand (_20715_, _20714_, _05848_);
  and (_20716_, _20366_, _05840_);
  nor (_20717_, _20716_, _18101_);
  nand (_20718_, _20717_, _20715_);
  and (_20719_, _18101_, _02752_);
  nor (_20720_, _20719_, _05862_);
  nand (_20722_, _20720_, _20718_);
  and (_20723_, _20366_, _05862_);
  not (_20724_, _20723_);
  and (_20725_, _20724_, _20722_);
  nand (_20726_, _20725_, _27788_);
  or (_20727_, _27788_, \oc8051_golden_model_1.PC [7]);
  and (_20728_, _20727_, _27053_);
  and (_28967_, _20728_, _20726_);
  nor (_20729_, _05846_, _02503_);
  nor (_20730_, _05786_, _02503_);
  nor (_20732_, _20364_, \oc8051_golden_model_1.PC [8]);
  and (_20733_, _20364_, \oc8051_golden_model_1.PC [8]);
  nor (_20734_, _20733_, _20732_);
  nor (_20735_, _20734_, _01930_);
  nor (_20736_, _20734_, _05389_);
  not (_20737_, _20734_);
  and (_20738_, _20737_, _01944_);
  and (_20739_, _20737_, _05325_);
  and (_20740_, _03073_, _02656_);
  and (_20741_, _20737_, _05297_);
  and (_20743_, _02577_, _02529_);
  and (_20744_, _20737_, _05225_);
  and (_20745_, _20737_, _05194_);
  nor (_20746_, _05177_, _02528_);
  nor (_20747_, _03187_, _17919_);
  and (_20748_, _03176_, _02528_);
  and (_20749_, _03162_, _02528_);
  and (_20750_, _03150_, _02528_);
  or (_20751_, _20734_, _04522_);
  and (_20752_, _04505_, _02528_);
  and (_20754_, _05903_, \oc8051_golden_model_1.PC [8]);
  and (_20755_, _20754_, _04521_);
  or (_20756_, _20755_, _18582_);
  and (_20757_, _20756_, _04503_);
  or (_20758_, _20757_, _20752_);
  and (_20759_, _20758_, _20751_);
  nand (_20760_, _04521_, _18144_);
  and (_20761_, _20760_, _20734_);
  nor (_20762_, _03406_, _04527_);
  not (_20763_, _20762_);
  and (_20765_, _03154_, _02528_);
  or (_20766_, _20765_, _20763_);
  or (_20767_, _20766_, _20761_);
  nor (_20768_, _20767_, _20759_);
  and (_20769_, _04540_, _02528_);
  and (_20770_, _02533_, _02526_);
  nor (_20771_, _20770_, _02534_);
  and (_20772_, _20771_, _04537_);
  or (_20773_, _20772_, _20769_);
  nor (_20774_, _20773_, _04539_);
  nor (_20776_, _20774_, _20768_);
  nor (_20777_, _20776_, _04545_);
  and (_20778_, _20737_, _04545_);
  or (_20779_, _20778_, _02661_);
  nor (_20780_, _20779_, _20777_);
  nor (_20781_, _03077_, _03071_);
  nor (_20782_, _20781_, _03078_);
  not (_20783_, _20782_);
  and (_20784_, _20783_, _04987_);
  and (_20785_, _04985_, _03074_);
  or (_20787_, _20785_, _02662_);
  nor (_20788_, _20787_, _20784_);
  or (_20789_, _20788_, _04992_);
  nor (_20790_, _20789_, _20780_);
  and (_20791_, _20737_, _04992_);
  nor (_20792_, _20791_, _03150_);
  not (_20793_, _20792_);
  nor (_20794_, _20793_, _20790_);
  nor (_20795_, _20794_, _20750_);
  nor (_20796_, _20795_, _07558_);
  and (_20798_, _20796_, _03365_);
  or (_20799_, _20798_, _05000_);
  nor (_20800_, _20799_, _20749_);
  and (_20801_, _20737_, _05000_);
  nor (_20802_, _20801_, _03168_);
  not (_20803_, _20802_);
  nor (_20804_, _20803_, _20800_);
  and (_20805_, _03168_, _02528_);
  nor (_20806_, _20805_, _05009_);
  not (_20807_, _20806_);
  nor (_20809_, _20807_, _20804_);
  and (_20810_, _20737_, _05009_);
  nor (_20811_, _20810_, _03176_);
  not (_20812_, _20811_);
  nor (_20813_, _20812_, _20809_);
  or (_20814_, _20813_, _20748_);
  nand (_20815_, _20814_, _20747_);
  and (_20816_, _03187_, _02528_);
  nor (_20817_, _20816_, _04498_);
  and (_20818_, _20817_, _20815_);
  nor (_20820_, _20783_, _04494_);
  not (_20821_, _20820_);
  and (_20822_, _04494_, _03073_);
  nor (_20823_, _20822_, _04499_);
  and (_20824_, _20823_, _20821_);
  nor (_20825_, _20824_, _20818_);
  or (_20826_, _20825_, _02675_);
  and (_20827_, _04275_, _03073_);
  and (_20828_, _20782_, _04277_);
  or (_20829_, _20828_, _03107_);
  or (_20831_, _20829_, _20827_);
  nand (_20832_, _20831_, _20826_);
  or (_20833_, _20832_, _02664_);
  and (_20834_, _05157_, _03073_);
  nor (_20835_, _20783_, _05157_);
  nor (_20836_, _20835_, _20834_);
  or (_20837_, _20836_, _03387_);
  and (_20838_, _20837_, _20833_);
  or (_20839_, _20838_, _02673_);
  and (_20840_, _03073_, _02630_);
  and (_20842_, _20782_, _19401_);
  or (_20843_, _20842_, _20840_);
  and (_20844_, _20843_, _02673_);
  nor (_20845_, _20844_, _02598_);
  nand (_20846_, _20845_, _20839_);
  and (_20847_, _20737_, _02598_);
  nor (_20848_, _20847_, _03144_);
  nand (_20849_, _20848_, _20846_);
  and (_20850_, _03144_, _02528_);
  not (_20851_, _20850_);
  and (_20853_, _20851_, _05178_);
  and (_20854_, _20853_, _20849_);
  or (_20855_, _20854_, _20746_);
  nand (_20856_, _20855_, _05186_);
  and (_20857_, _20737_, _05185_);
  nor (_20858_, _20857_, _03205_);
  nand (_20859_, _20858_, _20856_);
  and (_20860_, _03205_, _02528_);
  nor (_20861_, _20860_, _17956_);
  nand (_20862_, _20861_, _20859_);
  nand (_20864_, _20862_, _18677_);
  and (_20865_, _03203_, _02528_);
  nor (_20866_, _20865_, _05194_);
  and (_20867_, _20866_, _20864_);
  or (_20868_, _20867_, _20745_);
  nand (_20869_, _20868_, _05203_);
  and (_20870_, _05199_, _02529_);
  nor (_20871_, _20870_, _02047_);
  nand (_20872_, _20871_, _20869_);
  nor (_20873_, _20737_, _01985_);
  nor (_20875_, _20873_, _03140_);
  nand (_20876_, _20875_, _20872_);
  nor (_20877_, _02670_, _02025_);
  not (_20878_, _20877_);
  and (_20879_, _03140_, _02529_);
  nor (_20880_, _20879_, _20878_);
  nand (_20881_, _20880_, _20876_);
  and (_20882_, _03073_, _02670_);
  nor (_20883_, _20882_, _05217_);
  nand (_20884_, _20883_, _20881_);
  and (_20886_, _05217_, _02529_);
  nor (_20887_, _20886_, _02024_);
  nand (_20888_, _20887_, _20884_);
  and (_20889_, _03073_, _02024_);
  nor (_20890_, _20889_, _05225_);
  and (_20891_, _20890_, _20888_);
  nor (_20892_, _20891_, _20744_);
  or (_20893_, _20892_, _03135_);
  nor (_20894_, _05233_, _01960_);
  nand (_20895_, _03135_, _02529_);
  and (_20897_, _20895_, _20894_);
  nand (_20898_, _20897_, _20893_);
  and (_20899_, _20771_, _05233_);
  nor (_20900_, _20899_, _02577_);
  and (_20901_, _20900_, _20898_);
  or (_20902_, _20901_, _20743_);
  nand (_20903_, _20902_, _05245_);
  and (_20904_, _03074_, _02575_);
  nor (_20905_, _20904_, _05243_);
  nand (_20906_, _20905_, _20903_);
  and (_20908_, _05243_, _02528_);
  nor (_20909_, _20908_, _02573_);
  nand (_20910_, _20909_, _20906_);
  and (_20911_, _05277_, _05254_);
  nor (_20912_, _20911_, _05278_);
  nor (_20913_, _20912_, _02574_);
  nor (_20914_, _20913_, _03134_);
  nand (_20915_, _20914_, _20910_);
  and (_20916_, _03134_, _02528_);
  nor (_20917_, _20916_, _01967_);
  nand (_20919_, _20917_, _20915_);
  nand (_20920_, _20919_, _05291_);
  and (_20921_, _02528_, _01953_);
  and (_20922_, _20771_, _02568_);
  or (_20923_, _20922_, _20921_);
  and (_20924_, _20923_, _02567_);
  nor (_20925_, _20924_, _05297_);
  and (_20926_, _20925_, _20920_);
  or (_20927_, _20926_, _20741_);
  nand (_20928_, _20927_, _05306_);
  and (_20930_, _05302_, _02529_);
  nor (_20931_, _20930_, _02656_);
  and (_20932_, _20931_, _20928_);
  or (_20933_, _20932_, _20740_);
  nand (_20934_, _20933_, _03252_);
  and (_20935_, _03251_, _02528_);
  nor (_20936_, _20935_, _01974_);
  nand (_20937_, _20936_, _20934_);
  nand (_20938_, _20937_, _05316_);
  and (_20939_, _02528_, _02568_);
  and (_20941_, _20771_, _01953_);
  or (_20942_, _20941_, _20939_);
  and (_20943_, _20942_, _05315_);
  nor (_20944_, _20943_, _05325_);
  and (_20945_, _20944_, _20938_);
  or (_20946_, _20945_, _20739_);
  nand (_20947_, _20946_, _05333_);
  and (_20948_, _05329_, _02529_);
  nor (_20949_, _20948_, _02669_);
  nand (_20950_, _20949_, _20947_);
  and (_20952_, _03073_, _02669_);
  nor (_20953_, _20952_, _03243_);
  nand (_20954_, _20953_, _20950_);
  and (_20955_, _03243_, _02529_);
  nor (_20956_, _05342_, _01965_);
  not (_20957_, _20956_);
  nor (_20958_, _20957_, _20955_);
  nand (_20959_, _20958_, _20954_);
  nor (_20960_, _20771_, \oc8051_golden_model_1.PSW [7]);
  nor (_20961_, _02528_, _05348_);
  nor (_20963_, _20961_, _05343_);
  not (_20964_, _20963_);
  nor (_20965_, _20964_, _20960_);
  nor (_20966_, _20965_, _01944_);
  and (_20967_, _20966_, _20959_);
  or (_20968_, _20967_, _20738_);
  nand (_20969_, _20968_, _05358_);
  and (_20970_, _05355_, _02529_);
  nor (_20971_, _20970_, _02654_);
  and (_20972_, _20971_, _20969_);
  and (_20974_, _03073_, _02654_);
  or (_20975_, _20974_, _03239_);
  or (_20976_, _20975_, _20972_);
  and (_20977_, _03239_, _02529_);
  nor (_20978_, _05367_, _01957_);
  not (_20979_, _20978_);
  nor (_20980_, _20979_, _20977_);
  nand (_20981_, _20980_, _20976_);
  and (_20982_, _02528_, _05348_);
  and (_20983_, _20771_, \oc8051_golden_model_1.PSW [7]);
  or (_20985_, _20983_, _20982_);
  and (_20986_, _20985_, _05367_);
  nor (_20987_, _20986_, _05391_);
  and (_20988_, _20987_, _20981_);
  or (_20989_, _20988_, _20736_);
  nand (_20990_, _20989_, _05398_);
  and (_20991_, _05393_, _02529_);
  nor (_20992_, _20991_, _05396_);
  and (_20993_, _20992_, _20990_);
  and (_20994_, _20734_, _05396_);
  or (_20996_, _20994_, _20993_);
  nand (_20997_, _20996_, _06612_);
  and (_20998_, _03716_, _03109_);
  nor (_20999_, _20998_, _01936_);
  nand (_21000_, _20999_, _20997_);
  nand (_21001_, _21000_, _03267_);
  nor (_21002_, _05702_, _03073_);
  and (_21003_, _20783_, _05702_);
  or (_21004_, _21003_, _03267_);
  nor (_21005_, _21004_, _21002_);
  nor (_21007_, _21005_, _05412_);
  and (_21008_, _21007_, _21001_);
  or (_21009_, _21008_, _20735_);
  nand (_21010_, _21009_, _05728_);
  and (_21011_, _05720_, _02529_);
  nor (_21012_, _21011_, _05724_);
  and (_21013_, _21012_, _21010_);
  and (_21014_, _20734_, _05724_);
  or (_21015_, _21014_, _21013_);
  nand (_21016_, _21015_, _03126_);
  and (_21018_, _03716_, _03108_);
  nor (_21019_, _21018_, _01899_);
  nand (_21020_, _21019_, _21016_);
  nand (_21021_, _21020_, _03125_);
  and (_21022_, _05702_, _03074_);
  nor (_21023_, _20782_, _05702_);
  nor (_21024_, _21023_, _21022_);
  and (_21025_, _21024_, _02647_);
  nor (_21026_, _21025_, _05764_);
  nand (_21027_, _21026_, _21021_);
  and (_21029_, _20737_, _05764_);
  nor (_21030_, _21029_, _03123_);
  nand (_21031_, _21030_, _21027_);
  and (_21032_, _03123_, _02528_);
  nor (_21033_, _21032_, _05780_);
  nand (_21034_, _21033_, _21031_);
  and (_21035_, _20737_, _05780_);
  nor (_21036_, _21035_, _02646_);
  and (_21037_, _21036_, _21034_);
  or (_21038_, _21037_, _20730_);
  nor (_21040_, _02650_, _01971_);
  nand (_21041_, _21040_, _21038_);
  and (_21042_, _21024_, _02650_);
  nor (_21043_, _21042_, _05826_);
  nand (_21044_, _21043_, _21041_);
  nor (_21045_, _20734_, _05824_);
  nor (_21046_, _21045_, _03121_);
  nand (_21047_, _21046_, _21044_);
  and (_21048_, _03121_, _02528_);
  nor (_21049_, _21048_, _05840_);
  nand (_21051_, _21049_, _21047_);
  and (_21052_, _20737_, _05840_);
  nor (_21053_, _21052_, _02649_);
  and (_21054_, _21053_, _21051_);
  or (_21055_, _21054_, _20729_);
  nor (_21056_, _05862_, _01955_);
  and (_21057_, _21056_, _21055_);
  and (_21058_, _20734_, _05862_);
  or (_21059_, _21058_, _21057_);
  or (_21060_, _21059_, _27789_);
  or (_21062_, _27788_, \oc8051_golden_model_1.PC [8]);
  and (_21063_, _21062_, _27053_);
  and (_28968_, _21063_, _21060_);
  nor (_21064_, _05786_, _02471_);
  not (_21065_, \oc8051_golden_model_1.PC [9]);
  and (_21066_, _02208_, _01900_);
  and (_21067_, _21066_, \oc8051_golden_model_1.PC [8]);
  nor (_21068_, _21067_, _21065_);
  and (_21069_, _21067_, _21065_);
  or (_21070_, _21069_, _21068_);
  nor (_21072_, _21070_, _01930_);
  nor (_21073_, _21070_, _05389_);
  and (_21074_, _02793_, _02654_);
  not (_21075_, _21070_);
  and (_21076_, _21075_, _01944_);
  and (_21077_, _02793_, _02669_);
  and (_21078_, _21075_, _05325_);
  and (_21079_, _02793_, _02656_);
  and (_21080_, _21075_, _05297_);
  and (_21081_, _02577_, _02252_);
  and (_21083_, _03135_, _02251_);
  and (_21084_, _03203_, _02251_);
  nor (_21085_, _03203_, _17956_);
  and (_21086_, _21075_, _02598_);
  and (_21087_, _03162_, _02251_);
  nor (_21088_, _03078_, _03075_);
  and (_21089_, _21088_, _02797_);
  nor (_21090_, _21088_, _02797_);
  nor (_21091_, _21090_, _21089_);
  not (_21092_, _21091_);
  and (_21094_, _21092_, _04987_);
  and (_21095_, _04985_, _02793_);
  or (_21096_, _21095_, _02662_);
  or (_21097_, _21096_, _21094_);
  and (_21098_, _04540_, _02251_);
  nor (_21099_, _02534_, _02530_);
  and (_21100_, _21099_, _02255_);
  nor (_21101_, _21099_, _02255_);
  nor (_21102_, _21101_, _21100_);
  nor (_21103_, _21102_, _04540_);
  or (_21105_, _21103_, _21098_);
  nor (_21106_, _21105_, _04539_);
  and (_21107_, _04505_, _02251_);
  nor (_21108_, _04505_, _21065_);
  and (_21109_, _21108_, _04521_);
  or (_21110_, _21109_, _18582_);
  and (_21111_, _21110_, _04503_);
  or (_21112_, _21111_, _21107_);
  or (_21113_, _21070_, _04522_);
  and (_21114_, _21113_, _21112_);
  and (_21116_, _21070_, _20760_);
  and (_21117_, _03154_, _02251_);
  or (_21118_, _21117_, _20763_);
  or (_21119_, _21118_, _21116_);
  nor (_21120_, _21119_, _21114_);
  or (_21121_, _21120_, _04545_);
  nor (_21122_, _21121_, _21106_);
  and (_21123_, _21070_, _04545_);
  or (_21124_, _21123_, _02661_);
  or (_21125_, _21124_, _21122_);
  and (_21127_, _21125_, _21097_);
  nor (_21128_, _21127_, _04992_);
  and (_21129_, _21075_, _04992_);
  nor (_21130_, _21129_, _03150_);
  not (_21131_, _21130_);
  nor (_21132_, _21131_, _21128_);
  and (_21133_, _03150_, _02251_);
  or (_21134_, _21133_, _07558_);
  nor (_21135_, _21134_, _21132_);
  nor (_21136_, _21135_, _03162_);
  or (_21138_, _21136_, _05000_);
  nor (_21139_, _21138_, _21087_);
  and (_21140_, _21075_, _05000_);
  nor (_21141_, _21140_, _03168_);
  not (_21142_, _21141_);
  or (_21143_, _21142_, _21139_);
  and (_21144_, _03168_, _02251_);
  nor (_21145_, _21144_, _05009_);
  nand (_21146_, _21145_, _21143_);
  and (_21147_, _21075_, _05009_);
  nor (_21149_, _21147_, _03176_);
  nand (_21150_, _21149_, _21146_);
  and (_21151_, _03176_, _02251_);
  nor (_21152_, _21151_, _17919_);
  nand (_21153_, _21152_, _21150_);
  nand (_21154_, _21153_, _03430_);
  and (_21155_, _03187_, _02251_);
  nor (_21156_, _21155_, _04498_);
  and (_21157_, _21156_, _21154_);
  and (_21158_, _04494_, _02793_);
  nor (_21160_, _21091_, _04494_);
  or (_21161_, _21160_, _04499_);
  nor (_21162_, _21161_, _21158_);
  nor (_21163_, _21162_, _21157_);
  or (_21164_, _21163_, _02675_);
  and (_21165_, _04275_, _02793_);
  and (_21166_, _21092_, _04277_);
  or (_21167_, _21166_, _03107_);
  or (_21168_, _21167_, _21165_);
  nand (_21169_, _21168_, _21164_);
  or (_21171_, _21169_, _02664_);
  and (_21172_, _05157_, _02793_);
  nor (_21173_, _21091_, _05157_);
  nor (_21174_, _21173_, _21172_);
  or (_21175_, _21174_, _03387_);
  and (_21176_, _21175_, _21171_);
  or (_21177_, _21176_, _02673_);
  and (_21178_, _02793_, _02630_);
  nor (_21179_, _21091_, _02630_);
  or (_21180_, _21179_, _21178_);
  and (_21182_, _21180_, _02673_);
  nor (_21183_, _21182_, _02598_);
  and (_21184_, _21183_, _21177_);
  or (_21185_, _21184_, _21086_);
  and (_21186_, _21185_, _05168_);
  and (_21187_, _05178_, _02251_);
  nor (_21188_, _21187_, _05179_);
  or (_21189_, _21188_, _21186_);
  nor (_21190_, _05177_, _02252_);
  nor (_21191_, _21190_, _05185_);
  nand (_21193_, _21191_, _21189_);
  and (_21194_, _21075_, _05185_);
  nor (_21195_, _21194_, _03205_);
  and (_21196_, _21195_, _21193_);
  and (_21197_, _03205_, _02251_);
  or (_21198_, _21197_, _21196_);
  and (_21199_, _21198_, _21085_);
  or (_21200_, _21199_, _21084_);
  nand (_21201_, _21200_, _05195_);
  and (_21202_, _21070_, _05194_);
  nor (_21204_, _21202_, _05199_);
  nand (_21205_, _21204_, _21201_);
  and (_21206_, _05199_, _02252_);
  nor (_21207_, _21206_, _02047_);
  nand (_21208_, _21207_, _21205_);
  nor (_21209_, _21075_, _01985_);
  nor (_21210_, _21209_, _03140_);
  nand (_21211_, _21210_, _21208_);
  and (_21212_, _03140_, _02252_);
  nor (_21213_, _21212_, _20878_);
  nand (_21215_, _21213_, _21211_);
  and (_21216_, _02793_, _02670_);
  nor (_21217_, _21216_, _05217_);
  nand (_21218_, _21217_, _21215_);
  and (_21219_, _05217_, _02252_);
  nor (_21220_, _21219_, _02024_);
  nand (_21221_, _21220_, _21218_);
  and (_21222_, _02793_, _02024_);
  nor (_21223_, _21222_, _05225_);
  nand (_21224_, _21223_, _21221_);
  and (_21226_, _21075_, _05225_);
  nor (_21227_, _21226_, _03135_);
  and (_21228_, _21227_, _21224_);
  or (_21229_, _21228_, _21083_);
  nand (_21230_, _21229_, _20894_);
  nor (_21231_, _21102_, _05234_);
  nor (_21232_, _21231_, _02577_);
  and (_21233_, _21232_, _21230_);
  or (_21234_, _21233_, _21081_);
  nand (_21235_, _21234_, _05245_);
  and (_21237_, _02794_, _02575_);
  nor (_21238_, _21237_, _05243_);
  nand (_21239_, _21238_, _21235_);
  and (_21240_, _05243_, _02251_);
  nor (_21241_, _21240_, _02573_);
  nand (_21242_, _21241_, _21239_);
  nor (_21243_, _05278_, \oc8051_golden_model_1.DPH [1]);
  nor (_21244_, _21243_, _05279_);
  nor (_21245_, _21244_, _02574_);
  nor (_21246_, _21245_, _03134_);
  nand (_21248_, _21246_, _21242_);
  and (_21249_, _03134_, _02251_);
  nor (_21250_, _21249_, _01967_);
  nand (_21251_, _21250_, _21248_);
  nand (_21252_, _21251_, _05291_);
  and (_21253_, _21102_, _02568_);
  nor (_21254_, _02251_, _02568_);
  nor (_21255_, _21254_, _05291_);
  not (_21256_, _21255_);
  nor (_21257_, _21256_, _21253_);
  nor (_21259_, _21257_, _05297_);
  and (_21260_, _21259_, _21252_);
  or (_21261_, _21260_, _21080_);
  nand (_21262_, _21261_, _05306_);
  and (_21263_, _05302_, _02252_);
  nor (_21264_, _21263_, _02656_);
  and (_21265_, _21264_, _21262_);
  or (_21266_, _21265_, _21079_);
  nand (_21267_, _21266_, _03252_);
  and (_21268_, _03251_, _02251_);
  nor (_21270_, _21268_, _01974_);
  nand (_21271_, _21270_, _21267_);
  nand (_21272_, _21271_, _05316_);
  and (_21273_, _02251_, _02568_);
  nor (_21274_, _21102_, _02568_);
  or (_21275_, _21274_, _21273_);
  and (_21276_, _21275_, _05315_);
  nor (_21277_, _21276_, _05325_);
  and (_21278_, _21277_, _21272_);
  or (_21279_, _21278_, _21078_);
  nand (_21281_, _21279_, _05333_);
  and (_21282_, _05329_, _02252_);
  nor (_21283_, _21282_, _02669_);
  and (_21284_, _21283_, _21281_);
  or (_21285_, _21284_, _21077_);
  nand (_21286_, _21285_, _03244_);
  and (_21287_, _03243_, _02251_);
  nor (_21288_, _21287_, _01965_);
  nand (_21289_, _21288_, _21286_);
  nand (_21290_, _21289_, _05343_);
  and (_21292_, _21102_, _05348_);
  nor (_21293_, _02251_, _05348_);
  nor (_21294_, _21293_, _05343_);
  not (_21295_, _21294_);
  nor (_21296_, _21295_, _21292_);
  nor (_21297_, _21296_, _01944_);
  and (_21298_, _21297_, _21290_);
  or (_21299_, _21298_, _21076_);
  nand (_21300_, _21299_, _05358_);
  and (_21301_, _05355_, _02252_);
  nor (_21303_, _21301_, _02654_);
  and (_21304_, _21303_, _21300_);
  or (_21305_, _21304_, _21074_);
  nand (_21306_, _21305_, _05883_);
  and (_21307_, _03239_, _02251_);
  nor (_21308_, _21307_, _01957_);
  nand (_21309_, _21308_, _21306_);
  nand (_21310_, _21309_, _05368_);
  and (_21311_, _02251_, _05348_);
  nor (_21312_, _21102_, _05348_);
  or (_21314_, _21312_, _21311_);
  and (_21315_, _21314_, _05367_);
  nor (_21316_, _21315_, _05391_);
  and (_21317_, _21316_, _21310_);
  or (_21318_, _21317_, _21073_);
  nand (_21319_, _21318_, _05398_);
  and (_21320_, _05393_, _02252_);
  nor (_21321_, _21320_, _05396_);
  nand (_21322_, _21321_, _21319_);
  and (_21323_, _21070_, _05396_);
  nor (_21325_, _21323_, _03109_);
  nand (_21326_, _21325_, _21322_);
  nor (_21327_, _02653_, _01936_);
  not (_21328_, _21327_);
  and (_21329_, _03777_, _03109_);
  nor (_21330_, _21329_, _21328_);
  nand (_21331_, _21330_, _21326_);
  nor (_21332_, _05702_, _02793_);
  and (_21333_, _21091_, _05702_);
  or (_21334_, _21333_, _03267_);
  nor (_21336_, _21334_, _21332_);
  nor (_21337_, _21336_, _05412_);
  and (_21338_, _21337_, _21331_);
  or (_21339_, _21338_, _21072_);
  nand (_21340_, _21339_, _05728_);
  and (_21341_, _05720_, _02252_);
  nor (_21342_, _21341_, _05724_);
  nand (_21343_, _21342_, _21340_);
  and (_21344_, _21070_, _05724_);
  nor (_21345_, _21344_, _03108_);
  nand (_21347_, _21345_, _21343_);
  nor (_21348_, _02647_, _01899_);
  not (_21349_, _21348_);
  and (_21350_, _03777_, _03108_);
  nor (_21351_, _21350_, _21349_);
  nand (_21352_, _21351_, _21347_);
  and (_21353_, _05702_, _02794_);
  nor (_21354_, _21092_, _05702_);
  nor (_21355_, _21354_, _21353_);
  and (_21356_, _21355_, _02647_);
  nor (_21358_, _21356_, _05764_);
  nand (_21359_, _21358_, _21352_);
  and (_21360_, _21075_, _05764_);
  nor (_21361_, _21360_, _03123_);
  nand (_21362_, _21361_, _21359_);
  and (_21363_, _03123_, _02251_);
  nor (_21364_, _21363_, _05780_);
  nand (_21365_, _21364_, _21362_);
  and (_21366_, _21075_, _05780_);
  nor (_21367_, _21366_, _02646_);
  and (_21369_, _21367_, _21365_);
  or (_21370_, _21369_, _21064_);
  nand (_21371_, _21370_, _21040_);
  and (_21372_, _21355_, _02650_);
  nor (_21373_, _21372_, _05826_);
  nand (_21374_, _21373_, _21371_);
  nor (_21375_, _21070_, _05824_);
  nor (_21376_, _21375_, _03121_);
  nand (_21377_, _21376_, _21374_);
  and (_21378_, _03121_, _02251_);
  nor (_21380_, _21378_, _05840_);
  nand (_21381_, _21380_, _21377_);
  and (_21382_, _21075_, _05840_);
  nor (_21383_, _21382_, _02649_);
  and (_21384_, _21383_, _21381_);
  nor (_21385_, _05846_, _02471_);
  or (_21386_, _21385_, _21384_);
  nand (_21387_, _21386_, _21056_);
  and (_21388_, _21070_, _05862_);
  not (_21389_, _21388_);
  and (_21391_, _21389_, _21387_);
  nand (_21392_, _21391_, _27788_);
  or (_21393_, _27788_, \oc8051_golden_model_1.PC [9]);
  and (_21394_, _21393_, _27053_);
  and (_28969_, _21394_, _21392_);
  nor (_21395_, _01906_, \oc8051_golden_model_1.PC [10]);
  nor (_21396_, _21395_, _01907_);
  and (_21397_, _21396_, _05862_);
  not (_21398_, _21397_);
  and (_21399_, _02649_, _02439_);
  nor (_21401_, _21396_, _05824_);
  and (_21402_, _02646_, _02439_);
  not (_21403_, _21396_);
  and (_21404_, _21403_, _05764_);
  and (_21405_, _02778_, _02654_);
  and (_21406_, _02778_, _02669_);
  and (_21407_, _02778_, _02656_);
  and (_21408_, _21396_, _05225_);
  and (_21409_, _21403_, _05000_);
  nor (_21410_, _21403_, _04996_);
  and (_21412_, _04540_, _02238_);
  not (_21413_, _02248_);
  nor (_21414_, _02538_, _02535_);
  nor (_21415_, _21414_, _21413_);
  and (_21416_, _21414_, _21413_);
  nor (_21417_, _21416_, _21415_);
  nand (_21418_, _21417_, _04537_);
  nand (_21419_, _21418_, _03406_);
  or (_21420_, _21419_, _21412_);
  and (_21421_, _21396_, _04502_);
  not (_21423_, _04510_);
  and (_21424_, _04521_, _21423_);
  or (_21425_, _21396_, _21424_);
  or (_21426_, _04520_, \oc8051_golden_model_1.PC [10]);
  or (_21427_, _04512_, _04505_);
  or (_21428_, _21427_, _21426_);
  or (_21429_, _21428_, _18582_);
  and (_21430_, _21429_, _21425_);
  or (_21431_, _21430_, _03154_);
  nor (_21432_, _04505_, _03154_);
  or (_21434_, _21432_, _02238_);
  and (_21435_, _21434_, _18144_);
  and (_21436_, _21435_, _21431_);
  or (_21437_, _21436_, _20763_);
  nor (_21438_, _21437_, _21421_);
  nor (_21439_, _04545_, _02661_);
  not (_21440_, _21439_);
  nor (_21441_, _21440_, _21438_);
  nand (_21442_, _21441_, _21420_);
  or (_21443_, _04987_, _02777_);
  not (_21445_, _02790_);
  nor (_21446_, _03082_, _03079_);
  nor (_21447_, _21446_, _21445_);
  and (_21448_, _21446_, _21445_);
  nor (_21449_, _21448_, _21447_);
  or (_21450_, _21449_, _04985_);
  and (_21451_, _21450_, _02661_);
  nand (_21452_, _21451_, _21443_);
  nand (_21453_, _21452_, _21442_);
  and (_21454_, _21453_, _18134_);
  or (_21456_, _21454_, _21410_);
  nand (_21457_, _21456_, _03163_);
  nor (_21458_, _03163_, _02239_);
  nor (_21459_, _05000_, _07558_);
  not (_21460_, _21459_);
  nor (_21461_, _21460_, _21458_);
  and (_21462_, _21461_, _21457_);
  or (_21463_, _21462_, _21409_);
  nand (_21464_, _21463_, _03179_);
  and (_21465_, _03168_, _02239_);
  nor (_21467_, _21465_, _05009_);
  and (_21468_, _21467_, _21464_);
  and (_21469_, _21396_, _05009_);
  or (_21470_, _21469_, _21468_);
  nand (_21471_, _21470_, _03177_);
  and (_21472_, _21471_, _01990_);
  or (_21473_, _21472_, _03187_);
  or (_21474_, _03428_, _02239_);
  and (_21475_, _21474_, _04499_);
  and (_21476_, _21475_, _21473_);
  not (_21478_, _21449_);
  nor (_21479_, _21478_, _04494_);
  and (_21480_, _04494_, _02777_);
  or (_21481_, _21480_, _04499_);
  nor (_21482_, _21481_, _21479_);
  nor (_21483_, _21482_, _21476_);
  or (_21484_, _21483_, _02675_);
  and (_21485_, _04275_, _02777_);
  and (_21486_, _21449_, _04277_);
  or (_21487_, _21486_, _03107_);
  or (_21489_, _21487_, _21485_);
  nand (_21490_, _21489_, _21484_);
  or (_21491_, _21490_, _02664_);
  and (_21492_, _05157_, _02777_);
  nor (_21493_, _21478_, _05157_);
  nor (_21494_, _21493_, _21492_);
  or (_21495_, _21494_, _03387_);
  and (_21496_, _21495_, _21491_);
  or (_21497_, _21496_, _02673_);
  nand (_21498_, _02777_, _02630_);
  nand (_21500_, _21449_, _19401_);
  and (_21501_, _21500_, _21498_);
  or (_21502_, _21501_, _05024_);
  and (_21503_, _21502_, _21497_);
  or (_21504_, _21503_, _02598_);
  nand (_21505_, _21396_, _02598_);
  and (_21506_, _21505_, _21504_);
  nor (_21507_, _21506_, _03144_);
  and (_21508_, _03144_, _02238_);
  nor (_21509_, _21508_, _21507_);
  and (_21511_, _21509_, _05178_);
  nor (_21512_, _05177_, _02238_);
  or (_21513_, _21512_, _21511_);
  nand (_21514_, _21513_, _05186_);
  and (_21515_, _21403_, _05185_);
  nor (_21516_, _21515_, _03205_);
  nand (_21517_, _21516_, _21514_);
  nand (_21518_, _21517_, _01993_);
  nand (_21519_, _21518_, _18677_);
  nor (_21520_, _03207_, _02239_);
  nor (_21522_, _21520_, _05194_);
  nand (_21523_, _21522_, _21519_);
  and (_21524_, _21403_, _05194_);
  nor (_21525_, _21524_, _05199_);
  and (_21526_, _21525_, _21523_);
  and (_21527_, _05199_, _02238_);
  or (_21528_, _21527_, _02047_);
  or (_21529_, _21528_, _21526_);
  nor (_21530_, _21396_, _01985_);
  nor (_21531_, _21530_, _03140_);
  nand (_21533_, _21531_, _21529_);
  and (_21534_, _03140_, _02238_);
  nor (_21535_, _21534_, _20878_);
  nand (_21536_, _21535_, _21533_);
  and (_21537_, _02778_, _02670_);
  nor (_21538_, _21537_, _05217_);
  nand (_21539_, _21538_, _21536_);
  and (_21540_, _05217_, _02238_);
  nor (_21541_, _21540_, _02024_);
  nand (_21542_, _21541_, _21539_);
  and (_21544_, _02778_, _02024_);
  nor (_21545_, _21544_, _05225_);
  and (_21546_, _21545_, _21542_);
  or (_21547_, _21546_, _21408_);
  nand (_21548_, _21547_, _03462_);
  and (_21549_, _03135_, _02238_);
  not (_21550_, _21549_);
  and (_21551_, _21550_, _20894_);
  nand (_21552_, _21551_, _21548_);
  nor (_21553_, _21417_, _05234_);
  nor (_21555_, _21553_, _02577_);
  and (_21556_, _21555_, _21552_);
  and (_21557_, _02577_, _02238_);
  or (_21558_, _21557_, _02575_);
  or (_21559_, _21558_, _21556_);
  and (_21560_, _02778_, _02575_);
  nor (_21561_, _21560_, _05243_);
  nand (_21562_, _21561_, _21559_);
  and (_21563_, _05243_, _02238_);
  nor (_21564_, _21563_, _02573_);
  nand (_21566_, _21564_, _21562_);
  nor (_21567_, _05279_, \oc8051_golden_model_1.DPH [2]);
  nor (_21568_, _21567_, _05280_);
  nor (_21569_, _21568_, _02574_);
  nor (_21570_, _21569_, _03134_);
  and (_21571_, _21570_, _21566_);
  and (_21572_, _03134_, _02238_);
  or (_21573_, _21572_, _21571_);
  nor (_21574_, _02567_, _01967_);
  nand (_21575_, _21574_, _21573_);
  nor (_21577_, _21417_, _01953_);
  nor (_21578_, _02238_, _02568_);
  nor (_21579_, _21578_, _05291_);
  not (_21580_, _21579_);
  nor (_21581_, _21580_, _21577_);
  nor (_21582_, _21581_, _05297_);
  nand (_21583_, _21582_, _21575_);
  and (_21584_, _21403_, _05297_);
  nor (_21585_, _21584_, _05302_);
  nand (_21586_, _21585_, _21583_);
  and (_21588_, _05302_, _02238_);
  nor (_21589_, _21588_, _02656_);
  and (_21590_, _21589_, _21586_);
  or (_21591_, _21590_, _21407_);
  or (_21592_, _21591_, _03251_);
  nand (_21593_, _03251_, _02238_);
  and (_21594_, _21593_, _21592_);
  or (_21595_, _21594_, _01974_);
  or (_21596_, _21595_, _05315_);
  nor (_21597_, _21417_, _02568_);
  nor (_21599_, _02238_, _01953_);
  nor (_21600_, _21599_, _05316_);
  not (_21601_, _21600_);
  nor (_21602_, _21601_, _21597_);
  nor (_21603_, _21602_, _05325_);
  nand (_21604_, _21603_, _21596_);
  and (_21605_, _21403_, _05325_);
  nor (_21606_, _21605_, _05329_);
  nand (_21607_, _21606_, _21604_);
  and (_21608_, _05329_, _02238_);
  nor (_21610_, _21608_, _02669_);
  and (_21611_, _21610_, _21607_);
  or (_21612_, _21611_, _21406_);
  nand (_21613_, _21612_, _03244_);
  and (_21614_, _03243_, _02239_);
  nor (_21615_, _21614_, _20957_);
  nand (_21616_, _21615_, _21613_);
  nor (_21617_, _21417_, \oc8051_golden_model_1.PSW [7]);
  nor (_21618_, _02238_, _05348_);
  nor (_21619_, _21618_, _05343_);
  not (_21621_, _21619_);
  nor (_21622_, _21621_, _21617_);
  nor (_21623_, _21622_, _01944_);
  nand (_21624_, _21623_, _21616_);
  and (_21625_, _21403_, _01944_);
  nor (_21626_, _21625_, _05355_);
  nand (_21627_, _21626_, _21624_);
  and (_21628_, _05355_, _02238_);
  nor (_21629_, _21628_, _02654_);
  and (_21630_, _21629_, _21627_);
  or (_21632_, _21630_, _21405_);
  nand (_21633_, _21632_, _05883_);
  and (_21634_, _03239_, _02239_);
  nor (_21635_, _21634_, _20979_);
  nand (_21636_, _21635_, _21633_);
  and (_21637_, _02238_, _05348_);
  and (_21638_, _21417_, \oc8051_golden_model_1.PSW [7]);
  or (_21639_, _21638_, _21637_);
  and (_21640_, _21639_, _05367_);
  nor (_21641_, _21640_, _05391_);
  nand (_21643_, _21641_, _21636_);
  nor (_21644_, _21396_, _05389_);
  nor (_21645_, _21644_, _05393_);
  and (_21646_, _21645_, _21643_);
  and (_21647_, _05393_, _02238_);
  or (_21648_, _21647_, _21646_);
  and (_21649_, _21648_, _05397_);
  and (_21650_, _21396_, _05396_);
  or (_21651_, _21650_, _03109_);
  or (_21652_, _21651_, _21649_);
  and (_21654_, _03644_, _03109_);
  nor (_21655_, _21654_, _21328_);
  nand (_21656_, _21655_, _21652_);
  and (_21657_, _21478_, _05702_);
  nor (_21658_, _05702_, _02777_);
  or (_21659_, _21658_, _03267_);
  or (_21660_, _21659_, _21657_);
  and (_21661_, _21660_, _01930_);
  nand (_21662_, _21661_, _21656_);
  nor (_21663_, _21396_, _01930_);
  nor (_21665_, _21663_, _05720_);
  and (_21666_, _21665_, _21662_);
  and (_21667_, _05720_, _02238_);
  or (_21668_, _21667_, _21666_);
  and (_21669_, _21668_, _05726_);
  and (_21670_, _21396_, _05724_);
  or (_21671_, _21670_, _03108_);
  or (_21672_, _21671_, _21669_);
  and (_21673_, _03644_, _03108_);
  nor (_21674_, _21673_, _21349_);
  nand (_21676_, _21674_, _21672_);
  nor (_21677_, _21449_, _05702_);
  and (_21678_, _05702_, _02778_);
  nor (_21679_, _21678_, _21677_);
  and (_21680_, _21679_, _02647_);
  nor (_21681_, _21680_, _05764_);
  and (_21682_, _21681_, _21676_);
  or (_21683_, _21682_, _21404_);
  nand (_21684_, _21683_, _03124_);
  and (_21685_, _03123_, _02239_);
  nor (_21687_, _21685_, _05780_);
  nand (_21688_, _21687_, _21684_);
  and (_21689_, _21396_, _05780_);
  nor (_21690_, _21689_, _02646_);
  nand (_21691_, _21690_, _21688_);
  nand (_21692_, _21691_, _21040_);
  or (_21693_, _21692_, _21402_);
  and (_21694_, _21679_, _02650_);
  nor (_21695_, _21694_, _05826_);
  and (_21696_, _21695_, _21693_);
  or (_21698_, _21696_, _21401_);
  nand (_21699_, _21698_, _03513_);
  and (_21700_, _03121_, _02239_);
  nor (_21701_, _21700_, _05840_);
  nand (_21702_, _21701_, _21699_);
  and (_21703_, _21396_, _05840_);
  nor (_21704_, _21703_, _02649_);
  nand (_21705_, _21704_, _21702_);
  nand (_21706_, _21705_, _21056_);
  or (_21707_, _21706_, _21399_);
  and (_21709_, _21707_, _21398_);
  nand (_21710_, _21709_, _27788_);
  or (_21711_, _27788_, \oc8051_golden_model_1.PC [10]);
  and (_21712_, _21711_, _27053_);
  and (_28970_, _21712_, _21710_);
  nand (_21713_, _03859_, _03108_);
  nor (_21714_, _01907_, \oc8051_golden_model_1.PC [11]);
  nor (_21715_, _21714_, _01908_);
  or (_21716_, _21715_, _01930_);
  nand (_21717_, _03859_, _03109_);
  nor (_21719_, _21415_, _02240_);
  and (_21720_, _21719_, _02246_);
  nor (_21721_, _21719_, _02246_);
  or (_21722_, _21721_, _21720_);
  or (_21723_, _21722_, _05348_);
  or (_21724_, _02243_, \oc8051_golden_model_1.PSW [7]);
  and (_21725_, _21724_, _05367_);
  and (_21726_, _21725_, _21723_);
  or (_21727_, _21715_, _01945_);
  or (_21728_, _21722_, _02568_);
  or (_21730_, _02243_, _01953_);
  and (_21731_, _21730_, _05315_);
  and (_21732_, _21731_, _21728_);
  or (_21733_, _21715_, _05298_);
  or (_21734_, _08748_, _02243_);
  nor (_21735_, _21447_, _02779_);
  and (_21736_, _21735_, _02788_);
  nor (_21737_, _21735_, _02788_);
  or (_21738_, _21737_, _21736_);
  or (_21739_, _21738_, _02630_);
  nand (_21741_, _02785_, _02630_);
  and (_21742_, _21741_, _02673_);
  and (_21743_, _21742_, _21739_);
  and (_21744_, _21738_, _04277_);
  and (_21745_, _04275_, _02784_);
  or (_21746_, _21745_, _21744_);
  or (_21747_, _21746_, _03107_);
  or (_21748_, _21738_, _04494_);
  nand (_21749_, _04494_, _02785_);
  and (_21750_, _21749_, _21748_);
  or (_21752_, _21750_, _04499_);
  and (_21753_, _03168_, _02243_);
  or (_21754_, _21715_, _18144_);
  or (_21755_, _21715_, _21423_);
  or (_21756_, _21715_, _04521_);
  nor (_21757_, _04505_, \oc8051_golden_model_1.PC [11]);
  nand (_21758_, _21757_, _04521_);
  or (_21759_, _21758_, _17874_);
  and (_21760_, _21759_, _21756_);
  or (_21761_, _21760_, _04504_);
  and (_21763_, _21761_, _21755_);
  or (_21764_, _21763_, _03154_);
  and (_21765_, _21764_, _21754_);
  or (_21766_, _21765_, _04527_);
  and (_21767_, _04507_, _01998_);
  or (_21768_, _21767_, _02243_);
  and (_21769_, _21768_, _21766_);
  or (_21770_, _21769_, _03406_);
  and (_21771_, _21722_, _04537_);
  and (_21772_, _04540_, _02243_);
  or (_21774_, _21772_, _04539_);
  or (_21775_, _21774_, _21771_);
  and (_21776_, _21775_, _21770_);
  or (_21777_, _21776_, _04545_);
  and (_21778_, _21777_, _02662_);
  or (_21779_, _21738_, _04985_);
  or (_21780_, _04987_, _02784_);
  and (_21781_, _21780_, _02661_);
  and (_21782_, _21781_, _21779_);
  or (_21783_, _21782_, _04992_);
  or (_21785_, _21783_, _21778_);
  or (_21786_, _21715_, _04996_);
  and (_21787_, _21786_, _04995_);
  and (_21788_, _21787_, _21785_);
  not (_21789_, _04995_);
  and (_21790_, _21789_, _02243_);
  or (_21791_, _21790_, _05000_);
  or (_21792_, _21791_, _21788_);
  or (_21793_, _21715_, _05004_);
  and (_21794_, _21793_, _03179_);
  and (_21796_, _21794_, _21792_);
  or (_21797_, _21796_, _21753_);
  and (_21798_, _21797_, _05010_);
  nand (_21799_, _21715_, _05009_);
  nand (_21800_, _21799_, _05013_);
  or (_21801_, _21800_, _21798_);
  or (_21802_, _05013_, _02243_);
  and (_21803_, _21802_, _21801_);
  or (_21804_, _21803_, _04498_);
  and (_21805_, _21804_, _21752_);
  or (_21807_, _21805_, _02675_);
  and (_21808_, _21807_, _21747_);
  or (_21809_, _21808_, _02664_);
  and (_21810_, _05157_, _02784_);
  and (_21811_, _21738_, _05158_);
  or (_21812_, _21811_, _03387_);
  or (_21813_, _21812_, _21810_);
  and (_21814_, _21813_, _05024_);
  and (_21815_, _21814_, _21809_);
  or (_21816_, _21815_, _21743_);
  and (_21818_, _21816_, _02599_);
  nand (_21819_, _21715_, _02598_);
  nand (_21820_, _21819_, _05179_);
  or (_21821_, _21820_, _21818_);
  or (_21822_, _05179_, _02243_);
  and (_21823_, _21822_, _05186_);
  and (_21824_, _21823_, _21821_);
  and (_21825_, _21715_, _05185_);
  or (_21826_, _21825_, _05191_);
  or (_21827_, _21826_, _21824_);
  or (_21829_, _05190_, _02243_);
  and (_21830_, _21829_, _05195_);
  and (_21831_, _21830_, _21827_);
  and (_21832_, _21715_, _05194_);
  or (_21833_, _21832_, _05199_);
  or (_21834_, _21833_, _21831_);
  or (_21835_, _05203_, _02243_);
  and (_21836_, _21835_, _01985_);
  and (_21837_, _21836_, _21834_);
  nand (_21838_, _21715_, _02047_);
  nand (_21840_, _21838_, _05208_);
  or (_21841_, _21840_, _21837_);
  or (_21842_, _05208_, _02243_);
  and (_21843_, _21842_, _05212_);
  and (_21844_, _21843_, _21841_);
  and (_21845_, _02784_, _02670_);
  or (_21846_, _21845_, _05217_);
  or (_21847_, _21846_, _21844_);
  or (_21848_, _05220_, _02243_);
  and (_21849_, _21848_, _03139_);
  and (_21851_, _21849_, _21847_);
  or (_21852_, _05225_, _02784_);
  and (_21853_, _21852_, _17972_);
  or (_21854_, _21853_, _21851_);
  or (_21855_, _21715_, _05226_);
  and (_21856_, _21855_, _21854_);
  or (_21857_, _21856_, _05229_);
  or (_21858_, _05228_, _02243_);
  and (_21859_, _21858_, _05234_);
  and (_21860_, _21859_, _21857_);
  and (_21862_, _21722_, _05233_);
  or (_21863_, _21862_, _02577_);
  or (_21864_, _21863_, _21860_);
  and (_21865_, _21864_, _21734_);
  or (_21866_, _21865_, _02575_);
  nand (_21867_, _02785_, _02575_);
  and (_21868_, _21867_, _05244_);
  and (_21869_, _21868_, _21866_);
  and (_21870_, _05243_, _02243_);
  or (_21871_, _21870_, _21869_);
  and (_21873_, _21871_, _02574_);
  or (_21874_, _05280_, \oc8051_golden_model_1.DPH [3]);
  nor (_21875_, _05281_, _02574_);
  and (_21876_, _21875_, _21874_);
  or (_21877_, _21876_, _05253_);
  or (_21878_, _21877_, _21873_);
  or (_21879_, _05252_, _02243_);
  and (_21880_, _21879_, _05291_);
  and (_21881_, _21880_, _21878_);
  or (_21882_, _21722_, _01953_);
  or (_21884_, _02243_, _02568_);
  and (_21885_, _21884_, _02567_);
  and (_21886_, _21885_, _21882_);
  or (_21887_, _21886_, _05297_);
  or (_21888_, _21887_, _21881_);
  and (_21889_, _21888_, _21733_);
  or (_21890_, _21889_, _05302_);
  or (_21891_, _05306_, _02243_);
  and (_21892_, _21891_, _05305_);
  and (_21893_, _21892_, _21890_);
  nand (_21895_, _02784_, _02656_);
  nand (_21896_, _21895_, _05311_);
  or (_21897_, _21896_, _21893_);
  or (_21898_, _05311_, _02243_);
  and (_21899_, _21898_, _05316_);
  and (_21900_, _21899_, _21897_);
  or (_21901_, _21900_, _21732_);
  and (_21902_, _21901_, _05326_);
  and (_21903_, _21715_, _05325_);
  or (_21904_, _21903_, _05329_);
  or (_21906_, _21904_, _21902_);
  or (_21907_, _05333_, _02243_);
  and (_21908_, _21907_, _05332_);
  and (_21909_, _21908_, _21906_);
  nand (_21910_, _02784_, _02669_);
  nand (_21911_, _21910_, _05338_);
  or (_21912_, _21911_, _21909_);
  or (_21913_, _05338_, _02243_);
  and (_21914_, _21913_, _05343_);
  and (_21915_, _21914_, _21912_);
  or (_21917_, _21722_, \oc8051_golden_model_1.PSW [7]);
  or (_21918_, _02243_, _05348_);
  and (_21919_, _21918_, _05342_);
  and (_21920_, _21919_, _21917_);
  or (_21921_, _21920_, _01944_);
  or (_21922_, _21921_, _21915_);
  and (_21923_, _21922_, _21727_);
  or (_21924_, _21923_, _05355_);
  or (_21925_, _05358_, _02243_);
  and (_21926_, _21925_, _05357_);
  and (_21928_, _21926_, _21924_);
  nand (_21929_, _02784_, _02654_);
  nand (_21930_, _21929_, _05363_);
  or (_21931_, _21930_, _21928_);
  or (_21932_, _05363_, _02243_);
  and (_21933_, _21932_, _05368_);
  and (_21934_, _21933_, _21931_);
  or (_21935_, _21934_, _21726_);
  and (_21936_, _21935_, _05389_);
  and (_21937_, _21715_, _05391_);
  or (_21939_, _21937_, _05393_);
  or (_21940_, _21939_, _21936_);
  or (_21941_, _05398_, _02243_);
  and (_21942_, _21941_, _05397_);
  and (_21943_, _21942_, _21940_);
  and (_21944_, _21715_, _05396_);
  or (_21945_, _21944_, _03109_);
  or (_21946_, _21945_, _21943_);
  and (_21947_, _21946_, _21717_);
  or (_21948_, _21947_, _01936_);
  or (_21950_, _02243_, _05408_);
  and (_21951_, _21950_, _03267_);
  and (_21952_, _21951_, _21948_);
  or (_21953_, _21738_, _05704_);
  or (_21954_, _05702_, _02784_);
  and (_21955_, _21954_, _02653_);
  and (_21956_, _21955_, _21953_);
  or (_21957_, _21956_, _05412_);
  or (_21958_, _21957_, _21952_);
  and (_21959_, _21958_, _21716_);
  or (_21961_, _21959_, _05720_);
  or (_21962_, _05728_, _02243_);
  and (_21963_, _21962_, _05726_);
  and (_21964_, _21963_, _21961_);
  and (_21965_, _21715_, _05724_);
  or (_21966_, _21965_, _03108_);
  or (_21967_, _21966_, _21964_);
  and (_21968_, _21967_, _21713_);
  or (_21969_, _21968_, _01899_);
  or (_21970_, _02243_, _05748_);
  and (_21972_, _21970_, _03125_);
  and (_21973_, _21972_, _21969_);
  or (_21974_, _21738_, _05702_);
  nand (_21975_, _05702_, _02785_);
  and (_21976_, _21975_, _21974_);
  and (_21977_, _21976_, _02647_);
  or (_21978_, _21977_, _05764_);
  or (_21979_, _21978_, _21973_);
  or (_21980_, _21715_, _05770_);
  and (_21981_, _21980_, _03124_);
  and (_21983_, _21981_, _21979_);
  and (_21984_, _03123_, _02243_);
  or (_21985_, _21984_, _05780_);
  or (_21986_, _21985_, _21983_);
  or (_21987_, _21715_, _05788_);
  and (_21988_, _21987_, _05786_);
  and (_21989_, _21988_, _21986_);
  and (_21990_, _02646_, _02405_);
  or (_21991_, _21990_, _01971_);
  or (_21992_, _21991_, _21989_);
  or (_21994_, _02243_, _05802_);
  and (_21995_, _21994_, _03122_);
  and (_21996_, _21995_, _21992_);
  and (_21997_, _21976_, _02650_);
  or (_21998_, _21997_, _05826_);
  or (_21999_, _21998_, _21996_);
  or (_22000_, _21715_, _05824_);
  and (_22001_, _22000_, _03513_);
  and (_22002_, _22001_, _21999_);
  and (_22003_, _03121_, _02243_);
  or (_22005_, _22003_, _05840_);
  or (_22006_, _22005_, _22002_);
  or (_22007_, _21715_, _05848_);
  and (_22008_, _22007_, _05846_);
  and (_22009_, _22008_, _22006_);
  and (_22010_, _02649_, _02405_);
  or (_22011_, _22010_, _01955_);
  or (_22012_, _22011_, _22009_);
  or (_22013_, _02243_, _01956_);
  and (_22014_, _22013_, _05864_);
  and (_22016_, _22014_, _22012_);
  and (_22017_, _21715_, _05862_);
  or (_22018_, _22017_, _22016_);
  or (_22019_, _22018_, _27789_);
  or (_22020_, _27788_, \oc8051_golden_model_1.PC [11]);
  and (_22021_, _22020_, _27053_);
  and (_28971_, _22021_, _22019_);
  and (_22022_, _02234_, _05348_);
  and (_22023_, _02545_, _02542_);
  nor (_22024_, _22023_, _02546_);
  and (_22026_, _22024_, \oc8051_golden_model_1.PSW [7]);
  or (_22027_, _22026_, _22022_);
  and (_22028_, _22027_, _05367_);
  and (_22029_, _02577_, _02235_);
  and (_22030_, _02773_, _02024_);
  and (_22031_, _05157_, _02773_);
  and (_22032_, _03089_, _03086_);
  nor (_22033_, _22032_, _03090_);
  not (_22034_, _22033_);
  nor (_22035_, _22034_, _05157_);
  nor (_22037_, _22035_, _22031_);
  or (_22038_, _22037_, _03387_);
  and (_22039_, _22033_, _04277_);
  and (_22040_, _04275_, _02773_);
  or (_22041_, _22040_, _22039_);
  nor (_22042_, _22041_, _03107_);
  and (_22043_, _04494_, _02773_);
  nor (_22044_, _22034_, _04494_);
  or (_22045_, _22044_, _22043_);
  nor (_22046_, _22045_, _04499_);
  and (_22048_, _20364_, _02206_);
  and (_22049_, _22048_, \oc8051_golden_model_1.PC [11]);
  and (_22050_, _22049_, \oc8051_golden_model_1.PC [12]);
  nor (_22051_, _22049_, \oc8051_golden_model_1.PC [12]);
  nor (_22052_, _22051_, _22050_);
  nor (_22053_, _22052_, _04996_);
  or (_22054_, _21767_, _02234_);
  not (_22055_, _22052_);
  and (_22056_, _22055_, _04502_);
  nor (_22057_, _22052_, _21424_);
  nor (_22059_, _04504_, \oc8051_golden_model_1.PC [12]);
  and (_22060_, _22059_, _05903_);
  and (_22061_, _22060_, _04523_);
  or (_22062_, _22061_, _22057_);
  and (_22063_, _22062_, _04503_);
  nor (_22064_, _22063_, _22056_);
  or (_22065_, _22064_, _04527_);
  and (_22066_, _22065_, _22054_);
  nor (_22067_, _22066_, _03406_);
  and (_22068_, _04540_, _02234_);
  and (_22070_, _22024_, _04537_);
  or (_22071_, _22070_, _22068_);
  nor (_22072_, _22071_, _04539_);
  nor (_22073_, _22072_, _22067_);
  nor (_22074_, _22073_, _04545_);
  nor (_22075_, _22074_, _02661_);
  not (_22076_, _22075_);
  and (_22077_, _22033_, _04987_);
  and (_22078_, _04985_, _02773_);
  nor (_22079_, _22078_, _22077_);
  nor (_22081_, _22079_, _02662_);
  nor (_22082_, _22081_, _04992_);
  and (_22083_, _22082_, _22076_);
  nor (_22084_, _22083_, _22053_);
  nor (_22085_, _22084_, _21789_);
  nor (_22086_, _04995_, _02234_);
  nor (_22087_, _22086_, _05000_);
  not (_22088_, _22087_);
  nor (_22089_, _22088_, _22085_);
  and (_22090_, _22052_, _05000_);
  nor (_22092_, _22090_, _03168_);
  not (_22093_, _22092_);
  nor (_22094_, _22093_, _22089_);
  and (_22095_, _03168_, _02235_);
  nor (_22096_, _22095_, _05009_);
  not (_22097_, _22096_);
  nor (_22098_, _22097_, _22094_);
  and (_22099_, _22052_, _05009_);
  nor (_22100_, _22099_, _05014_);
  not (_22101_, _22100_);
  nor (_22103_, _22101_, _22098_);
  nor (_22104_, _05013_, _02234_);
  nor (_22105_, _22104_, _22103_);
  nor (_22106_, _22105_, _04498_);
  nor (_22107_, _22106_, _22046_);
  nor (_22108_, _22107_, _02675_);
  nor (_22109_, _22108_, _22042_);
  nand (_22110_, _22109_, _03387_);
  and (_22111_, _22110_, _22038_);
  or (_22112_, _22111_, _02673_);
  nand (_22114_, _02773_, _02630_);
  nand (_22115_, _22033_, _19401_);
  and (_22116_, _22115_, _22114_);
  or (_22117_, _22116_, _05024_);
  nand (_22118_, _22117_, _22112_);
  nand (_22119_, _22118_, _02599_);
  and (_22120_, _22052_, _02598_);
  not (_22121_, _22120_);
  and (_22122_, _22121_, _05179_);
  nand (_22123_, _22122_, _22119_);
  nor (_22125_, _05179_, _02234_);
  nor (_22126_, _22125_, _05185_);
  nand (_22127_, _22126_, _22123_);
  and (_22128_, _22052_, _05185_);
  nor (_22129_, _22128_, _05191_);
  nand (_22130_, _22129_, _22127_);
  nor (_22131_, _05190_, _02234_);
  nor (_22132_, _22131_, _05194_);
  nand (_22133_, _22132_, _22130_);
  and (_22134_, _22052_, _05194_);
  nor (_22136_, _22134_, _05199_);
  nand (_22137_, _22136_, _22133_);
  and (_22138_, _05199_, _02235_);
  nor (_22139_, _22138_, _02047_);
  nand (_22140_, _22139_, _22137_);
  nor (_22141_, _22055_, _01985_);
  nor (_22142_, _22141_, _05209_);
  nand (_22143_, _22142_, _22140_);
  nor (_22144_, _05208_, _02234_);
  nor (_22145_, _22144_, _02670_);
  nand (_22147_, _22145_, _22143_);
  and (_22148_, _02773_, _02670_);
  nor (_22149_, _22148_, _05217_);
  nand (_22150_, _22149_, _22147_);
  and (_22151_, _05217_, _02235_);
  nor (_22152_, _22151_, _02024_);
  and (_22153_, _22152_, _22150_);
  or (_22154_, _22153_, _22030_);
  nand (_22155_, _22154_, _05226_);
  and (_22156_, _22052_, _05225_);
  nor (_22158_, _22156_, _05229_);
  nand (_22159_, _22158_, _22155_);
  nor (_22160_, _05228_, _02234_);
  nor (_22161_, _22160_, _05233_);
  nand (_22162_, _22161_, _22159_);
  and (_22163_, _22024_, _05233_);
  nor (_22164_, _22163_, _02577_);
  and (_22165_, _22164_, _22162_);
  or (_22166_, _22165_, _22029_);
  nand (_22167_, _22166_, _05245_);
  and (_22169_, _02774_, _02575_);
  nor (_22170_, _22169_, _05243_);
  and (_22171_, _22170_, _22167_);
  and (_22172_, _05243_, _02234_);
  or (_22173_, _22172_, _22171_);
  nand (_22174_, _22173_, _02574_);
  nor (_22175_, _05281_, \oc8051_golden_model_1.DPH [4]);
  or (_22176_, _05282_, _02574_);
  or (_22177_, _22176_, _22175_);
  and (_22178_, _22177_, _05252_);
  nand (_22180_, _22178_, _22174_);
  nor (_22181_, _05252_, _02234_);
  nor (_22182_, _22181_, _02567_);
  nand (_22183_, _22182_, _22180_);
  nand (_22184_, _02234_, _01953_);
  nand (_22185_, _22024_, _02568_);
  and (_22186_, _22185_, _22184_);
  or (_22187_, _22186_, _05291_);
  nand (_22188_, _22187_, _22183_);
  nand (_22189_, _22188_, _05298_);
  and (_22191_, _22052_, _05297_);
  nor (_22192_, _22191_, _05302_);
  nand (_22193_, _22192_, _22189_);
  and (_22194_, _05302_, _02235_);
  nor (_22195_, _22194_, _02656_);
  nand (_22196_, _22195_, _22193_);
  and (_22197_, _02773_, _02656_);
  nor (_22198_, _22197_, _05312_);
  nand (_22199_, _22198_, _22196_);
  nor (_22200_, _05311_, _02234_);
  nor (_22202_, _22200_, _05315_);
  nand (_22203_, _22202_, _22199_);
  nand (_22204_, _02234_, _02568_);
  nand (_22205_, _22024_, _01953_);
  and (_22206_, _22205_, _22204_);
  or (_22207_, _22206_, _05316_);
  nand (_22208_, _22207_, _22203_);
  nand (_22209_, _22208_, _05326_);
  and (_22210_, _22052_, _05325_);
  nor (_22211_, _22210_, _05329_);
  nand (_22213_, _22211_, _22209_);
  and (_22214_, _05329_, _02235_);
  nor (_22215_, _22214_, _02669_);
  nand (_22216_, _22215_, _22213_);
  and (_22217_, _02773_, _02669_);
  nor (_22218_, _22217_, _05339_);
  nand (_22219_, _22218_, _22216_);
  nor (_22220_, _05338_, _02234_);
  nor (_22221_, _22220_, _05342_);
  nand (_22222_, _22221_, _22219_);
  nand (_22224_, _02234_, \oc8051_golden_model_1.PSW [7]);
  nand (_22225_, _22024_, _05348_);
  and (_22226_, _22225_, _22224_);
  or (_22227_, _22226_, _05343_);
  nand (_22228_, _22227_, _22222_);
  nand (_22229_, _22228_, _01945_);
  and (_22230_, _22052_, _01944_);
  nor (_22231_, _22230_, _05355_);
  nand (_22232_, _22231_, _22229_);
  and (_22233_, _05355_, _02235_);
  nor (_22235_, _22233_, _02654_);
  nand (_22236_, _22235_, _22232_);
  and (_22237_, _02773_, _02654_);
  nor (_22238_, _22237_, _05364_);
  nand (_22239_, _22238_, _22236_);
  nor (_22240_, _05363_, _02234_);
  nor (_22241_, _22240_, _05367_);
  and (_22242_, _22241_, _22239_);
  or (_22243_, _22242_, _22028_);
  nand (_22244_, _22243_, _05389_);
  nor (_22246_, _22055_, _05389_);
  nor (_22247_, _22246_, _05393_);
  nand (_22248_, _22247_, _22244_);
  and (_22249_, _05393_, _02235_);
  nor (_22250_, _22249_, _05396_);
  nand (_22251_, _22250_, _22248_);
  and (_22252_, _22052_, _05396_);
  nor (_22253_, _22252_, _03109_);
  and (_22254_, _22253_, _22251_);
  and (_22255_, _04325_, _03109_);
  or (_22257_, _22255_, _22254_);
  nand (_22258_, _22257_, _05408_);
  and (_22259_, _02235_, _01936_);
  nor (_22260_, _22259_, _02653_);
  and (_22261_, _22260_, _22258_);
  and (_22262_, _22033_, _05702_);
  nor (_22263_, _05702_, _02774_);
  nor (_22264_, _22263_, _22262_);
  nor (_22265_, _22264_, _03267_);
  or (_22266_, _22265_, _22261_);
  nand (_22268_, _22266_, _01930_);
  nor (_22269_, _22055_, _01930_);
  nor (_22270_, _22269_, _05720_);
  nand (_22271_, _22270_, _22268_);
  and (_22272_, _05720_, _02235_);
  nor (_22273_, _22272_, _05724_);
  nand (_22274_, _22273_, _22271_);
  and (_22275_, _22052_, _05724_);
  nor (_22276_, _22275_, _03108_);
  nand (_22277_, _22276_, _22274_);
  and (_22279_, _04325_, _03108_);
  nor (_22280_, _22279_, _01899_);
  and (_22281_, _22280_, _22277_);
  and (_22282_, _02234_, _01899_);
  or (_22283_, _22282_, _02647_);
  or (_22284_, _22283_, _22281_);
  nor (_22285_, _22033_, _05702_);
  and (_22286_, _05702_, _02774_);
  nor (_22287_, _22286_, _22285_);
  nor (_22288_, _22287_, _03125_);
  nor (_22290_, _22288_, _05764_);
  and (_22291_, _22290_, _22284_);
  and (_22292_, _22052_, _05764_);
  or (_22293_, _22292_, _03123_);
  nor (_22294_, _22293_, _22291_);
  and (_22295_, _03123_, _02235_);
  or (_22296_, _22295_, _22294_);
  and (_22297_, _22296_, _05788_);
  and (_22298_, _22055_, _05780_);
  or (_22299_, _22298_, _22297_);
  nand (_22301_, _22299_, _05786_);
  and (_22302_, _02646_, _02370_);
  nor (_22303_, _22302_, _01971_);
  and (_22304_, _22303_, _22301_);
  and (_22305_, _02234_, _01971_);
  or (_22306_, _22305_, _02650_);
  nor (_22307_, _22306_, _22304_);
  nor (_22308_, _22287_, _03122_);
  or (_22309_, _22308_, _22307_);
  and (_22310_, _22309_, _05824_);
  nor (_22312_, _22052_, _05824_);
  or (_22313_, _22312_, _22310_);
  nand (_22314_, _22313_, _03513_);
  and (_22315_, _03121_, _02235_);
  nor (_22316_, _22315_, _05840_);
  nand (_22317_, _22316_, _22314_);
  and (_22318_, _22052_, _05840_);
  nor (_22319_, _22318_, _02649_);
  and (_22320_, _22319_, _22317_);
  and (_22321_, _02649_, _02370_);
  or (_22323_, _22321_, _22320_);
  nand (_22324_, _22323_, _01956_);
  and (_22325_, _02235_, _01955_);
  nor (_22326_, _22325_, _05862_);
  nand (_22327_, _22326_, _22324_);
  and (_22328_, _22052_, _05862_);
  not (_22329_, _22328_);
  and (_22330_, _22329_, _22327_);
  nand (_22331_, _22330_, _27788_);
  or (_22332_, _27788_, \oc8051_golden_model_1.PC [12]);
  and (_22334_, _22332_, _27053_);
  and (_28972_, _22334_, _22331_);
  nand (_22335_, _04480_, _03108_);
  nor (_22336_, _01909_, \oc8051_golden_model_1.PC [13]);
  nor (_22337_, _22336_, _01910_);
  or (_22338_, _22337_, _01930_);
  or (_22339_, _22337_, _01945_);
  or (_22340_, _22337_, _05326_);
  or (_22341_, _22337_, _05298_);
  or (_22342_, _08748_, _02230_);
  or (_22344_, _02771_, _02770_);
  nand (_22345_, _22344_, _03091_);
  or (_22346_, _22344_, _03091_);
  and (_22347_, _22346_, _22345_);
  and (_22348_, _22347_, _04277_);
  and (_22349_, _04275_, _02768_);
  or (_22350_, _22349_, _22348_);
  or (_22351_, _22350_, _03107_);
  or (_22352_, _22347_, _04494_);
  nand (_22353_, _04494_, _02769_);
  and (_22355_, _22353_, _22352_);
  or (_22356_, _22355_, _04499_);
  and (_22357_, _03168_, _02230_);
  or (_22358_, _21767_, _02230_);
  or (_22359_, _22337_, _04523_);
  or (_22360_, _04520_, _04502_);
  or (_22361_, _22360_, _21427_);
  nand (_22362_, _01988_, _02761_);
  or (_22363_, _22362_, _04511_);
  or (_22364_, _22363_, _22361_);
  and (_22366_, _22364_, _22359_);
  or (_22367_, _22366_, _04527_);
  and (_22368_, _22367_, _22358_);
  or (_22369_, _22368_, _03406_);
  or (_22370_, _02232_, _02231_);
  nand (_22371_, _22370_, _02547_);
  or (_22372_, _22370_, _02547_);
  and (_22373_, _22372_, _22371_);
  and (_22374_, _22373_, _04537_);
  and (_22375_, _04540_, _02230_);
  or (_22377_, _22375_, _04539_);
  or (_22378_, _22377_, _22374_);
  and (_22379_, _22378_, _22369_);
  or (_22380_, _22379_, _04545_);
  and (_22381_, _22380_, _02662_);
  or (_22382_, _22347_, _04985_);
  or (_22383_, _04987_, _02768_);
  and (_22384_, _22383_, _02661_);
  and (_22385_, _22384_, _22382_);
  or (_22386_, _22385_, _04992_);
  or (_22388_, _22386_, _22381_);
  or (_22389_, _22337_, _04996_);
  and (_22390_, _22389_, _04995_);
  and (_22391_, _22390_, _22388_);
  and (_22392_, _21789_, _02230_);
  or (_22393_, _22392_, _05000_);
  or (_22394_, _22393_, _22391_);
  or (_22395_, _22337_, _05004_);
  and (_22396_, _22395_, _03179_);
  and (_22397_, _22396_, _22394_);
  or (_22399_, _22397_, _22357_);
  and (_22400_, _22399_, _05010_);
  nand (_22401_, _22337_, _05009_);
  nand (_22402_, _22401_, _05013_);
  or (_22403_, _22402_, _22400_);
  or (_22404_, _05013_, _02230_);
  and (_22405_, _22404_, _22403_);
  or (_22406_, _22405_, _04498_);
  and (_22407_, _22406_, _22356_);
  or (_22408_, _22407_, _02675_);
  and (_22410_, _22408_, _22351_);
  or (_22411_, _22410_, _02664_);
  and (_22412_, _22347_, _05158_);
  and (_22413_, _05157_, _02768_);
  or (_22414_, _22413_, _03387_);
  or (_22415_, _22414_, _22412_);
  and (_22416_, _22415_, _05024_);
  and (_22417_, _22416_, _22411_);
  or (_22418_, _22347_, _02630_);
  nand (_22419_, _02769_, _02630_);
  and (_22421_, _22419_, _02673_);
  and (_22422_, _22421_, _22418_);
  or (_22423_, _22422_, _22417_);
  and (_22424_, _22423_, _02599_);
  nand (_22425_, _22337_, _02598_);
  nand (_22426_, _22425_, _05179_);
  or (_22427_, _22426_, _22424_);
  or (_22428_, _05179_, _02230_);
  and (_22429_, _22428_, _05186_);
  and (_22430_, _22429_, _22427_);
  and (_22432_, _22337_, _05185_);
  or (_22433_, _22432_, _05191_);
  or (_22434_, _22433_, _22430_);
  or (_22435_, _05190_, _02230_);
  and (_22436_, _22435_, _05195_);
  and (_22437_, _22436_, _22434_);
  and (_22438_, _22337_, _05194_);
  or (_22439_, _22438_, _05199_);
  or (_22440_, _22439_, _22437_);
  or (_22441_, _05203_, _02230_);
  and (_22443_, _22441_, _01985_);
  and (_22444_, _22443_, _22440_);
  and (_22445_, _22337_, _02047_);
  or (_22446_, _22445_, _05209_);
  or (_22447_, _22446_, _22444_);
  or (_22448_, _05208_, _02230_);
  and (_22449_, _22448_, _05212_);
  and (_22450_, _22449_, _22447_);
  and (_22451_, _02768_, _02670_);
  or (_22452_, _22451_, _05217_);
  or (_22454_, _22452_, _22450_);
  or (_22455_, _05220_, _02230_);
  and (_22456_, _22455_, _03139_);
  and (_22457_, _22456_, _22454_);
  or (_22458_, _05225_, _02768_);
  and (_22459_, _22458_, _17972_);
  or (_22460_, _22459_, _22457_);
  or (_22461_, _22337_, _05226_);
  and (_22462_, _22461_, _22460_);
  or (_22463_, _22462_, _05229_);
  or (_22465_, _05228_, _02230_);
  and (_22466_, _22465_, _05234_);
  and (_22467_, _22466_, _22463_);
  and (_22468_, _22373_, _05233_);
  or (_22469_, _22468_, _02577_);
  or (_22470_, _22469_, _22467_);
  and (_22471_, _22470_, _22342_);
  or (_22472_, _22471_, _02575_);
  nand (_22473_, _02769_, _02575_);
  and (_22474_, _22473_, _05244_);
  and (_22476_, _22474_, _22472_);
  and (_22477_, _05243_, _02230_);
  or (_22478_, _22477_, _22476_);
  and (_22479_, _22478_, _02574_);
  or (_22480_, _05282_, \oc8051_golden_model_1.DPH [5]);
  nor (_22481_, _05283_, _02574_);
  and (_22482_, _22481_, _22480_);
  or (_22483_, _22482_, _05253_);
  or (_22484_, _22483_, _22479_);
  or (_22485_, _05252_, _02230_);
  and (_22487_, _22485_, _05291_);
  and (_22488_, _22487_, _22484_);
  or (_22489_, _22373_, _01953_);
  or (_22490_, _02230_, _02568_);
  and (_22491_, _22490_, _02567_);
  and (_22492_, _22491_, _22489_);
  or (_22493_, _22492_, _05297_);
  or (_22494_, _22493_, _22488_);
  and (_22495_, _22494_, _22341_);
  or (_22496_, _22495_, _05302_);
  or (_22498_, _05306_, _02230_);
  and (_22499_, _22498_, _05305_);
  and (_22500_, _22499_, _22496_);
  nand (_22501_, _02768_, _02656_);
  nand (_22502_, _22501_, _05311_);
  or (_22503_, _22502_, _22500_);
  or (_22504_, _05311_, _02230_);
  and (_22505_, _22504_, _05316_);
  and (_22506_, _22505_, _22503_);
  or (_22507_, _22373_, _02568_);
  or (_22509_, _02230_, _01953_);
  and (_22510_, _22509_, _05315_);
  and (_22511_, _22510_, _22507_);
  or (_22512_, _22511_, _05325_);
  or (_22513_, _22512_, _22506_);
  and (_22514_, _22513_, _22340_);
  or (_22515_, _22514_, _05329_);
  or (_22516_, _05333_, _02230_);
  and (_22517_, _22516_, _05332_);
  and (_22518_, _22517_, _22515_);
  nand (_22520_, _02768_, _02669_);
  nand (_22521_, _22520_, _05338_);
  or (_22522_, _22521_, _22518_);
  or (_22523_, _05338_, _02230_);
  and (_22524_, _22523_, _05343_);
  and (_22525_, _22524_, _22522_);
  or (_22526_, _22373_, \oc8051_golden_model_1.PSW [7]);
  or (_22527_, _02230_, _05348_);
  and (_22528_, _22527_, _05342_);
  and (_22529_, _22528_, _22526_);
  or (_22531_, _22529_, _01944_);
  or (_22532_, _22531_, _22525_);
  and (_22533_, _22532_, _22339_);
  or (_22534_, _22533_, _05355_);
  or (_22535_, _05358_, _02230_);
  and (_22536_, _22535_, _05357_);
  and (_22537_, _22536_, _22534_);
  nand (_22538_, _02768_, _02654_);
  nand (_22539_, _22538_, _05363_);
  or (_22540_, _22539_, _22537_);
  or (_22542_, _05363_, _02230_);
  and (_22543_, _22542_, _05368_);
  and (_22544_, _22543_, _22540_);
  or (_22545_, _22373_, _05348_);
  or (_22546_, _02230_, \oc8051_golden_model_1.PSW [7]);
  and (_22547_, _22546_, _05367_);
  and (_22548_, _22547_, _22545_);
  or (_22549_, _22548_, _22544_);
  and (_22550_, _22549_, _05389_);
  and (_22551_, _22337_, _05391_);
  or (_22553_, _22551_, _05393_);
  or (_22554_, _22553_, _22550_);
  or (_22555_, _05398_, _02230_);
  and (_22556_, _22555_, _05397_);
  and (_22557_, _22556_, _22554_);
  and (_22558_, _22337_, _05396_);
  or (_22559_, _22558_, _03109_);
  or (_22560_, _22559_, _22557_);
  nand (_22561_, _04480_, _03109_);
  and (_22562_, _22561_, _22560_);
  or (_22564_, _22562_, _01936_);
  or (_22565_, _02230_, _05408_);
  and (_22566_, _22565_, _03267_);
  and (_22567_, _22566_, _22564_);
  or (_22568_, _22347_, _05704_);
  or (_22569_, _05702_, _02768_);
  and (_22570_, _22569_, _02653_);
  and (_22571_, _22570_, _22568_);
  or (_22572_, _22571_, _05412_);
  or (_22573_, _22572_, _22567_);
  and (_22575_, _22573_, _22338_);
  or (_22576_, _22575_, _05720_);
  or (_22577_, _05728_, _02230_);
  and (_22578_, _22577_, _05726_);
  and (_22579_, _22578_, _22576_);
  and (_22580_, _22337_, _05724_);
  or (_22581_, _22580_, _03108_);
  or (_22582_, _22581_, _22579_);
  and (_22583_, _22582_, _22335_);
  or (_22584_, _22583_, _01899_);
  or (_22586_, _02230_, _05748_);
  and (_22587_, _22586_, _03125_);
  and (_22588_, _22587_, _22584_);
  nand (_22589_, _05702_, _02769_);
  or (_22590_, _22347_, _05702_);
  and (_22591_, _22590_, _22589_);
  and (_22592_, _22591_, _02647_);
  or (_22593_, _22592_, _05764_);
  or (_22594_, _22593_, _22588_);
  or (_22595_, _22337_, _05770_);
  and (_22597_, _22595_, _03124_);
  and (_22598_, _22597_, _22594_);
  and (_22599_, _03123_, _02230_);
  or (_22600_, _22599_, _05780_);
  or (_22601_, _22600_, _22598_);
  or (_22602_, _22337_, _05788_);
  and (_22603_, _22602_, _05786_);
  and (_22604_, _22603_, _22601_);
  nor (_22605_, _05786_, _02333_);
  or (_22606_, _22605_, _01971_);
  or (_22608_, _22606_, _22604_);
  or (_22609_, _02230_, _05802_);
  and (_22610_, _22609_, _03122_);
  and (_22611_, _22610_, _22608_);
  and (_22612_, _22591_, _02650_);
  or (_22613_, _22612_, _05826_);
  or (_22614_, _22613_, _22611_);
  or (_22615_, _22337_, _05824_);
  and (_22616_, _22615_, _03513_);
  and (_22617_, _22616_, _22614_);
  and (_22619_, _03121_, _02230_);
  or (_22620_, _22619_, _05840_);
  or (_22621_, _22620_, _22617_);
  or (_22622_, _22337_, _05848_);
  and (_22623_, _22622_, _05846_);
  and (_22624_, _22623_, _22621_);
  nand (_22625_, _02333_, _01956_);
  and (_22626_, _22625_, _18101_);
  or (_22627_, _22626_, _22624_);
  or (_22628_, _02230_, _01956_);
  and (_22630_, _22628_, _05864_);
  and (_22631_, _22630_, _22627_);
  and (_22632_, _22337_, _05862_);
  or (_22633_, _22632_, _22631_);
  or (_22634_, _22633_, _27789_);
  or (_22635_, _27788_, \oc8051_golden_model_1.PC [13]);
  and (_22636_, _22635_, _27053_);
  and (_28973_, _22636_, _22634_);
  and (_22637_, _03121_, _02217_);
  nor (_22638_, _05363_, _02217_);
  nor (_22640_, _05338_, _02217_);
  nor (_22641_, _05311_, _02217_);
  and (_22642_, _05157_, _02755_);
  and (_22643_, _03093_, _02760_);
  nor (_22644_, _22643_, _03094_);
  not (_22645_, _22644_);
  nor (_22646_, _22645_, _05157_);
  nor (_22647_, _22646_, _22642_);
  or (_22648_, _22647_, _03387_);
  and (_22649_, _04275_, _02755_);
  and (_22651_, _22644_, _04277_);
  nor (_22652_, _22651_, _22649_);
  nand (_22653_, _22652_, _02675_);
  and (_22654_, _04494_, _02755_);
  nor (_22655_, _22645_, _04494_);
  or (_22656_, _22655_, _22654_);
  nor (_22657_, _22656_, _04499_);
  nor (_22658_, _01910_, \oc8051_golden_model_1.PC [14]);
  nor (_22659_, _22658_, _01911_);
  and (_22660_, _22659_, _05009_);
  nor (_22662_, _22659_, _05004_);
  and (_22663_, _22659_, _04545_);
  or (_22664_, _04537_, _02217_);
  and (_22665_, _02549_, _02221_);
  nor (_22666_, _22665_, _02550_);
  nand (_22667_, _22666_, _04537_);
  and (_22668_, _22667_, _03406_);
  nand (_22669_, _22668_, _22664_);
  or (_22670_, _21767_, _02216_);
  or (_22671_, _22659_, _21424_);
  nand (_22673_, _04522_, _05903_);
  nor (_22674_, _04504_, \oc8051_golden_model_1.PC [14]);
  nand (_22675_, _22674_, _04521_);
  or (_22676_, _22675_, _22673_);
  and (_22677_, _22676_, _22671_);
  or (_22678_, _22677_, _03154_);
  or (_22679_, _22659_, _18144_);
  and (_22680_, _22679_, _22678_);
  or (_22681_, _22680_, _04527_);
  and (_22682_, _22681_, _22670_);
  nor (_22684_, _22682_, _03406_);
  nor (_22685_, _22684_, _04545_);
  and (_22686_, _22685_, _22669_);
  or (_22687_, _22686_, _22663_);
  nand (_22688_, _22687_, _02662_);
  nand (_22689_, _04985_, _02755_);
  or (_22690_, _22645_, _04985_);
  nand (_22691_, _22690_, _22689_);
  nand (_22692_, _22691_, _02661_);
  and (_22693_, _22692_, _18134_);
  nand (_22695_, _22693_, _22688_);
  nor (_22696_, _22659_, _18134_);
  nor (_22697_, _22696_, _21789_);
  nand (_22698_, _22697_, _22695_);
  nor (_22699_, _04995_, _02217_);
  nor (_22700_, _22699_, _05000_);
  and (_22701_, _22700_, _22698_);
  or (_22702_, _22701_, _22662_);
  nand (_22703_, _22702_, _03179_);
  and (_22704_, _03168_, _02217_);
  nor (_22706_, _22704_, _05009_);
  and (_22707_, _22706_, _22703_);
  or (_22708_, _22707_, _22660_);
  nand (_22709_, _22708_, _05013_);
  nor (_22710_, _05013_, _02217_);
  nor (_22711_, _22710_, _04498_);
  and (_22712_, _22711_, _22709_);
  or (_22713_, _22712_, _22657_);
  nand (_22714_, _22713_, _03107_);
  nand (_22715_, _22714_, _22653_);
  or (_22717_, _22715_, _02664_);
  and (_22718_, _22717_, _22648_);
  or (_22719_, _22718_, _02673_);
  nor (_22720_, _22644_, _02630_);
  and (_22721_, _02756_, _02630_);
  nor (_22722_, _22721_, _05024_);
  not (_22723_, _22722_);
  nor (_22724_, _22723_, _22720_);
  nor (_22725_, _22724_, _02598_);
  and (_22726_, _22725_, _22719_);
  nor (_22728_, _22659_, _02599_);
  or (_22729_, _22728_, _22726_);
  and (_22730_, _22729_, _05179_);
  nor (_22731_, _05179_, _02216_);
  or (_22732_, _22731_, _22730_);
  nand (_22733_, _22732_, _05186_);
  not (_22734_, _22659_);
  and (_22735_, _22734_, _05185_);
  nor (_22736_, _22735_, _05191_);
  nand (_22737_, _22736_, _22733_);
  nor (_22739_, _05190_, _02217_);
  nor (_22740_, _22739_, _05194_);
  nand (_22741_, _22740_, _22737_);
  nor (_22742_, _22659_, _05195_);
  nor (_22743_, _22742_, _05199_);
  and (_22744_, _22743_, _22741_);
  and (_22745_, _05199_, _02216_);
  or (_22746_, _22745_, _02047_);
  or (_22747_, _22746_, _22744_);
  nor (_22748_, _22659_, _01985_);
  nor (_22750_, _22748_, _05209_);
  nand (_22751_, _22750_, _22747_);
  nor (_22752_, _05208_, _02217_);
  nor (_22753_, _22752_, _02670_);
  nand (_22754_, _22753_, _22751_);
  and (_22755_, _02756_, _02670_);
  nor (_22756_, _22755_, _05217_);
  and (_22757_, _22756_, _22754_);
  and (_22758_, _05217_, _02216_);
  or (_22759_, _22758_, _02024_);
  or (_22761_, _22759_, _22757_);
  and (_22762_, _02756_, _02024_);
  nor (_22763_, _22762_, _05225_);
  nand (_22764_, _22763_, _22761_);
  and (_22765_, _22659_, _05225_);
  nor (_22766_, _22765_, _05229_);
  nand (_22767_, _22766_, _22764_);
  nor (_22768_, _05228_, _02216_);
  nor (_22769_, _22768_, _05233_);
  and (_22770_, _22769_, _22767_);
  and (_22772_, _22666_, _05233_);
  nor (_22773_, _22772_, _22770_);
  or (_22774_, _22773_, _02577_);
  nand (_22775_, _02577_, _02216_);
  and (_22776_, _22775_, _05245_);
  nand (_22777_, _22776_, _22774_);
  and (_22778_, _02756_, _02575_);
  nor (_22779_, _22778_, _05243_);
  nand (_22780_, _22779_, _22777_);
  and (_22781_, _05243_, _02216_);
  nor (_22783_, _22781_, _02573_);
  nand (_22784_, _22783_, _22780_);
  nor (_22785_, _05283_, \oc8051_golden_model_1.DPH [6]);
  nor (_22786_, _22785_, _05284_);
  nor (_22787_, _22786_, _02574_);
  nor (_22788_, _22787_, _05253_);
  and (_22789_, _22788_, _22784_);
  nor (_22790_, _05252_, _02217_);
  or (_22791_, _22790_, _22789_);
  nand (_22792_, _22791_, _05291_);
  and (_22794_, _02216_, _01953_);
  and (_22795_, _22666_, _02568_);
  or (_22796_, _22795_, _22794_);
  and (_22797_, _22796_, _02567_);
  nor (_22798_, _22797_, _05297_);
  nand (_22799_, _22798_, _22792_);
  nor (_22800_, _22659_, _05298_);
  nor (_22801_, _22800_, _05302_);
  nand (_22802_, _22801_, _22799_);
  and (_22803_, _05302_, _02216_);
  nor (_22805_, _22803_, _02656_);
  nand (_22806_, _22805_, _22802_);
  and (_22807_, _02756_, _02656_);
  nor (_22808_, _22807_, _05312_);
  and (_22809_, _22808_, _22806_);
  or (_22810_, _22809_, _22641_);
  nand (_22811_, _22810_, _05316_);
  and (_22812_, _02216_, _02568_);
  and (_22813_, _22666_, _01953_);
  or (_22814_, _22813_, _22812_);
  and (_22816_, _22814_, _05315_);
  nor (_22817_, _22816_, _05325_);
  nand (_22818_, _22817_, _22811_);
  nor (_22819_, _22659_, _05326_);
  nor (_22820_, _22819_, _05329_);
  nand (_22821_, _22820_, _22818_);
  and (_22822_, _05329_, _02216_);
  nor (_22823_, _22822_, _02669_);
  nand (_22824_, _22823_, _22821_);
  and (_22825_, _02756_, _02669_);
  nor (_22827_, _22825_, _05339_);
  and (_22828_, _22827_, _22824_);
  or (_22829_, _22828_, _22640_);
  nand (_22830_, _22829_, _05343_);
  nor (_22831_, _22666_, \oc8051_golden_model_1.PSW [7]);
  nor (_22832_, _02216_, _05348_);
  nor (_22833_, _22832_, _05343_);
  not (_22834_, _22833_);
  nor (_22835_, _22834_, _22831_);
  nor (_22836_, _22835_, _01944_);
  nand (_22838_, _22836_, _22830_);
  nor (_22839_, _22659_, _01945_);
  nor (_22840_, _22839_, _05355_);
  nand (_22841_, _22840_, _22838_);
  and (_22842_, _05355_, _02216_);
  nor (_22843_, _22842_, _02654_);
  nand (_22844_, _22843_, _22841_);
  and (_22845_, _02756_, _02654_);
  nor (_22846_, _22845_, _05364_);
  and (_22847_, _22846_, _22844_);
  or (_22849_, _22847_, _22638_);
  nand (_22850_, _22849_, _05368_);
  nor (_22851_, _22666_, _05348_);
  nor (_22852_, _02216_, \oc8051_golden_model_1.PSW [7]);
  nor (_22853_, _22852_, _05368_);
  not (_22854_, _22853_);
  nor (_22855_, _22854_, _22851_);
  nor (_22856_, _22855_, _05391_);
  nand (_22857_, _22856_, _22850_);
  nor (_22858_, _22659_, _05389_);
  nor (_22860_, _22858_, _05393_);
  and (_22861_, _22860_, _22857_);
  and (_22862_, _05393_, _02216_);
  or (_22863_, _22862_, _22861_);
  and (_22864_, _22863_, _05397_);
  and (_22865_, _22659_, _05396_);
  or (_22866_, _22865_, _22864_);
  and (_22867_, _22866_, _06612_);
  nor (_22868_, _04373_, _06612_);
  or (_22869_, _22868_, _01936_);
  or (_22871_, _22869_, _22867_);
  and (_22872_, _02217_, _01936_);
  nor (_22873_, _22872_, _02653_);
  nand (_22874_, _22873_, _22871_);
  and (_22875_, _22645_, _05702_);
  nor (_22876_, _05702_, _02755_);
  or (_22877_, _22876_, _03267_);
  nor (_22878_, _22877_, _22875_);
  nor (_22879_, _22878_, _05412_);
  nand (_22880_, _22879_, _22874_);
  nor (_22882_, _22659_, _01930_);
  nor (_22883_, _22882_, _05720_);
  and (_22884_, _22883_, _22880_);
  and (_22885_, _05720_, _02216_);
  or (_22886_, _22885_, _22884_);
  and (_22887_, _22886_, _05726_);
  and (_22888_, _22659_, _05724_);
  or (_22889_, _22888_, _03108_);
  or (_22890_, _22889_, _22887_);
  and (_22891_, _04373_, _03108_);
  nor (_22893_, _22891_, _01899_);
  and (_22894_, _22893_, _22890_);
  and (_22895_, _02216_, _01899_);
  or (_22896_, _22895_, _02647_);
  nor (_22897_, _22896_, _22894_);
  and (_22898_, _05702_, _02756_);
  nor (_22899_, _22644_, _05702_);
  nor (_22900_, _22899_, _22898_);
  nor (_22901_, _22900_, _03125_);
  or (_22902_, _22901_, _22897_);
  and (_22904_, _22902_, _05770_);
  nor (_22905_, _22659_, _05770_);
  or (_22906_, _22905_, _22904_);
  nand (_22907_, _22906_, _03124_);
  and (_22908_, _03123_, _02217_);
  nor (_22909_, _22908_, _05780_);
  nand (_22910_, _22909_, _22907_);
  and (_22911_, _22659_, _05780_);
  nor (_22912_, _22911_, _02646_);
  nand (_22913_, _22912_, _22910_);
  and (_22915_, _02646_, _02295_);
  nor (_22916_, _22915_, _01971_);
  nand (_22917_, _22916_, _22913_);
  and (_22918_, _02216_, _01971_);
  nor (_22919_, _22918_, _02650_);
  nand (_22920_, _22919_, _22917_);
  nor (_22921_, _22900_, _03122_);
  nor (_22922_, _22921_, _05826_);
  nand (_22923_, _22922_, _22920_);
  nor (_22924_, _22734_, _05824_);
  nor (_22926_, _22924_, _03121_);
  and (_22927_, _22926_, _22923_);
  or (_22928_, _22927_, _22637_);
  nand (_22929_, _22928_, _05848_);
  nor (_22930_, _22659_, _05848_);
  nor (_22931_, _22930_, _02649_);
  and (_22932_, _22931_, _22929_);
  and (_22933_, _02295_, _01956_);
  nor (_22934_, _22933_, _18100_);
  or (_22935_, _22934_, _22932_);
  and (_22937_, _02217_, _01955_);
  nor (_22938_, _22937_, _05862_);
  and (_22939_, _22938_, _22935_);
  and (_22940_, _22659_, _05862_);
  or (_22941_, _22940_, _22939_);
  or (_22942_, _22941_, _27789_);
  or (_22943_, _27788_, \oc8051_golden_model_1.PC [14]);
  and (_22944_, _22943_, _27053_);
  and (_28974_, _22944_, _22942_);
  and (_22945_, _27789_, \oc8051_golden_model_1.P0INREG [0]);
  or (_22947_, _22945_, _28129_);
  and (_28975_, _22947_, _27053_);
  and (_22948_, _27789_, \oc8051_golden_model_1.P0INREG [1]);
  or (_22949_, _22948_, _28111_);
  and (_28976_, _22949_, _27053_);
  and (_22950_, _27789_, \oc8051_golden_model_1.P0INREG [2]);
  or (_22951_, _22950_, _28085_);
  and (_28979_, _22951_, _27053_);
  and (_22952_, _27789_, \oc8051_golden_model_1.P0INREG [3]);
  or (_22953_, _22952_, _28140_);
  and (_28980_, _22953_, _27053_);
  and (_22955_, _27789_, \oc8051_golden_model_1.P0INREG [4]);
  or (_22956_, _22955_, _28121_);
  and (_28981_, _22956_, _27053_);
  and (_22957_, _27789_, \oc8051_golden_model_1.P0INREG [5]);
  or (_22958_, _22957_, _28103_);
  and (_28982_, _22958_, _27053_);
  and (_22959_, _27789_, \oc8051_golden_model_1.P0INREG [6]);
  or (_22960_, _22959_, _28093_);
  and (_28983_, _22960_, _27053_);
  and (_22962_, _27789_, \oc8051_golden_model_1.P1INREG [0]);
  or (_22963_, _22962_, _27847_);
  and (_28986_, _22963_, _27053_);
  and (_22964_, _27789_, \oc8051_golden_model_1.P1INREG [1]);
  or (_22965_, _22964_, _27809_);
  and (_28987_, _22965_, _27053_);
  and (_22966_, _27789_, \oc8051_golden_model_1.P1INREG [2]);
  or (_22967_, _22966_, _27799_);
  and (_28988_, _22967_, _27053_);
  and (_22968_, _27789_, \oc8051_golden_model_1.P1INREG [3]);
  or (_22970_, _22968_, _27837_);
  and (_28989_, _22970_, _27053_);
  and (_22971_, _27789_, \oc8051_golden_model_1.P1INREG [4]);
  or (_22972_, _22971_, _27856_);
  and (_28990_, _22972_, _27053_);
  and (_22973_, _27789_, \oc8051_golden_model_1.P1INREG [5]);
  or (_22974_, _22973_, _27818_);
  and (_28991_, _22974_, _27053_);
  and (_22975_, _27789_, \oc8051_golden_model_1.P1INREG [6]);
  or (_22976_, _22975_, _27791_);
  and (_28992_, _22976_, _27053_);
  and (_22978_, _27789_, \oc8051_golden_model_1.P2INREG [0]);
  or (_22979_, _22978_, _28062_);
  and (_28993_, _22979_, _27053_);
  and (_22980_, _27789_, \oc8051_golden_model_1.P2INREG [1]);
  or (_22981_, _22980_, _27998_);
  and (_28994_, _22981_, _27053_);
  and (_22982_, _27789_, \oc8051_golden_model_1.P2INREG [2]);
  or (_22983_, _22982_, _27985_);
  and (_28995_, _22983_, _27053_);
  and (_22985_, _27789_, \oc8051_golden_model_1.P2INREG [3]);
  or (_22986_, _22985_, _28050_);
  and (_28996_, _22986_, _27053_);
  and (_22987_, _27789_, \oc8051_golden_model_1.P2INREG [4]);
  or (_22988_, _22987_, _28070_);
  and (_28999_, _22988_, _27053_);
  and (_22989_, _27789_, \oc8051_golden_model_1.P2INREG [5]);
  or (_22990_, _22989_, _28014_);
  and (_29000_, _22990_, _27053_);
  and (_22991_, _27789_, \oc8051_golden_model_1.P2INREG [6]);
  or (_22993_, _22991_, _27977_);
  and (_29001_, _22993_, _27053_);
  and (_22994_, _27789_, \oc8051_golden_model_1.P3INREG [0]);
  or (_22995_, _22994_, _28171_);
  and (_29004_, _22995_, _27053_);
  and (_22996_, _27789_, \oc8051_golden_model_1.P3INREG [1]);
  or (_22997_, _22996_, _28228_);
  and (_29005_, _22997_, _27053_);
  and (_22998_, _27789_, \oc8051_golden_model_1.P3INREG [2]);
  or (_22999_, _22998_, _28210_);
  and (_29006_, _22999_, _27053_);
  and (_23001_, _27789_, \oc8051_golden_model_1.P3INREG [3]);
  or (_23002_, _23001_, _28190_);
  and (_29007_, _23002_, _27053_);
  and (_23003_, _27789_, \oc8051_golden_model_1.P3INREG [4]);
  or (_23004_, _23003_, _28163_);
  and (_29008_, _23004_, _27053_);
  and (_23005_, _27789_, \oc8051_golden_model_1.P3INREG [5]);
  or (_23006_, _23005_, _28220_);
  and (_29009_, _23006_, _27053_);
  and (_23008_, _27789_, \oc8051_golden_model_1.P3INREG [6]);
  or (_23009_, _23008_, _28201_);
  and (_29010_, _23009_, _27053_);
  nor (_00006_[6], _28203_, rst);
  nor (_00006_[5], _28221_, rst);
  nor (_00006_[4], _28164_, rst);
  nor (_00006_[3], _28191_, rst);
  nor (_00006_[2], _28211_, rst);
  nor (_00006_[1], _28229_, rst);
  nor (_00006_[0], _28172_, rst);
  nor (_00005_[6], _27978_, rst);
  nor (_00005_[5], _28016_, rst);
  nor (_00005_[4], _28071_, rst);
  nor (_00005_[3], _28052_, rst);
  nor (_00005_[2], _27986_, rst);
  nor (_00005_[1], _28000_, rst);
  nor (_00005_[0], _28063_, rst);
  nor (_00004_[6], _27792_, rst);
  nor (_00004_[5], _27819_, rst);
  nor (_00004_[4], _27857_, rst);
  nor (_00004_[3], _27838_, rst);
  nor (_00004_[2], _27800_, rst);
  nor (_00004_[1], _27810_, rst);
  nor (_00004_[0], _27848_, rst);
  nor (_00002_[6], _28094_, rst);
  nor (_00002_[5], _28104_, rst);
  nor (_00002_[4], _28122_, rst);
  nor (_00002_[3], _28141_, rst);
  nor (_00002_[2], _28086_, rst);
  nor (_00002_[1], _28112_, rst);
  nor (_00002_[0], _28130_, rst);
  nor (_00004_[7], _27830_, rst);
  nor (_00005_[7], _28036_, rst);
  nor (_00006_[7], _28183_, rst);
  nor (_23013_, _11298_, _10582_);
  nor (_23014_, _14684_, _13201_);
  and (_23015_, _23014_, _23013_);
  nor (_23016_, _06857_, _06599_);
  nor (_23017_, _07245_, _07137_);
  and (_23018_, _23017_, _23016_);
  or (_23020_, _13513_, _11610_);
  nor (_23021_, _23020_, _14996_);
  and (_23022_, _12896_, _10993_);
  nand (_23023_, _23022_, _14379_);
  nor (_23024_, _23023_, _06135_);
  nor (_23025_, _06300_, _06217_);
  and (_23026_, _23025_, _23024_);
  nor (_23027_, _16572_, _16253_);
  nor (_23028_, _16803_, _16650_);
  and (_23029_, _23028_, _23027_);
  nor (_23031_, _15699_, _15545_);
  nor (_23032_, _16100_, _15859_);
  and (_23033_, _23032_, _23031_);
  and (_23034_, _23033_, _23029_);
  or (_23035_, _17402_, _17234_);
  or (_23036_, _23035_, _17839_);
  nor (_23037_, _23036_, _12061_);
  and (_23038_, _23037_, _23034_);
  nor (_23039_, _16410_, _16332_);
  nor (_23040_, _15779_, _15225_);
  and (_23042_, _23040_, _23039_);
  nor (_23043_, _16175_, _15621_);
  nor (_23044_, _17315_, _16725_);
  and (_23045_, _23044_, _23043_);
  nor (_23046_, \oc8051_golden_model_1.IE [1], \oc8051_golden_model_1.IE [0]);
  nor (_23047_, \oc8051_golden_model_1.IE [3], \oc8051_golden_model_1.IE [2]);
  and (_23048_, _23047_, _23046_);
  nor (_23049_, \oc8051_golden_model_1.IP [4], \oc8051_golden_model_1.IP [3]);
  nor (_23050_, \oc8051_golden_model_1.IP [6], \oc8051_golden_model_1.IP [5]);
  and (_23051_, _23050_, _23049_);
  and (_23053_, _23051_, _23048_);
  nor (_23054_, \oc8051_golden_model_1.SBUF [3], \oc8051_golden_model_1.SBUF [2]);
  nor (_23055_, \oc8051_golden_model_1.SBUF [4], \oc8051_golden_model_1.SBUF [1]);
  and (_23056_, _23055_, _23054_);
  nor (_23057_, \oc8051_golden_model_1.IE [5], \oc8051_golden_model_1.IE [4]);
  nor (_23058_, \oc8051_golden_model_1.SBUF [0], \oc8051_golden_model_1.IE [6]);
  and (_23059_, _23058_, _23057_);
  and (_23060_, _23059_, _23056_);
  and (_23061_, _23060_, _23053_);
  nor (_23062_, \oc8051_golden_model_1.IE [7], \oc8051_golden_model_1.IP [7]);
  nor (_23064_, \oc8051_golden_model_1.SCON [7], \oc8051_golden_model_1.SBUF [7]);
  nor (_23065_, \oc8051_golden_model_1.TL1 [7], \oc8051_golden_model_1.TH1 [7]);
  and (_23066_, _23065_, _23064_);
  and (_23067_, _23066_, _23062_);
  nor (_23068_, \oc8051_golden_model_1.IP [1], \oc8051_golden_model_1.IP [0]);
  nor (_23069_, \oc8051_golden_model_1.IP [2], \oc8051_golden_model_1.PCON [7]);
  and (_23070_, _23069_, _23068_);
  nor (_23071_, \oc8051_golden_model_1.TL0 [7], \oc8051_golden_model_1.TH0 [7]);
  nor (_23072_, \oc8051_golden_model_1.TCON [7], \oc8051_golden_model_1.TMOD [7]);
  and (_23073_, _23072_, _23071_);
  and (_23075_, _23073_, _23070_);
  and (_23076_, _23075_, _23067_);
  and (_23077_, _23076_, _23061_);
  nor (_23078_, \oc8051_golden_model_1.TL1 [1], \oc8051_golden_model_1.TL1 [0]);
  nor (_23079_, \oc8051_golden_model_1.TL1 [3], \oc8051_golden_model_1.TL1 [2]);
  and (_23080_, _23079_, _23078_);
  nor (_23081_, \oc8051_golden_model_1.TL1 [5], \oc8051_golden_model_1.TL1 [4]);
  nor (_23082_, \oc8051_golden_model_1.TH0 [0], \oc8051_golden_model_1.TL1 [6]);
  and (_23083_, _23082_, _23081_);
  and (_23084_, _23083_, _23080_);
  nor (_23086_, \oc8051_golden_model_1.TL0 [1], \oc8051_golden_model_1.TL0 [0]);
  nor (_23087_, \oc8051_golden_model_1.TH0 [6], \oc8051_golden_model_1.TH0 [5]);
  and (_23088_, _23087_, _23086_);
  nor (_23089_, \oc8051_golden_model_1.TH0 [2], \oc8051_golden_model_1.TH0 [1]);
  nor (_23090_, \oc8051_golden_model_1.TH0 [4], \oc8051_golden_model_1.TH0 [3]);
  and (_23091_, _23090_, _23089_);
  and (_23092_, _23091_, _23088_);
  and (_23093_, _23092_, _23084_);
  nor (_23094_, \oc8051_golden_model_1.SCON [3], \oc8051_golden_model_1.SCON [2]);
  nor (_23095_, \oc8051_golden_model_1.SCON [5], \oc8051_golden_model_1.SCON [4]);
  and (_23097_, _23095_, _23094_);
  nor (_23098_, \oc8051_golden_model_1.SCON [1], \oc8051_golden_model_1.SCON [0]);
  nor (_23099_, \oc8051_golden_model_1.SBUF [6], \oc8051_golden_model_1.SBUF [5]);
  and (_23100_, _23099_, _23098_);
  and (_23101_, _23100_, _23097_);
  nor (_23102_, \oc8051_golden_model_1.TH1 [5], \oc8051_golden_model_1.TH1 [4]);
  nor (_23103_, \oc8051_golden_model_1.TH1 [6], \oc8051_golden_model_1.TH1 [3]);
  and (_23104_, _23103_, _23102_);
  nor (_23105_, \oc8051_golden_model_1.TH1 [0], \oc8051_golden_model_1.SCON [6]);
  nor (_23106_, \oc8051_golden_model_1.TH1 [2], \oc8051_golden_model_1.TH1 [1]);
  and (_23108_, _23106_, _23105_);
  and (_23109_, _23108_, _23104_);
  and (_23110_, _23109_, _23101_);
  and (_23111_, _23110_, _23093_);
  nor (_23112_, \oc8051_golden_model_1.PCON [6], \oc8051_golden_model_1.PCON [5]);
  and (_23113_, _23112_, regs_always_zero);
  nor (_23114_, \oc8051_golden_model_1.PCON [3], \oc8051_golden_model_1.PCON [2]);
  nor (_23115_, \oc8051_golden_model_1.PCON [4], \oc8051_golden_model_1.PCON [1]);
  and (_23116_, _23115_, _23114_);
  nor (_23117_, \oc8051_golden_model_1.TCON [5], \oc8051_golden_model_1.TCON [4]);
  nor (_23119_, \oc8051_golden_model_1.PCON [0], \oc8051_golden_model_1.TCON [6]);
  and (_23120_, _23119_, _23117_);
  and (_23121_, _23120_, _23116_);
  and (_23122_, _23121_, _23113_);
  nor (_23123_, \oc8051_golden_model_1.TMOD [1], \oc8051_golden_model_1.TMOD [0]);
  nor (_23124_, \oc8051_golden_model_1.TMOD [2], \oc8051_golden_model_1.TL0 [6]);
  and (_23125_, _23124_, _23123_);
  nor (_23126_, \oc8051_golden_model_1.TL0 [3], \oc8051_golden_model_1.TL0 [2]);
  nor (_23127_, \oc8051_golden_model_1.TL0 [5], \oc8051_golden_model_1.TL0 [4]);
  and (_23128_, _23127_, _23126_);
  and (_23130_, _23128_, _23125_);
  and (_23131_, \oc8051_golden_model_1.TCON [1], _14284_);
  nor (_23132_, \oc8051_golden_model_1.TCON [3], \oc8051_golden_model_1.TCON [2]);
  and (_23133_, _23132_, _23131_);
  nor (_23134_, \oc8051_golden_model_1.TMOD [4], \oc8051_golden_model_1.TMOD [3]);
  nor (_23135_, \oc8051_golden_model_1.TMOD [6], \oc8051_golden_model_1.TMOD [5]);
  and (_23136_, _23135_, _23134_);
  and (_23137_, _23136_, _23133_);
  and (_23138_, _23137_, _23130_);
  and (_23139_, _23138_, _23122_);
  and (_23141_, _23139_, _23111_);
  nand (_23142_, _23141_, _23077_);
  nor (_23143_, _23142_, _11742_);
  nor (_23144_, _15068_, _12321_);
  and (_23145_, _23144_, _23143_);
  and (_23146_, _23145_, _23045_);
  nor (_23147_, _12478_, _11900_);
  and (_23148_, _23147_, _23146_);
  and (_23149_, _23148_, _23042_);
  nor (_23150_, _16969_, _16884_);
  nor (_23152_, _17575_, _17489_);
  and (_23153_, _23152_, _23150_);
  and (_23154_, _23153_, _10274_);
  and (_23155_, _23154_, _23149_);
  nor (_23156_, _12798_, _12558_);
  nor (_23157_, _15305_, _15146_);
  and (_23158_, _23157_, _23156_);
  nor (_23159_, _11980_, _11820_);
  nor (_23160_, _12399_, _12247_);
  and (_23161_, _23160_, _23159_);
  and (_23163_, _23161_, _23158_);
  and (_23164_, _23163_, _23155_);
  and (_23165_, _23164_, _23038_);
  and (_23166_, _23165_, _23026_);
  nor (_23167_, _06470_, _06385_);
  nor (_23168_, _07022_, _06940_);
  and (_23169_, _23168_, _23167_);
  not (_23170_, _12995_);
  and (_23171_, _14478_, _23170_);
  nor (_23172_, _11092_, _10376_);
  and (_23174_, _23172_, _23171_);
  and (_23175_, _23174_, _23169_);
  and (_23176_, _23175_, _23166_);
  nor (_23177_, _17148_, _17059_);
  nor (_23178_, _17752_, _17663_);
  and (_23179_, _23178_, _23177_);
  nor (_23180_, _15940_, _15467_);
  nor (_23181_, _16491_, _16021_);
  and (_23182_, _23181_, _23180_);
  nor (_23183_, _12638_, _12156_);
  nor (_23185_, _15385_, _12720_);
  and (_23186_, _23185_, _23183_);
  and (_23187_, _23186_, _23182_);
  nand (_23188_, _23187_, _23179_);
  nor (_23189_, _23188_, _10894_);
  and (_23190_, _23189_, _23176_);
  and (_23191_, _23190_, _23021_);
  and (_23192_, _23191_, _23018_);
  and (_23193_, _23192_, _23015_);
  nor (_23194_, _14893_, _14788_);
  nor (_23196_, _14581_, _13410_);
  and (_23197_, _23196_, _23194_);
  nor (_23198_, _11507_, _11402_);
  nor (_23199_, _13305_, _13098_);
  and (_23200_, _23199_, _23198_);
  nor (_23201_, _10686_, _10479_);
  nor (_23202_, _11195_, _10791_);
  and (_23203_, _23202_, _23201_);
  and (_23204_, _23203_, _23200_);
  and (_23205_, _23204_, _23197_);
  and (_23207_, _23205_, _23193_);
  or (_00009_, _23207_, rst);
  and (_23208_, ABINPUT008[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nor (_23209_, ABINPUT008[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_23210_, _23209_, _23208_);
  nand (_23211_, ABINPUT008[2], _24460_);
  or (_23212_, ABINPUT008[6], _24505_);
  and (_23213_, _23212_, _23211_);
  and (_23214_, _23213_, _23210_);
  and (_23215_, ABINPUT008[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor (_23217_, ABINPUT008[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_23218_, _23217_, _23215_);
  or (_23219_, ABINPUT008[2], _24460_);
  and (_23220_, _23219_, _27053_);
  and (_23221_, _23220_, _23218_);
  and (_23222_, _23221_, _23214_);
  nand (_23223_, ABINPUT008[6], _24505_);
  or (_23224_, ABINPUT008[4], _25809_);
  or (_23225_, ABINPUT008[7], _24435_);
  and (_23226_, _23225_, _23224_);
  and (_23228_, _23226_, _23223_);
  and (_23229_, ABINPUT008[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_23230_, ABINPUT008[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_23231_, _23230_, _23229_);
  nand (_23232_, ABINPUT008[4], _25809_);
  nand (_23233_, ABINPUT008[7], _24435_);
  and (_23234_, _23233_, _23232_);
  and (_23235_, _23234_, _23231_);
  and (_23236_, _23235_, _23228_);
  and (_00007_, _23236_, _23222_);
  nand (_23238_, _14280_, _24332_);
  or (_23239_, _14280_, _24332_);
  and (_23240_, _23239_, _23238_);
  or (_23241_, _13811_, _24308_);
  nand (_23242_, _13811_, _24308_);
  and (_23243_, _23242_, _23241_);
  or (_23244_, _13921_, _25652_);
  nand (_23245_, _13921_, _25652_);
  and (_23246_, _23245_, _23244_);
  and (_23247_, _23246_, _23243_);
  nand (_23249_, _14041_, _25833_);
  or (_23250_, _14041_, _25833_);
  or (_23251_, _13588_, _24296_);
  nand (_23252_, _13588_, _24296_);
  and (_23253_, _23252_, _23251_);
  and (_23254_, _23253_, _27053_);
  or (_23255_, _13700_, _25884_);
  nand (_23256_, _13700_, _25884_);
  and (_23257_, _23256_, _23255_);
  and (_23258_, _23257_, _23254_);
  and (_23260_, _23258_, _23250_);
  and (_23261_, _23260_, _23249_);
  and (_23262_, _23261_, _23247_);
  not (_23263_, _24326_);
  nand (_23264_, _14161_, _23263_);
  or (_23265_, _06749_, _25615_);
  and (_23266_, _23265_, _23264_);
  or (_23267_, _14161_, _23263_);
  nand (_23268_, _06749_, _25615_);
  and (_23269_, _23268_, _23267_);
  and (_23271_, _23269_, _23266_);
  and (_23272_, _23271_, _23262_);
  and (_00008_, _23272_, _23240_);
  nand (_23273_, _18534_, _29665_);
  or (_23274_, _18534_, _29665_);
  or (_23275_, _20357_, _29685_);
  or (_23276_, _20725_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_23277_, _20725_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_23278_, _23277_, _23276_);
  and (_23279_, _23278_, _23275_);
  nand (_23281_, _19632_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_23282_, _19632_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_23283_, _20000_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_23284_, _21059_, _29693_);
  or (_23285_, _21059_, _29693_);
  and (_23286_, _21391_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_23287_, _21391_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_23288_, _05874_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_23289_, _05874_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_23290_, _23289_, _23288_);
  nand (_23292_, _22941_, _29712_);
  or (_23293_, _22941_, _29712_);
  nand (_23294_, _23293_, _23292_);
  nor (_23295_, _23294_, _23290_);
  or (_23296_, _21709_, _29178_);
  nand (_23297_, _21709_, _29178_);
  nand (_23298_, _23297_, _23296_);
  nor (_23299_, _22633_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_23300_, _22633_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_23301_, _23300_, _23299_);
  not (_23303_, _23301_);
  and (_23304_, _22018_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_23305_, _22018_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_23306_, _23305_, _23304_);
  nor (_23307_, _18111_, _29661_);
  and (_23308_, _18111_, _29661_);
  nor (_23309_, _23308_, _23307_);
  nor (_23310_, _23309_, _23306_);
  and (_23311_, _23310_, _23303_);
  and (_23312_, _23311_, _23298_);
  and (_23314_, _23312_, _23295_);
  nand (_23315_, _22330_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_23316_, _22330_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_23317_, _23316_, _23315_);
  and (_23318_, _23317_, _23314_);
  nand (_23319_, _23318_, _23287_);
  nor (_23320_, _23319_, _23286_);
  nand (_23321_, _23320_, _23285_);
  nor (_23322_, _23321_, _23284_);
  and (_23323_, _23322_, _23283_);
  and (_23325_, _23323_, _23282_);
  and (_23326_, _23325_, _23281_);
  nand (_23327_, _20357_, _29685_);
  nand (_23328_, _19270_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_23329_, _20000_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_23330_, _19270_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_23331_, _23330_, _23329_);
  and (_23332_, _23331_, _23328_);
  and (_23333_, _23332_, _23327_);
  and (_23334_, _23333_, _23326_);
  and (_23336_, _23334_, _23279_);
  nand (_23337_, _18910_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_23338_, _18910_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_23339_, _23338_, _23337_);
  and (_23340_, _23339_, _23336_);
  and (_23341_, _23340_, _23274_);
  nand (_23342_, _23341_, _23273_);
  nand (_23343_, _23207_, _00001_);
  nor (_00003_, _23343_, _23342_);
  and (_23344_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor (_23346_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_23347_, _23346_, _23344_);
  and (_23348_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor (_23349_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_23350_, _23349_, _23348_);
  and (_23351_, _23350_, _23347_);
  or (_23352_, \oc8051_golden_model_1.P3 [2], _25008_);
  or (_23353_, _11647_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_23354_, _23353_, _23352_);
  or (_23355_, \oc8051_golden_model_1.P3 [0], _24981_);
  or (_23357_, _11645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_23358_, _23357_, _23355_);
  and (_23359_, _23358_, _23354_);
  and (_23360_, _23359_, _23351_);
  or (_23361_, _11631_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_23362_, \oc8051_golden_model_1.P1 [6], _24869_);
  and (_23363_, _23362_, _23361_);
  or (_23364_, _11628_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_23365_, \oc8051_golden_model_1.P1 [4], _24841_);
  and (_23366_, _23365_, _23364_);
  and (_23368_, _23366_, _23363_);
  and (_23369_, \oc8051_golden_model_1.P1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_23370_, \oc8051_golden_model_1.P1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_23371_, _23370_, _23369_);
  and (_23372_, \oc8051_golden_model_1.P2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_23373_, \oc8051_golden_model_1.P2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_23374_, _23373_, _23372_);
  and (_23375_, _23374_, _23371_);
  and (_23376_, _23375_, _23368_);
  and (_23377_, _23376_, _23360_);
  and (_23379_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_23380_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_23381_, _23380_, _23379_);
  and (_23382_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nor (_23383_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_23384_, _23383_, _23382_);
  and (_23385_, _23384_, _23381_);
  or (_23386_, \oc8051_golden_model_1.P3 [7], _24678_);
  or (_23387_, _11656_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_23388_, _07027_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_23390_, _23388_, _23387_);
  and (_23391_, _23390_, _23386_);
  or (_23392_, \oc8051_golden_model_1.P3 [6], _25064_);
  or (_23393_, _11653_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_23394_, _23393_, _23392_);
  or (_23395_, \oc8051_golden_model_1.P3 [4], _25036_);
  or (_23396_, _11650_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_23397_, _23396_, _23395_);
  and (_23398_, _23397_, _23394_);
  and (_23399_, _23398_, _23391_);
  and (_23401_, _23399_, _23385_);
  or (_23402_, \oc8051_golden_model_1.P2 [6], _24966_);
  or (_23403_, _11642_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_23404_, _23403_, _23402_);
  or (_23405_, _11639_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_23406_, \oc8051_golden_model_1.P2 [4], _24938_);
  and (_23407_, _23406_, _23405_);
  and (_23408_, _23407_, _23404_);
  and (_23409_, \oc8051_golden_model_1.P2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_23410_, \oc8051_golden_model_1.P2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_23412_, _23410_, _23409_);
  and (_23413_, \oc8051_golden_model_1.P3 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_23414_, \oc8051_golden_model_1.P3 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_23415_, _23414_, _23413_);
  and (_23416_, _23415_, _23412_);
  and (_23417_, _23416_, _23408_);
  and (_23418_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_23419_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_23420_, _23419_, _23418_);
  and (_23421_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_23423_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_23424_, _23423_, _23421_);
  and (_23425_, _23424_, _23420_);
  or (_23426_, \oc8051_golden_model_1.P2 [2], _24911_);
  or (_23427_, _11636_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_23428_, _23427_, _23426_);
  or (_23429_, _11634_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_23430_, \oc8051_golden_model_1.P2 [0], _24883_);
  and (_23431_, _23430_, _23429_);
  and (_23432_, _23431_, _23428_);
  and (_23434_, _23432_, _23425_);
  and (_23435_, _23434_, _23417_);
  and (_23436_, _23435_, _23401_);
  and (_23437_, _23436_, _23377_);
  nand (_23438_, ABINPUT009[84], _26383_);
  or (_23439_, ABINPUT009[86], _26393_);
  and (_23440_, _23439_, _23438_);
  or (_23441_, ABINPUT009[84], _26383_);
  nand (_23442_, ABINPUT009[82], _26378_);
  and (_23443_, _23442_, _23441_);
  and (_23445_, _23443_, _23440_);
  and (_23446_, ABINPUT009[87], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nor (_23447_, ABINPUT009[87], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_23448_, _23447_, _23446_);
  and (_23449_, ABINPUT009[89], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_23450_, ABINPUT009[89], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_23451_, _23450_, _23449_);
  and (_23452_, _23451_, _23448_);
  and (_23453_, _23452_, _23445_);
  and (_23454_, ABINPUT009[75], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_23456_, ABINPUT009[75], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_23457_, _23456_, _23454_);
  and (_23458_, ABINPUT009[77], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_23459_, ABINPUT009[77], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_23460_, _23459_, _23458_);
  and (_23461_, _23460_, _23457_);
  nand (_23462_, ABINPUT009[78], _26366_);
  or (_23463_, ABINPUT009[80], _26371_);
  and (_23464_, _23463_, _23462_);
  or (_23465_, ABINPUT009[82], _26378_);
  nand (_23467_, ABINPUT009[80], _26371_);
  and (_23468_, _23467_, _23465_);
  and (_23469_, _23468_, _23464_);
  and (_23470_, _23469_, _23461_);
  and (_23471_, _23470_, _23453_);
  and (_23472_, ABINPUT009[101], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_23473_, ABINPUT009[101], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_23474_, _23473_, _23472_);
  nand (_23475_, ABINPUT009[100], _26456_);
  or (_23476_, ABINPUT009[102], _26463_);
  and (_23478_, _23476_, _23475_);
  and (_23479_, _23478_, _23474_);
  and (_23480_, ABINPUT009[99], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_23481_, ABINPUT009[99], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_23482_, _23481_, _23480_);
  or (_23483_, ABINPUT009[100], _26456_);
  nand (_23484_, ABINPUT009[98], _26450_);
  and (_23485_, _23484_, _23483_);
  and (_23486_, _23485_, _23482_);
  and (_23487_, _23486_, _23479_);
  nor (_23489_, ABINPUT009[95], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_23490_, ABINPUT009[95], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_23491_, _23490_, _23489_);
  nor (_23492_, ABINPUT009[97], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and (_23493_, ABINPUT009[97], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_23494_, _23493_, _23492_);
  and (_23495_, _23494_, _23491_);
  nand (_23496_, ABINPUT009[92], _26433_);
  or (_23497_, ABINPUT009[94], _26438_);
  and (_23498_, _23497_, _23496_);
  or (_23500_, ABINPUT009[92], _26433_);
  nand (_23501_, ABINPUT009[90], _26427_);
  and (_23502_, _23501_, _23500_);
  and (_23503_, _23502_, _23498_);
  and (_23504_, _23503_, _23495_);
  and (_23505_, _23504_, _23487_);
  nor (_23506_, ABINPUT009[83], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_23507_, ABINPUT009[83], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_23508_, _23507_, _23506_);
  and (_23509_, ABINPUT009[85], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_23511_, ABINPUT009[85], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_23512_, _23511_, _23509_);
  and (_23513_, _23512_, _23508_);
  nand (_23514_, ABINPUT009[88], _26413_);
  or (_23515_, ABINPUT009[90], _26427_);
  and (_23516_, _23515_, _23514_);
  nand (_23517_, ABINPUT009[86], _26393_);
  or (_23518_, ABINPUT009[88], _26413_);
  and (_23519_, _23518_, _23517_);
  and (_23520_, _23519_, _23516_);
  and (_23522_, _23520_, _23513_);
  or (_23523_, ABINPUT009[78], _26366_);
  nand (_23524_, ABINPUT009[76], _26361_);
  and (_23525_, _23524_, _23523_);
  or (_23526_, ABINPUT009[76], _26361_);
  nand (_23527_, ABINPUT009[74], _26355_);
  and (_23528_, _23527_, _23526_);
  and (_23529_, _23528_, _23525_);
  and (_23530_, ABINPUT009[81], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_23531_, ABINPUT009[81], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_23533_, _23531_, _23530_);
  and (_23534_, ABINPUT009[79], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_23535_, ABINPUT009[79], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_23536_, _23535_, _23534_);
  and (_23537_, _23536_, _23533_);
  and (_23538_, _23537_, _23529_);
  and (_23539_, _23538_, _23522_);
  and (_23540_, ABINPUT009[103], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nor (_23541_, ABINPUT009[103], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_23542_, _23541_, _23540_);
  and (_23544_, ABINPUT009[105], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_23545_, ABINPUT009[105], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_23546_, _23545_, _23544_);
  and (_23547_, _23546_, _23542_);
  nand (_23548_, ABINPUT009[104], _26475_);
  or (_23549_, ABINPUT009[106], _26491_);
  and (_23550_, _23549_, _23548_);
  or (_23551_, ABINPUT009[104], _26475_);
  nand (_23552_, ABINPUT009[102], _26463_);
  and (_23553_, _23552_, _23551_);
  and (_23555_, _23553_, _23550_);
  and (_23556_, _23555_, _23547_);
  and (_23557_, ABINPUT009[91], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_23558_, ABINPUT009[91], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_23559_, _23558_, _23557_);
  and (_23560_, ABINPUT009[93], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_23561_, ABINPUT009[93], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_23562_, _23561_, _23560_);
  and (_23563_, _23562_, _23559_);
  nand (_23564_, ABINPUT009[96], _26443_);
  or (_23566_, ABINPUT009[98], _26450_);
  and (_23567_, _23566_, _23564_);
  or (_23568_, ABINPUT009[96], _26443_);
  nand (_23569_, ABINPUT009[94], _26438_);
  and (_23570_, _23569_, _23568_);
  and (_23571_, _23570_, _23567_);
  and (_23572_, _23571_, _23563_);
  and (_23573_, _23572_, _23556_);
  and (_23574_, _23573_, _23539_);
  and (_23575_, _23574_, _23505_);
  and (_23577_, _23575_, _23471_);
  and (_23578_, _23577_, _23437_);
  and (_23579_, ABINPUT009[119], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nor (_23580_, ABINPUT009[119], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_23581_, _23580_, _23579_);
  and (_23582_, ABINPUT009[121], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_23583_, ABINPUT009[121], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_23584_, _23583_, _23582_);
  and (_23585_, _23584_, _23581_);
  nand (_23586_, ABINPUT009[120], _26541_);
  or (_23588_, ABINPUT009[122], _26547_);
  and (_23589_, _23588_, _23586_);
  nand (_23590_, ABINPUT009[118], _26536_);
  or (_23591_, ABINPUT009[120], _26541_);
  and (_23592_, _23591_, _23590_);
  and (_23593_, _23592_, _23589_);
  and (_23594_, _23593_, _23585_);
  and (_23595_, ABINPUT009[117], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_23596_, ABINPUT009[117], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_23597_, _23596_, _23595_);
  or (_23599_, ABINPUT009[118], _26536_);
  nand (_23600_, ABINPUT009[116], _26531_);
  and (_23601_, _23600_, _23599_);
  and (_23602_, _23601_, _23597_);
  and (_23603_, ABINPUT009[115], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_23604_, ABINPUT009[115], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_23605_, _23604_, _23603_);
  or (_23606_, ABINPUT009[116], _26531_);
  nand (_23607_, ABINPUT009[114], _26525_);
  and (_23608_, _23607_, _23606_);
  and (_23610_, _23608_, _23605_);
  and (_23611_, _23610_, _23602_);
  and (_23612_, _23611_, _23594_);
  and (_23613_, ABINPUT009[109], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_23614_, ABINPUT009[109], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_23615_, _23614_, _23613_);
  and (_23616_, ABINPUT009[107], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_23617_, ABINPUT009[107], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_23618_, _23617_, _23616_);
  and (_23619_, _23618_, _23615_);
  nand (_23621_, ABINPUT009[108], _26505_);
  or (_23622_, ABINPUT009[110], _26513_);
  and (_23623_, _23622_, _23621_);
  or (_23624_, ABINPUT009[108], _26505_);
  nand (_23625_, ABINPUT009[106], _26491_);
  and (_23626_, _23625_, _23624_);
  and (_23627_, _23626_, _23623_);
  and (_23628_, _23627_, _23619_);
  nor (_23629_, ABINPUT009[111], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_23630_, ABINPUT009[111], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_23632_, _23630_, _23629_);
  nor (_23633_, ABINPUT009[113], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_23634_, ABINPUT009[113], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_23635_, _23634_, _23633_);
  or (_23636_, ABINPUT009[114], _26525_);
  nand (_23637_, ABINPUT009[112], _26518_);
  and (_23638_, _23637_, _23636_);
  and (_23639_, _23638_, _23635_);
  and (_23640_, _23639_, _23632_);
  and (_23641_, _23640_, _23628_);
  and (_23643_, _23641_, _23612_);
  or (_23644_, \oc8051_golden_model_1.P0 [6], _24778_);
  or (_23645_, _11620_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_23646_, _23645_, _23644_);
  or (_23647_, _11617_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_23648_, \oc8051_golden_model_1.P0 [4], _24752_);
  and (_23649_, _23648_, _23647_);
  and (_23650_, _23649_, _23646_);
  nor (_23651_, \oc8051_golden_model_1.P1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_23652_, \oc8051_golden_model_1.P1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_23654_, _23652_, _23651_);
  and (_23655_, \oc8051_golden_model_1.P0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_23656_, \oc8051_golden_model_1.P0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_23657_, _23656_, _23655_);
  and (_23658_, _23657_, _23654_);
  and (_23659_, _23658_, _23650_);
  and (_23660_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_23661_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_23662_, _23661_, _23660_);
  and (_23663_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_23665_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_23666_, _23665_, _23663_);
  and (_23667_, _23666_, _23662_);
  or (_23668_, \oc8051_golden_model_1.P1 [2], _24813_);
  or (_23669_, _11625_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_23670_, _23669_, _23668_);
  or (_23671_, _11623_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_23672_, \oc8051_golden_model_1.P1 [0], _24786_);
  and (_23673_, _23672_, _23671_);
  and (_23674_, _23673_, _23670_);
  and (_23676_, _23674_, _23667_);
  and (_23677_, _23676_, _23659_);
  and (_23678_, ABINPUT009[123], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_23679_, ABINPUT009[123], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_23680_, _23679_, _23678_);
  and (_23681_, ABINPUT009[125], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_23682_, ABINPUT009[125], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_23683_, _23682_, _23681_);
  and (_23684_, _23683_, _23680_);
  nand (_23685_, ABINPUT009[124], _26552_);
  or (_23687_, ABINPUT009[126], _26558_);
  and (_23688_, _23687_, _23685_);
  nand (_23689_, ABINPUT009[122], _26547_);
  or (_23690_, ABINPUT009[124], _26552_);
  and (_23691_, _23690_, _23689_);
  and (_23692_, _23691_, _23688_);
  and (_23693_, _23692_, _23684_);
  nor (_23694_, ABINPUT009[127], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_23695_, ABINPUT009[127], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_23696_, _23695_, _23694_);
  nor (_23698_, \oc8051_golden_model_1.P0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_23699_, \oc8051_golden_model_1.P0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_23700_, _23699_, _23698_);
  or (_23701_, _11614_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_23702_, \oc8051_golden_model_1.P0 [2], _24723_);
  and (_23703_, _23702_, _23701_);
  and (_23704_, _23703_, _23700_);
  and (_23705_, _23704_, _23696_);
  and (_23706_, _23705_, _23693_);
  and (_23707_, _23706_, _23677_);
  and (_23709_, _23707_, _23643_);
  or (_23710_, \oc8051_golden_model_1.P0 [0], _24699_);
  nand (_23711_, ABINPUT009[126], _26558_);
  and (_23712_, _23711_, _23710_);
  or (_23713_, ABINPUT009[112], _26518_);
  nand (_23714_, ABINPUT009[110], _26513_);
  and (_23715_, _23714_, _23713_);
  and (_23716_, _23715_, _23712_);
  and (_23717_, _23716_, _23709_);
  or (_23718_, ABINPUT009[72], _26348_);
  nand (_23720_, ABINPUT009[70], _26343_);
  and (_23721_, _23720_, _23718_);
  nor (_23722_, ABINPUT009[67], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_23723_, ABINPUT009[67], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_23724_, _23723_, _23722_);
  and (_23725_, ABINPUT009[69], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_23726_, ABINPUT009[69], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_23727_, _23726_, _23725_);
  and (_23728_, _23727_, _23724_);
  or (_23729_, ABINPUT009[70], _26343_);
  nand (_23731_, ABINPUT009[68], _26337_);
  and (_23732_, _23731_, _23729_);
  or (_23733_, ABINPUT009[68], _26337_);
  nand (_23734_, ABINPUT009[66], _26331_);
  and (_23735_, _23734_, _23733_);
  and (_23736_, _23735_, _23732_);
  and (_23737_, _23736_, _23728_);
  and (_23738_, ABINPUT009[71], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_23739_, ABINPUT009[71], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_23740_, _23739_, _23738_);
  and (_23742_, ABINPUT009[73], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_23743_, ABINPUT009[73], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_23744_, _23743_, _23742_);
  nand (_23745_, ABINPUT009[72], _26348_);
  or (_23746_, ABINPUT009[74], _26355_);
  and (_23747_, _23746_, _23745_);
  and (_23748_, _23747_, _23744_);
  and (_23749_, _23748_, _23740_);
  and (_23750_, _23749_, _23737_);
  and (_23751_, _23750_, _23721_);
  and (_23753_, ABINPUT009[51], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_23754_, ABINPUT009[51], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_23755_, _23754_, _23753_);
  nor (_23756_, ABINPUT009[53], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and (_23757_, ABINPUT009[53], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_23758_, _23757_, _23756_);
  and (_23759_, _23758_, _23755_);
  or (_23760_, ABINPUT009[54], _26294_);
  nand (_23761_, ABINPUT009[52], _26288_);
  and (_23762_, _23761_, _23760_);
  nand (_23764_, ABINPUT009[50], _26281_);
  or (_23765_, ABINPUT009[52], _26288_);
  and (_23766_, _23765_, _23764_);
  and (_23767_, _23766_, _23762_);
  and (_23768_, _23767_, _23759_);
  and (_23769_, ABINPUT009[55], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_23770_, ABINPUT009[55], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_23771_, _23770_, _23769_);
  and (_23772_, ABINPUT009[57], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_23773_, ABINPUT009[57], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_23775_, _23773_, _23772_);
  nand (_23776_, ABINPUT009[56], _26299_);
  or (_23777_, ABINPUT009[58], _26306_);
  and (_23778_, _23777_, _23776_);
  and (_23779_, _23778_, _23775_);
  and (_23780_, _23779_, _23771_);
  and (_23781_, _23780_, _23768_);
  nor (_23782_, ABINPUT009[45], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_23783_, ABINPUT009[45], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_23784_, _23783_, _23782_);
  and (_23786_, ABINPUT009[43], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_23787_, ABINPUT009[43], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_23788_, _23787_, _23786_);
  and (_23789_, _23788_, _23784_);
  or (_23790_, ABINPUT009[46], _26268_);
  nand (_23791_, ABINPUT009[44], _26261_);
  and (_23792_, _23791_, _23790_);
  or (_23793_, ABINPUT009[44], _26261_);
  nand (_23794_, ABINPUT009[42], _26254_);
  and (_23795_, _23794_, _23793_);
  and (_23797_, _23795_, _23792_);
  and (_23798_, _23797_, _23789_);
  and (_23799_, ABINPUT009[47], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor (_23800_, ABINPUT009[47], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_23801_, _23800_, _23799_);
  and (_23802_, ABINPUT009[49], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor (_23803_, ABINPUT009[49], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_23804_, _23803_, _23802_);
  or (_23805_, ABINPUT009[50], _26281_);
  nand (_23806_, ABINPUT009[48], _26273_);
  and (_23808_, _23806_, _23805_);
  and (_23809_, _23808_, _23804_);
  and (_23810_, _23809_, _23801_);
  and (_23811_, _23810_, _23798_);
  and (_23812_, _23811_, _23781_);
  and (_23813_, _23812_, _23751_);
  and (_23814_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_23815_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_23816_, _23815_, _23814_);
  nand (_23817_, _11659_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_23819_, _11659_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_23820_, _23819_, _23817_);
  and (_23821_, _23820_, _23816_);
  or (_23822_, \oc8051_golden_model_1.PSW [4], _25809_);
  or (_23823_, _11663_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_23824_, _23823_, _23822_);
  or (_23825_, \oc8051_golden_model_1.PSW [3], _25583_);
  or (_23826_, _03159_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_23827_, _23826_, _23825_);
  and (_23828_, _23827_, _23824_);
  and (_23830_, _23828_, _23821_);
  or (_23831_, _05348_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_23832_, \oc8051_golden_model_1.PSW [7], _24435_);
  and (_23833_, _23832_, _23831_);
  and (_23834_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_23835_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_23836_, _23835_, _23834_);
  nand (_23837_, _11665_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_23838_, _11665_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_23839_, _23838_, _23837_);
  and (_23841_, _23839_, _23836_);
  and (_23842_, _23841_, _23833_);
  and (_23843_, _23842_, _23830_);
  or (_23844_, _23843_, property_valid_psw_1_r);
  and (_23845_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nor (_23846_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_23847_, _23846_, _23845_);
  and (_23848_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nor (_23849_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  or (_23850_, _23849_, _23848_);
  and (_23852_, _23850_, _23847_);
  or (_23853_, \oc8051_golden_model_1.DPH [2], _28519_);
  or (_23854_, _05254_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_23855_, _23854_, _23853_);
  or (_23856_, _10168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_23857_, \oc8051_golden_model_1.DPH [0], _28434_);
  and (_23858_, _23857_, _23856_);
  and (_23859_, _23858_, _23855_);
  and (_23860_, _23859_, _23852_);
  nor (_23861_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_23863_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_23864_, _23863_, _23861_);
  or (_23865_, _10147_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_23866_, \oc8051_golden_model_1.B [6], _19723_);
  and (_23867_, _23866_, _23865_);
  and (_23868_, _23867_, _23864_);
  nor (_23869_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_23870_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_23871_, _23870_, _23869_);
  or (_23872_, \oc8051_golden_model_1.B [4], _19383_);
  or (_23874_, _10144_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_23875_, _23874_, _23872_);
  and (_23876_, _23875_, _23871_);
  and (_23877_, _23876_, _23868_);
  and (_23878_, _23877_, _23860_);
  nor (_23879_, \oc8051_golden_model_1.DPL [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_23880_, \oc8051_golden_model_1.DPL [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  or (_23881_, _23880_, _23879_);
  and (_23882_, \oc8051_golden_model_1.B [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor (_23883_, \oc8051_golden_model_1.B [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_23885_, _23883_, _23882_);
  and (_23886_, _23885_, _23881_);
  nand (_23887_, _10162_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  or (_23888_, _10159_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_23889_, _23888_, _23887_);
  or (_23890_, _10150_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_23891_, _10159_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_23892_, _23891_, _23890_);
  and (_23893_, _23892_, _23889_);
  and (_23894_, _23893_, _23886_);
  nand (_23896_, _10168_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_23897_, _10165_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_23898_, _23897_, _23896_);
  or (_23899_, _10162_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_23900_, _10165_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_23901_, _23900_, _23899_);
  and (_23902_, _23901_, _23898_);
  and (_23903_, \oc8051_golden_model_1.DPL [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nor (_23904_, \oc8051_golden_model_1.DPL [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  or (_23905_, _23904_, _23903_);
  and (_23907_, \oc8051_golden_model_1.DPH [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_23908_, \oc8051_golden_model_1.DPH [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_23909_, _23908_, _23907_);
  and (_23910_, _23909_, _23905_);
  and (_23911_, _23910_, _23902_);
  and (_23912_, _23911_, _23894_);
  and (_23913_, _23912_, _23878_);
  or (_23914_, _10175_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_23915_, \oc8051_golden_model_1.DPH [6], _28703_);
  and (_23916_, _23915_, _23914_);
  or (_23918_, \oc8051_golden_model_1.DPH [4], _28612_);
  or (_23919_, _10172_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_23920_, _23919_, _23918_);
  and (_23921_, _23920_, _23916_);
  and (_23922_, \oc8051_golden_model_1.DPH [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_23923_, \oc8051_golden_model_1.DPH [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_23924_, _23923_, _23922_);
  and (_23925_, ABINPUT009[1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_23926_, ABINPUT009[1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_23927_, _23926_, _23925_);
  and (_23929_, _23927_, _23924_);
  and (_23930_, _23929_, _23921_);
  nor (_23931_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_23932_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_23933_, _23932_, _23931_);
  nor (_23934_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_23935_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_23936_, _23935_, _23934_);
  and (_23937_, _23936_, _23933_);
  or (_23938_, ABINPUT009[2], _26073_);
  nand (_23940_, ABINPUT009[0], _26034_);
  and (_23941_, _23940_, _23938_);
  or (_23942_, _10178_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_23943_, ABINPUT009[0], _26034_);
  and (_23944_, _23943_, _23942_);
  and (_23945_, _23944_, _23941_);
  and (_23946_, _23945_, _23937_);
  and (_23947_, _23946_, _23930_);
  nor (_23948_, ABINPUT009[3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_23949_, ABINPUT009[3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_23951_, _23949_, _23948_);
  and (_23952_, ABINPUT009[5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_23953_, ABINPUT009[5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_23954_, _23953_, _23952_);
  and (_23955_, _23954_, _23951_);
  or (_23956_, ABINPUT009[6], _26135_);
  nand (_23957_, ABINPUT009[4], _26105_);
  and (_23958_, _23957_, _23956_);
  or (_23959_, ABINPUT009[4], _26105_);
  nand (_23960_, ABINPUT009[2], _26073_);
  and (_23962_, _23960_, _23959_);
  and (_23963_, _23962_, _23958_);
  and (_23964_, _23963_, _23955_);
  and (_23965_, ABINPUT009[7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_23966_, ABINPUT009[7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_23967_, _23966_, _23965_);
  and (_23968_, ABINPUT009[9], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_23969_, ABINPUT009[9], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_23970_, _23969_, _23968_);
  or (_23971_, ABINPUT009[10], _26160_);
  nand (_23973_, ABINPUT009[8], _26152_);
  and (_23974_, _23973_, _23971_);
  and (_23975_, _23974_, _23970_);
  and (_23976_, _23975_, _23967_);
  and (_23977_, _23976_, _23964_);
  and (_23978_, _23977_, _23947_);
  and (_23979_, _23978_, _23913_);
  and (_23980_, _23979_, _23844_);
  and (_23981_, _23980_, _23813_);
  and (_23982_, _23981_, _23717_);
  and (_23984_, _23982_, _23578_);
  or (_23985_, _24288_, \oc8051_golden_model_1.SP [7]);
  nand (_23986_, _24288_, \oc8051_golden_model_1.SP [7]);
  and (_23987_, _23986_, _23985_);
  or (_23988_, _24332_, \oc8051_golden_model_1.SP [6]);
  nand (_23989_, _24332_, \oc8051_golden_model_1.SP [6]);
  and (_23990_, _23989_, _23988_);
  or (_23991_, _24326_, \oc8051_golden_model_1.SP [5]);
  nand (_23992_, _24326_, \oc8051_golden_model_1.SP [5]);
  and (_23993_, _23992_, _23991_);
  nand (_23995_, _24314_, \oc8051_golden_model_1.SP [3]);
  or (_23996_, _24314_, \oc8051_golden_model_1.SP [3]);
  and (_23997_, _23996_, _23995_);
  nand (_23998_, _24302_, \oc8051_golden_model_1.SP [1]);
  nand (_23999_, _24296_, \oc8051_golden_model_1.SP [0]);
  or (_24000_, _24296_, \oc8051_golden_model_1.SP [0]);
  and (_24001_, _24000_, _23999_);
  or (_24002_, _24302_, \oc8051_golden_model_1.SP [1]);
  and (_24003_, _24002_, _24001_);
  and (_24004_, _24003_, _23998_);
  or (_24006_, _24308_, \oc8051_golden_model_1.SP [2]);
  nand (_24007_, _24308_, \oc8051_golden_model_1.SP [2]);
  and (_24008_, _24007_, _24006_);
  and (_24009_, _24008_, _24004_);
  and (_24010_, _24009_, _23997_);
  or (_24011_, _24320_, \oc8051_golden_model_1.SP [4]);
  nand (_24012_, _24320_, \oc8051_golden_model_1.SP [4]);
  and (_24013_, _24012_, _24011_);
  and (_24014_, _24013_, _24010_);
  and (_24015_, _24014_, _23993_);
  and (_24017_, _24015_, _23990_);
  and (_24018_, _24017_, _23987_);
  or (_24019_, _24018_, property_valid_sp_1_r);
  nand (_24020_, ABINPUT009[6], _26135_);
  or (_24021_, ABINPUT009[8], _26152_);
  and (_24022_, _24021_, _24020_);
  or (_24023_, \oc8051_golden_model_1.B [0], _18595_);
  or (_24024_, _09265_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_24025_, _24024_, _24023_);
  or (_24026_, \oc8051_golden_model_1.ACC [0], _27945_);
  and (_24027_, _24026_, p1_valid_r);
  or (_24028_, _02059_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_24029_, \oc8051_golden_model_1.ACC [2], _24571_);
  and (_24030_, _24029_, _24028_);
  and (_24031_, _24030_, _24027_);
  and (_24032_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_24033_, \oc8051_golden_model_1.ACC [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_24034_, _24033_, _24032_);
  and (_24035_, _24034_, inst_finished_r);
  and (_24036_, _24035_, _24031_);
  nor (_24037_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_24038_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_24039_, _24038_, _24037_);
  and (_24040_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_24041_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_24042_, _24041_, _24040_);
  and (_24043_, _24042_, _24039_);
  or (_24044_, _08826_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_24045_, \oc8051_golden_model_1.ACC [6], _24614_);
  and (_24046_, _24045_, _24044_);
  or (_24048_, _08384_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_24049_, \oc8051_golden_model_1.ACC [4], _24592_);
  and (_24050_, _24049_, _24048_);
  and (_24051_, _24050_, _24046_);
  and (_24052_, _24051_, _24043_);
  and (_24053_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_24054_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_24055_, _24054_, _24053_);
  or (_24056_, _10141_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_24057_, \oc8051_golden_model_1.B [2], _19021_);
  and (_24059_, _24057_, _24056_);
  nor (_24060_, \oc8051_golden_model_1.B [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_24061_, \oc8051_golden_model_1.B [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_24062_, _24061_, _24060_);
  and (_24063_, _24062_, _24059_);
  and (_24064_, _24063_, _24055_);
  and (_24065_, _24064_, _24052_);
  and (_24066_, _24065_, _24036_);
  and (_24067_, _24066_, _24025_);
  and (_24068_, _24067_, _24022_);
  nand (_24070_, ABINPUT009[20], _26190_);
  or (_24071_, ABINPUT009[22], _26195_);
  and (_24072_, _24071_, _24070_);
  nand (_24073_, ABINPUT009[18], _26185_);
  or (_24074_, ABINPUT009[20], _26190_);
  and (_24075_, _24074_, _24073_);
  and (_24076_, _24075_, _24072_);
  nor (_24077_, ABINPUT009[25], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  and (_24078_, ABINPUT009[25], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_24079_, _24078_, _24077_);
  and (_24081_, ABINPUT009[23], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_24082_, ABINPUT009[23], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_24083_, _24082_, _24081_);
  and (_24084_, _24083_, _24079_);
  and (_24085_, _24084_, _24076_);
  and (_24086_, ABINPUT009[11], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_24087_, ABINPUT009[11], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_24088_, _24087_, _24086_);
  and (_24089_, ABINPUT009[13], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_24090_, ABINPUT009[13], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_24092_, _24090_, _24089_);
  and (_24093_, _24092_, _24088_);
  nand (_24094_, ABINPUT009[16], _26177_);
  or (_24095_, ABINPUT009[18], _26185_);
  and (_24096_, _24095_, _24094_);
  or (_24097_, ABINPUT009[16], _26177_);
  nand (_24098_, ABINPUT009[14], _26172_);
  and (_24099_, _24098_, _24097_);
  and (_24100_, _24099_, _24096_);
  and (_24101_, _24100_, _24093_);
  and (_24103_, _24101_, _24085_);
  nor (_24104_, ABINPUT009[37], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_24105_, ABINPUT009[37], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_24106_, _24105_, _24104_);
  and (_24107_, ABINPUT009[35], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_24108_, ABINPUT009[35], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_24109_, _24108_, _24107_);
  and (_24110_, _24109_, _24106_);
  nand (_24111_, ABINPUT009[38], _26241_);
  or (_24112_, ABINPUT009[40], _26246_);
  and (_24114_, _24112_, _24111_);
  or (_24115_, ABINPUT009[42], _26254_);
  nand (_24116_, ABINPUT009[40], _26246_);
  and (_24117_, _24116_, _24115_);
  and (_24118_, _24117_, _24114_);
  and (_24119_, _24118_, _24110_);
  nand (_24120_, ABINPUT009[28], _26212_);
  or (_24121_, ABINPUT009[30], _26217_);
  and (_24122_, _24121_, _24120_);
  or (_24123_, ABINPUT009[28], _26212_);
  nand (_24125_, ABINPUT009[26], _26207_);
  and (_24126_, _24125_, _24123_);
  and (_24127_, _24126_, _24122_);
  nor (_24128_, ABINPUT009[31], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_24129_, ABINPUT009[31], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_24130_, _24129_, _24128_);
  and (_24131_, ABINPUT009[33], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_24132_, ABINPUT009[33], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_24133_, _24132_, _24131_);
  and (_24134_, _24133_, _24130_);
  and (_24136_, _24134_, _24127_);
  and (_24137_, _24136_, _24119_);
  and (_24138_, _24137_, _24103_);
  nor (_24139_, ABINPUT009[19], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_24140_, ABINPUT009[19], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_24141_, _24140_, _24139_);
  and (_24142_, ABINPUT009[21], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_24143_, ABINPUT009[21], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_24144_, _24143_, _24142_);
  and (_24145_, _24144_, _24141_);
  nand (_24147_, ABINPUT009[24], _26200_);
  or (_24148_, ABINPUT009[26], _26207_);
  and (_24149_, _24148_, _24147_);
  nand (_24150_, ABINPUT009[22], _26195_);
  or (_24151_, ABINPUT009[24], _26200_);
  and (_24152_, _24151_, _24150_);
  and (_24153_, _24152_, _24149_);
  and (_24154_, _24153_, _24145_);
  nand (_24155_, ABINPUT009[12], _26166_);
  or (_24156_, ABINPUT009[14], _26172_);
  and (_24158_, _24156_, _24155_);
  nand (_24159_, ABINPUT009[10], _26160_);
  or (_24160_, ABINPUT009[12], _26166_);
  and (_24161_, _24160_, _24159_);
  and (_24162_, _24161_, _24158_);
  nor (_24163_, ABINPUT009[17], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_24164_, ABINPUT009[17], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_24165_, _24164_, _24163_);
  nor (_24166_, ABINPUT009[15], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_24167_, ABINPUT009[15], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_24169_, _24167_, _24166_);
  and (_24170_, _24169_, _24165_);
  and (_24171_, _24170_, _24162_);
  and (_24172_, _24171_, _24154_);
  nand (_24173_, ABINPUT009[36], _26235_);
  or (_24174_, ABINPUT009[38], _26241_);
  and (_24175_, _24174_, _24173_);
  nand (_24176_, ABINPUT009[34], _26230_);
  or (_24177_, ABINPUT009[36], _26235_);
  and (_24178_, _24177_, _24176_);
  and (_24180_, _24178_, _24175_);
  nor (_24181_, ABINPUT009[39], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_24182_, ABINPUT009[39], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_24183_, _24182_, _24181_);
  and (_24184_, ABINPUT009[41], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_24185_, ABINPUT009[41], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_24186_, _24185_, _24184_);
  and (_24187_, _24186_, _24183_);
  and (_24188_, _24187_, _24180_);
  nor (_24189_, ABINPUT009[27], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_24191_, ABINPUT009[27], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_24192_, _24191_, _24189_);
  nor (_24193_, ABINPUT009[29], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_24194_, ABINPUT009[29], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_24195_, _24194_, _24193_);
  and (_24196_, _24195_, _24192_);
  nand (_24197_, ABINPUT009[32], _26222_);
  or (_24198_, ABINPUT009[34], _26230_);
  and (_24199_, _24198_, _24197_);
  or (_24200_, ABINPUT009[32], _26222_);
  nand (_24202_, ABINPUT009[30], _26217_);
  and (_24203_, _24202_, _24200_);
  and (_24204_, _24203_, _24199_);
  and (_24205_, _24204_, _24196_);
  and (_24206_, _24205_, _24188_);
  and (_24207_, _24206_, _24172_);
  and (_24208_, _24207_, _24138_);
  or (_24209_, ABINPUT009[56], _26299_);
  nand (_24210_, ABINPUT009[54], _26294_);
  and (_24211_, _24210_, _24209_);
  or (_24213_, ABINPUT009[48], _26273_);
  nand (_24214_, ABINPUT009[46], _26268_);
  and (_24215_, _24214_, _24213_);
  and (_24216_, _24215_, _24211_);
  or (_24217_, ABINPUT009[62], _26318_);
  nand (_24218_, ABINPUT009[60], _26312_);
  and (_24219_, _24218_, _24217_);
  or (_24220_, ABINPUT009[60], _26312_);
  nand (_24221_, ABINPUT009[58], _26306_);
  and (_24222_, _24221_, _24220_);
  and (_24224_, _24222_, _24219_);
  and (_24225_, ABINPUT009[63], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_24226_, ABINPUT009[63], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_24227_, _24226_, _24225_);
  and (_24228_, ABINPUT009[65], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_24229_, ABINPUT009[65], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_24230_, _24229_, _24228_);
  and (_24231_, _24230_, _24227_);
  and (_24232_, ABINPUT009[59], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_24233_, ABINPUT009[59], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_24235_, _24233_, _24232_);
  and (_24236_, ABINPUT009[61], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor (_24237_, ABINPUT009[61], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_24238_, _24237_, _24236_);
  and (_24239_, _24238_, _24235_);
  nand (_24240_, ABINPUT009[64], _26323_);
  or (_24241_, ABINPUT009[66], _26331_);
  and (_24242_, _24241_, _24240_);
  nand (_24243_, ABINPUT009[62], _26318_);
  or (_24244_, ABINPUT009[64], _26323_);
  and (_24246_, _24244_, _24243_);
  and (_24247_, _24246_, _24242_);
  and (_24248_, _24247_, _24239_);
  and (_24249_, _24248_, _24231_);
  and (_24250_, _24249_, _24224_);
  and (_24251_, _24250_, _24216_);
  and (_24252_, _24251_, _24208_);
  and (_24253_, _24252_, _24068_);
  and (_24254_, _24253_, _24019_);
  and (_24255_, _24254_, _23984_);
  or (_24257_, _24255_, rst);
  and (_00000_, _24257_, _00009_);
  nor (_00002_[7], _28149_, rst);
  and (_24258_, _27788_, eq_state);
  and (_24259_, _24258_, _01954_);
  and (_24260_, _24259_, _02672_);
  and (property_invalid_pc, _24260_, _23342_);
  buf (_00064_, _27053_);
  buf (_00111_, _27053_);
  buf (_00161_, _27053_);
  buf (_00212_, _27053_);
  buf (_00264_, _27053_);
  buf (_00315_, _27053_);
  buf (_00365_, _27053_);
  buf (_00418_, _27053_);
  buf (_00470_, _27053_);
  buf (_00522_, _27053_);
  buf (_00573_, _27053_);
  buf (_00626_, _27053_);
  buf (_00678_, _27053_);
  buf (_00730_, _27053_);
  buf (_00782_, _27053_);
  buf (_00834_, _27053_);
  buf (_03145_, _00910_);
  buf (_03148_, _00914_);
  buf (_03182_, _00910_);
  buf (_03185_, _00914_);
  buf (_05659_, _01056_);
  buf (_05661_, _01059_);
  buf (_05663_, _01062_);
  buf (_05665_, _01065_);
  buf (_05667_, _01068_);
  buf (_05669_, _01071_);
  buf (_05671_, _01074_);
  buf (_05673_, _01077_);
  buf (_05675_, _01080_);
  buf (_05677_, _01083_);
  buf (_05679_, _01086_);
  buf (_05681_, _01089_);
  buf (_05683_, _01091_);
  buf (_05685_, _01094_);
  buf (_05779_, _01056_);
  buf (_05781_, _01059_);
  buf (_05783_, _01062_);
  buf (_05785_, _01065_);
  buf (_05787_, _01068_);
  buf (_05789_, _01071_);
  buf (_05791_, _01074_);
  buf (_05793_, _01077_);
  buf (_05795_, _01080_);
  buf (_05797_, _01083_);
  buf (_05799_, _01086_);
  buf (_05801_, _01089_);
  buf (_05803_, _01091_);
  buf (_05805_, _01094_);
  buf (_08171_, _01513_);
  buf (_08274_, _01513_);
  dff (p0in_reg[0], _00002_[0]);
  dff (p0in_reg[1], _00002_[1]);
  dff (p0in_reg[2], _00002_[2]);
  dff (p0in_reg[3], _00002_[3]);
  dff (p0in_reg[4], _00002_[4]);
  dff (p0in_reg[5], _00002_[5]);
  dff (p0in_reg[6], _00002_[6]);
  dff (p0in_reg[7], _00002_[7]);
  dff (p1in_reg[0], _00004_[0]);
  dff (p1in_reg[1], _00004_[1]);
  dff (p1in_reg[2], _00004_[2]);
  dff (p1in_reg[3], _00004_[3]);
  dff (p1in_reg[4], _00004_[4]);
  dff (p1in_reg[5], _00004_[5]);
  dff (p1in_reg[6], _00004_[6]);
  dff (p1in_reg[7], _00004_[7]);
  dff (p2in_reg[0], _00005_[0]);
  dff (p2in_reg[1], _00005_[1]);
  dff (p2in_reg[2], _00005_[2]);
  dff (p2in_reg[3], _00005_[3]);
  dff (p2in_reg[4], _00005_[4]);
  dff (p2in_reg[5], _00005_[5]);
  dff (p2in_reg[6], _00005_[6]);
  dff (p2in_reg[7], _00005_[7]);
  dff (p3in_reg[0], _00006_[0]);
  dff (p3in_reg[1], _00006_[1]);
  dff (p3in_reg[2], _00006_[2]);
  dff (p3in_reg[3], _00006_[3]);
  dff (p3in_reg[4], _00006_[4]);
  dff (p3in_reg[5], _00006_[5]);
  dff (p3in_reg[6], _00006_[6]);
  dff (p3in_reg[7], _00006_[7]);
  dff (inst_finished_r, _00001_);
  dff (regs_always_zero, _00009_);
  dff (property_valid_psw_1_r, _00007_);
  dff (property_valid_sp_1_r, _00008_);
  dff (p1_valid_r, _00003_);
  dff (eq_state, _00000_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _00088_);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _00090_);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _00092_);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _00094_);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _00096_);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _00098_);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _00100_);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _00062_);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _00064_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _00140_);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _00142_);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _00144_);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _00146_);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _00148_);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _00149_);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _00151_);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _00108_);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _00111_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _00603_);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _00605_);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _00607_);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _00609_);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _00611_);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _00613_);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _00615_);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _00571_);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _00573_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _00655_);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _00657_);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _00659_);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _00661_);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _00663_);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _00665_);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _00667_);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _00623_);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _00626_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _00707_);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _00709_);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _00711_);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _00713_);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _00715_);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _00717_);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _00719_);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _00675_);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _00678_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _00759_);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _00761_);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _00763_);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _00765_);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _00767_);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _00769_);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _00771_);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _00727_);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _00730_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _00811_);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _00813_);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _00815_);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _00817_);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _00819_);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _00821_);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _00823_);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _00779_);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _00782_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _00863_);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _00865_);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _00867_);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _00869_);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _00871_);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _00873_);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _00875_);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _00831_);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _00834_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _00190_);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _00192_);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _00194_);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _00196_);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _00198_);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _00200_);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _00202_);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _00158_);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _00161_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _00241_);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _00243_);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _00245_);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _00247_);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _00249_);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _00251_);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _00253_);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _00210_);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _00212_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _00292_);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _00294_);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _00296_);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _00298_);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _00300_);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _00302_);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _00304_);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _00261_);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _00264_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _00343_);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _00345_);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _00347_);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _00349_);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _00351_);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _00352_);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _00354_);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _00312_);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _00315_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _00395_);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _00397_);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _00399_);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _00401_);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _00403_);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _00405_);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _00407_);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _00362_);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _00365_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _00448_);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _00450_);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _00452_);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _00454_);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _00456_);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _00458_);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _00460_);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _00415_);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _00418_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _00499_);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _00501_);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _00503_);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _00505_);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _00507_);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _00509_);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _00511_);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _00467_);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _00470_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _00551_);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _00553_);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _00555_);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _00557_);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _00559_);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _00561_);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _00563_);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _00519_);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _00522_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _30702_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _30703_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _30704_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _30705_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _30706_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _30707_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _30708_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _30709_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _30758_[0]);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _30758_[1]);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _30758_[2]);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _30758_[3]);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _30758_[4]);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _30758_[5]);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _30758_[6]);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _30758_[7]);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _30757_[0]);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _30757_[1]);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _30757_[2]);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _30757_[3]);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _30757_[4]);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _30757_[5]);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _30757_[6]);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _30757_[7]);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _30756_[0]);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _30756_[1]);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _30756_[2]);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _30756_[3]);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _30756_[4]);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _30756_[5]);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _30756_[6]);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _30756_[7]);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _30755_[0]);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _30755_[1]);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _30755_[2]);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _30755_[3]);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _30755_[4]);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _30755_[5]);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _30755_[6]);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _30755_[7]);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _30754_[0]);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _30754_[1]);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _30754_[2]);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _30754_[3]);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _30754_[4]);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _30754_[5]);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _30754_[6]);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _30754_[7]);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _30710_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _30711_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _30712_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _30753_[3]);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _30753_[4]);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _30753_[5]);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _30753_[6]);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _30753_[7]);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _30745_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _30746_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _30747_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _30748_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _30749_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _30750_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _30751_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _30752_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _30737_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _30738_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _30739_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _30740_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _30741_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _30742_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _30743_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _30744_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _30729_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _30730_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _30731_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _30732_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _30733_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _30734_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _30735_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _30736_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _30721_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _30722_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _30723_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _30724_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _30725_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _30726_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _30727_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _30728_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _30762_[0]);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _30762_[1]);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _30762_[2]);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _30762_[3]);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _30762_[4]);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _30762_[5]);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _30762_[6]);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _30762_[7]);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _30761_[0]);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _30761_[1]);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _30761_[2]);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _30761_[3]);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _30761_[4]);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _30761_[5]);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _30761_[6]);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _30761_[7]);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _30760_[0]);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _30760_[1]);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _30760_[2]);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _30760_[3]);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _30760_[4]);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _30760_[5]);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _30760_[6]);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _30760_[7]);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _30759_[0]);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _30759_[1]);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _30759_[2]);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _30759_[3]);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _30759_[4]);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _30759_[5]);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _30759_[6]);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _30759_[7]);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _30713_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _30714_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _30715_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _30716_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _30717_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _30718_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _30719_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _30720_);
  dff (\oc8051_golden_model_1.B [0], _28763_);
  dff (\oc8051_golden_model_1.B [1], _28764_);
  dff (\oc8051_golden_model_1.B [2], _28767_);
  dff (\oc8051_golden_model_1.B [3], _28768_);
  dff (\oc8051_golden_model_1.B [4], _28769_);
  dff (\oc8051_golden_model_1.B [5], _28770_);
  dff (\oc8051_golden_model_1.B [6], _28771_);
  dff (\oc8051_golden_model_1.B [7], _26422_);
  dff (\oc8051_golden_model_1.ACC [0], _28773_);
  dff (\oc8051_golden_model_1.ACC [1], _28776_);
  dff (\oc8051_golden_model_1.ACC [2], _28777_);
  dff (\oc8051_golden_model_1.ACC [3], _28778_);
  dff (\oc8051_golden_model_1.ACC [4], _28779_);
  dff (\oc8051_golden_model_1.ACC [5], _28780_);
  dff (\oc8051_golden_model_1.ACC [6], _28781_);
  dff (\oc8051_golden_model_1.ACC [7], _26420_);
  dff (\oc8051_golden_model_1.DPL [0], _28783_);
  dff (\oc8051_golden_model_1.DPL [1], _28784_);
  dff (\oc8051_golden_model_1.DPL [2], _28785_);
  dff (\oc8051_golden_model_1.DPL [3], _28786_);
  dff (\oc8051_golden_model_1.DPL [4], _28787_);
  dff (\oc8051_golden_model_1.DPL [5], _28788_);
  dff (\oc8051_golden_model_1.DPL [6], _28789_);
  dff (\oc8051_golden_model_1.DPL [7], _26419_);
  dff (\oc8051_golden_model_1.DPH [0], _28794_);
  dff (\oc8051_golden_model_1.DPH [1], _28795_);
  dff (\oc8051_golden_model_1.DPH [2], _28796_);
  dff (\oc8051_golden_model_1.DPH [3], _28797_);
  dff (\oc8051_golden_model_1.DPH [4], _28798_);
  dff (\oc8051_golden_model_1.DPH [5], _28799_);
  dff (\oc8051_golden_model_1.DPH [6], _28800_);
  dff (\oc8051_golden_model_1.DPH [7], _26418_);
  dff (\oc8051_golden_model_1.IE [0], _28801_);
  dff (\oc8051_golden_model_1.IE [1], _28802_);
  dff (\oc8051_golden_model_1.IE [2], _28803_);
  dff (\oc8051_golden_model_1.IE [3], _28804_);
  dff (\oc8051_golden_model_1.IE [4], _28805_);
  dff (\oc8051_golden_model_1.IE [5], _28808_);
  dff (\oc8051_golden_model_1.IE [6], _28809_);
  dff (\oc8051_golden_model_1.IE [7], _26417_);
  dff (\oc8051_golden_model_1.IP [0], _28810_);
  dff (\oc8051_golden_model_1.IP [1], _28813_);
  dff (\oc8051_golden_model_1.IP [2], _28814_);
  dff (\oc8051_golden_model_1.IP [3], _28815_);
  dff (\oc8051_golden_model_1.IP [4], _28816_);
  dff (\oc8051_golden_model_1.IP [5], _28817_);
  dff (\oc8051_golden_model_1.IP [6], _28818_);
  dff (\oc8051_golden_model_1.IP [7], _26415_);
  dff (\oc8051_golden_model_1.P0 [0], _28821_);
  dff (\oc8051_golden_model_1.P0 [1], _28822_);
  dff (\oc8051_golden_model_1.P0 [2], _28823_);
  dff (\oc8051_golden_model_1.P0 [3], _28824_);
  dff (\oc8051_golden_model_1.P0 [4], _28825_);
  dff (\oc8051_golden_model_1.P0 [5], _28826_);
  dff (\oc8051_golden_model_1.P0 [6], _28827_);
  dff (\oc8051_golden_model_1.P0 [7], _26414_);
  dff (\oc8051_golden_model_1.P1 [0], _28830_);
  dff (\oc8051_golden_model_1.P1 [1], _28831_);
  dff (\oc8051_golden_model_1.P1 [2], _28832_);
  dff (\oc8051_golden_model_1.P1 [3], _28833_);
  dff (\oc8051_golden_model_1.P1 [4], _28834_);
  dff (\oc8051_golden_model_1.P1 [5], _28835_);
  dff (\oc8051_golden_model_1.P1 [6], _28836_);
  dff (\oc8051_golden_model_1.P1 [7], _26412_);
  dff (\oc8051_golden_model_1.P2 [0], _28841_);
  dff (\oc8051_golden_model_1.P2 [1], _28842_);
  dff (\oc8051_golden_model_1.P2 [2], _28843_);
  dff (\oc8051_golden_model_1.P2 [3], _28844_);
  dff (\oc8051_golden_model_1.P2 [4], _28845_);
  dff (\oc8051_golden_model_1.P2 [5], _28846_);
  dff (\oc8051_golden_model_1.P2 [6], _28847_);
  dff (\oc8051_golden_model_1.P2 [7], _26411_);
  dff (\oc8051_golden_model_1.P3 [0], _28850_);
  dff (\oc8051_golden_model_1.P3 [1], _28851_);
  dff (\oc8051_golden_model_1.P3 [2], _28852_);
  dff (\oc8051_golden_model_1.P3 [3], _28853_);
  dff (\oc8051_golden_model_1.P3 [4], _28854_);
  dff (\oc8051_golden_model_1.P3 [5], _28855_);
  dff (\oc8051_golden_model_1.P3 [6], _28856_);
  dff (\oc8051_golden_model_1.P3 [7], _26410_);
  dff (\oc8051_golden_model_1.PSW [0], _28859_);
  dff (\oc8051_golden_model_1.PSW [1], _28860_);
  dff (\oc8051_golden_model_1.PSW [2], _28861_);
  dff (\oc8051_golden_model_1.PSW [3], _28862_);
  dff (\oc8051_golden_model_1.PSW [4], _28863_);
  dff (\oc8051_golden_model_1.PSW [5], _28864_);
  dff (\oc8051_golden_model_1.PSW [6], _28867_);
  dff (\oc8051_golden_model_1.PSW [7], _26409_);
  dff (\oc8051_golden_model_1.PCON [0], _28868_);
  dff (\oc8051_golden_model_1.PCON [1], _28869_);
  dff (\oc8051_golden_model_1.PCON [2], _28872_);
  dff (\oc8051_golden_model_1.PCON [3], _28873_);
  dff (\oc8051_golden_model_1.PCON [4], _28874_);
  dff (\oc8051_golden_model_1.PCON [5], _28875_);
  dff (\oc8051_golden_model_1.PCON [6], _28876_);
  dff (\oc8051_golden_model_1.PCON [7], _26407_);
  dff (\oc8051_golden_model_1.SBUF [0], _28877_);
  dff (\oc8051_golden_model_1.SBUF [1], _28878_);
  dff (\oc8051_golden_model_1.SBUF [2], _28879_);
  dff (\oc8051_golden_model_1.SBUF [3], _28880_);
  dff (\oc8051_golden_model_1.SBUF [4], _28881_);
  dff (\oc8051_golden_model_1.SBUF [5], _28882_);
  dff (\oc8051_golden_model_1.SBUF [6], _28883_);
  dff (\oc8051_golden_model_1.SBUF [7], _26406_);
  dff (\oc8051_golden_model_1.SCON [0], _28886_);
  dff (\oc8051_golden_model_1.SCON [1], _28887_);
  dff (\oc8051_golden_model_1.SCON [2], _28888_);
  dff (\oc8051_golden_model_1.SCON [3], _28889_);
  dff (\oc8051_golden_model_1.SCON [4], _28892_);
  dff (\oc8051_golden_model_1.SCON [5], _28893_);
  dff (\oc8051_golden_model_1.SCON [6], _28894_);
  dff (\oc8051_golden_model_1.SCON [7], _26404_);
  dff (\oc8051_golden_model_1.SP [0], _28896_);
  dff (\oc8051_golden_model_1.SP [1], _28897_);
  dff (\oc8051_golden_model_1.SP [2], _28898_);
  dff (\oc8051_golden_model_1.SP [3], _28899_);
  dff (\oc8051_golden_model_1.SP [4], _28900_);
  dff (\oc8051_golden_model_1.SP [5], _28901_);
  dff (\oc8051_golden_model_1.SP [6], _28902_);
  dff (\oc8051_golden_model_1.SP [7], _26403_);
  dff (\oc8051_golden_model_1.TCON [0], _28905_);
  dff (\oc8051_golden_model_1.TCON [1], _28906_);
  dff (\oc8051_golden_model_1.TCON [2], _28907_);
  dff (\oc8051_golden_model_1.TCON [3], _28908_);
  dff (\oc8051_golden_model_1.TCON [4], _28909_);
  dff (\oc8051_golden_model_1.TCON [5], _28910_);
  dff (\oc8051_golden_model_1.TCON [6], _28912_);
  dff (\oc8051_golden_model_1.TCON [7], _26402_);
  dff (\oc8051_golden_model_1.TH0 [0], _28913_);
  dff (\oc8051_golden_model_1.TH0 [1], _28914_);
  dff (\oc8051_golden_model_1.TH0 [2], _28915_);
  dff (\oc8051_golden_model_1.TH0 [3], _28916_);
  dff (\oc8051_golden_model_1.TH0 [4], _28917_);
  dff (\oc8051_golden_model_1.TH0 [5], _28918_);
  dff (\oc8051_golden_model_1.TH0 [6], _28919_);
  dff (\oc8051_golden_model_1.TH0 [7], _26400_);
  dff (\oc8051_golden_model_1.TH1 [0], _28922_);
  dff (\oc8051_golden_model_1.TH1 [1], _28923_);
  dff (\oc8051_golden_model_1.TH1 [2], _28924_);
  dff (\oc8051_golden_model_1.TH1 [3], _28925_);
  dff (\oc8051_golden_model_1.TH1 [4], _28926_);
  dff (\oc8051_golden_model_1.TH1 [5], _28927_);
  dff (\oc8051_golden_model_1.TH1 [6], _28928_);
  dff (\oc8051_golden_model_1.TH1 [7], _26399_);
  dff (\oc8051_golden_model_1.TL0 [0], _28931_);
  dff (\oc8051_golden_model_1.TL0 [1], _28932_);
  dff (\oc8051_golden_model_1.TL0 [2], _28933_);
  dff (\oc8051_golden_model_1.TL0 [3], _28934_);
  dff (\oc8051_golden_model_1.TL0 [4], _28935_);
  dff (\oc8051_golden_model_1.TL0 [5], _28936_);
  dff (\oc8051_golden_model_1.TL0 [6], _28937_);
  dff (\oc8051_golden_model_1.TL0 [7], _26398_);
  dff (\oc8051_golden_model_1.TL1 [0], _28940_);
  dff (\oc8051_golden_model_1.TL1 [1], _28941_);
  dff (\oc8051_golden_model_1.TL1 [2], _28942_);
  dff (\oc8051_golden_model_1.TL1 [3], _28943_);
  dff (\oc8051_golden_model_1.TL1 [4], _28944_);
  dff (\oc8051_golden_model_1.TL1 [5], _28945_);
  dff (\oc8051_golden_model_1.TL1 [6], _28946_);
  dff (\oc8051_golden_model_1.TL1 [7], _26397_);
  dff (\oc8051_golden_model_1.TMOD [0], _28949_);
  dff (\oc8051_golden_model_1.TMOD [1], _28950_);
  dff (\oc8051_golden_model_1.TMOD [2], _28951_);
  dff (\oc8051_golden_model_1.TMOD [3], _28952_);
  dff (\oc8051_golden_model_1.TMOD [4], _28953_);
  dff (\oc8051_golden_model_1.TMOD [5], _28954_);
  dff (\oc8051_golden_model_1.TMOD [6], _28955_);
  dff (\oc8051_golden_model_1.TMOD [7], _26395_);
  dff (\oc8051_golden_model_1.PC [0], _28958_);
  dff (\oc8051_golden_model_1.PC [1], _28959_);
  dff (\oc8051_golden_model_1.PC [2], _28960_);
  dff (\oc8051_golden_model_1.PC [3], _28961_);
  dff (\oc8051_golden_model_1.PC [4], _28964_);
  dff (\oc8051_golden_model_1.PC [5], _28965_);
  dff (\oc8051_golden_model_1.PC [6], _28966_);
  dff (\oc8051_golden_model_1.PC [7], _28967_);
  dff (\oc8051_golden_model_1.PC [8], _28968_);
  dff (\oc8051_golden_model_1.PC [9], _28969_);
  dff (\oc8051_golden_model_1.PC [10], _28970_);
  dff (\oc8051_golden_model_1.PC [11], _28971_);
  dff (\oc8051_golden_model_1.PC [12], _28972_);
  dff (\oc8051_golden_model_1.PC [13], _28973_);
  dff (\oc8051_golden_model_1.PC [14], _28974_);
  dff (\oc8051_golden_model_1.PC [15], _26394_);
  dff (\oc8051_golden_model_1.P0INREG [0], _28975_);
  dff (\oc8051_golden_model_1.P0INREG [1], _28976_);
  dff (\oc8051_golden_model_1.P0INREG [2], _28979_);
  dff (\oc8051_golden_model_1.P0INREG [3], _28980_);
  dff (\oc8051_golden_model_1.P0INREG [4], _28981_);
  dff (\oc8051_golden_model_1.P0INREG [5], _28982_);
  dff (\oc8051_golden_model_1.P0INREG [6], _28983_);
  dff (\oc8051_golden_model_1.P0INREG [7], _26392_);
  dff (\oc8051_golden_model_1.P1INREG [0], _28986_);
  dff (\oc8051_golden_model_1.P1INREG [1], _28987_);
  dff (\oc8051_golden_model_1.P1INREG [2], _28988_);
  dff (\oc8051_golden_model_1.P1INREG [3], _28989_);
  dff (\oc8051_golden_model_1.P1INREG [4], _28990_);
  dff (\oc8051_golden_model_1.P1INREG [5], _28991_);
  dff (\oc8051_golden_model_1.P1INREG [6], _28992_);
  dff (\oc8051_golden_model_1.P1INREG [7], _26391_);
  dff (\oc8051_golden_model_1.P2INREG [0], _28993_);
  dff (\oc8051_golden_model_1.P2INREG [1], _28994_);
  dff (\oc8051_golden_model_1.P2INREG [2], _28995_);
  dff (\oc8051_golden_model_1.P2INREG [3], _28996_);
  dff (\oc8051_golden_model_1.P2INREG [4], _28999_);
  dff (\oc8051_golden_model_1.P2INREG [5], _29000_);
  dff (\oc8051_golden_model_1.P2INREG [6], _29001_);
  dff (\oc8051_golden_model_1.P2INREG [7], _26390_);
  dff (\oc8051_golden_model_1.P3INREG [0], _29004_);
  dff (\oc8051_golden_model_1.P3INREG [1], _29005_);
  dff (\oc8051_golden_model_1.P3INREG [2], _29006_);
  dff (\oc8051_golden_model_1.P3INREG [3], _29007_);
  dff (\oc8051_golden_model_1.P3INREG [4], _29008_);
  dff (\oc8051_golden_model_1.P3INREG [5], _29009_);
  dff (\oc8051_golden_model_1.P3INREG [6], _29010_);
  dff (\oc8051_golden_model_1.P3INREG [7], _26389_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _01036_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _01039_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _01042_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _01044_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _01047_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _01050_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _01053_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _00906_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _01056_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _01059_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _01062_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _01065_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _01068_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _01071_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _01074_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _00910_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _01077_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _01080_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _01083_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _01086_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _01089_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _01091_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _01094_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _00914_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _12189_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _12191_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _12105_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _12194_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _12197_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _12108_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _12200_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _12111_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _12203_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _12206_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _12209_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _12212_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _12215_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _12218_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _12221_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _12114_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _12117_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _25347_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _12120_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _25348_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _12123_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _25349_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _25350_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _12126_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _25351_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _25352_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _12129_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _25353_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _12132_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _25354_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _25355_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _25356_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _12135_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _25358_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _12138_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _12141_);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _08171_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _03604_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _03606_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _03608_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _03610_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _03612_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _03614_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _03616_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _03618_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _03620_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _03622_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _03624_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _03626_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _03628_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _03630_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _03632_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _02749_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _03664_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _03666_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _03668_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _03670_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _03672_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _03674_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _03676_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _03678_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _03680_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _03682_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _03684_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _03686_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _03688_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _03690_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _03692_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _02753_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _05565_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _05567_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _05569_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _05571_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _05573_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _05575_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _05577_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _05579_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _05581_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _05583_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _05585_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _05587_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _05589_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _05591_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _05593_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _05595_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _05597_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _05599_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _05601_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _05603_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _05605_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _05607_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _05609_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _05611_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _05613_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _05615_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _05617_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _05619_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _05621_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _05623_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _05625_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _03202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _03131_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _05628_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _05631_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _05634_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _05636_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _03138_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _05639_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _05642_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _05645_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _05648_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _05651_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _05654_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _05657_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _03142_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _05659_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _05661_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _05663_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _05665_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _05667_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _05669_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _05671_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _03145_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _05673_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _05675_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _05677_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _05679_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _05681_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _05683_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _05685_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _03148_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _03151_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _03155_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _05687_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _05689_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _05691_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _05693_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _05695_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _05697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _05699_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _03158_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _05701_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _05703_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _05705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _05707_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _05709_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _05711_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _05713_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _05715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _05717_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _05719_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _05721_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _05723_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _05725_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _05727_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _05729_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _03161_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _05731_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _05733_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _05735_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _05737_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _05739_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _05741_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _05743_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _05745_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _05747_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _05749_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _05751_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _05753_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _05755_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _05757_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _05759_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03164_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _03169_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _03175_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _03172_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _05761_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _05763_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _05765_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _05767_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _05769_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _05771_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _05773_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _03178_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _05775_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _05777_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _03180_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _05779_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _05781_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _05783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _05785_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _05787_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _05789_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _05791_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _03182_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _05793_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _05795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _05797_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _05799_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _05801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _05803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _05805_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _03185_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _03188_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _05807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _05809_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _05811_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _05813_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _05815_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _05817_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _05819_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03190_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _03193_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _03196_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _05821_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _05823_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _05825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _03199_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _05827_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _05829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _05831_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _05833_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _05835_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _05837_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _05839_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _05841_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _05843_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _05845_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _05847_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _05849_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _05851_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _05853_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _05855_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _05857_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _05859_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _05861_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _05863_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _05865_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _05867_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _05869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _05871_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _05873_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _05875_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _05877_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _05879_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _05881_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _05882_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _05884_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _05886_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _03204_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _05888_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _05890_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _05892_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _05894_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _05896_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _05898_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _05900_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _03206_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _03208_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _03210_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _05902_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _05904_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _05906_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _05908_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _05910_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _05912_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _05914_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _05916_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _05918_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _05920_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _05922_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _05924_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _05926_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _05928_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _05930_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _03212_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _03214_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _03216_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _03218_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _05932_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _05934_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _05936_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _05938_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _05940_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _05942_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _05944_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _05946_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _05948_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _05950_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _05952_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _05954_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _05956_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _05958_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _05960_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _03220_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _03222_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _08268_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _08429_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _08431_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _08433_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _08435_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _08437_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _08439_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _08441_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _08271_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _08274_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _08443_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _08445_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _08277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _28438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _28444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _28450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _28456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _28462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _28467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _28473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _28476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _28518_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _28522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _28526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _28530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _28534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _28538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _28542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _28545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _28484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _28488_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _28492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _28496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _28500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _28504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _28507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _28510_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _28585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _28589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _28593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _28597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _28600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _28604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _28608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _28611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _28551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _28554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _28558_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _28562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _28566_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _28570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _28574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _28577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _28743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _28744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _28746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _28750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _28754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _28758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _28762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _28772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _28713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _28717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _28721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _28725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _28729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _28733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _28736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _28739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _28679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _28683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _28687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _28690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _28694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _28698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _28702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _28705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _28647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _28651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _28655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _28659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _28663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _28667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _28671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _28674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _28616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _28620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _28624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _28628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _28632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _28636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _28640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _28643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _29118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _29122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _29126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _29130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _29134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _29138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _29142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _28150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _29086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _29090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _29094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _29098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _29102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _29106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _29110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _29113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _29057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _29061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _29065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _29069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _29072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _29074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _29078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _29081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _29025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _29029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _29033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _29037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _29041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _29045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _29049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _29052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _28921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _28939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _28957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _28978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _28998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _29012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _29016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _29019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _28791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _28807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _28820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _28838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _28849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _28866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _28885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _28895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _00044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _00046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _00048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _00049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _00051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _00053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _00055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _28138_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _01506_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _01508_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _02181_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _02183_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _02185_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _02187_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _02189_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _02191_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _02193_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _01510_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _01513_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _08829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _08840_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _08851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _08862_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _08873_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _08884_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _08895_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _07125_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _24640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _24650_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _24660_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _24671_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _24681_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _24692_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _24702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _05301_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _29419_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _29430_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _29441_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _29452_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _29463_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _29474_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _29485_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _28181_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _29496_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _29507_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _29518_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _29529_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _29540_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _29551_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _29562_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _28202_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _27053_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _27993_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _27995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _27997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _27999_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _28001_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _28003_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _28005_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _27056_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _28007_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _27058_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _27061_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _28009_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _28011_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _27064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _28013_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _28015_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _27066_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _28017_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _27068_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _28019_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _27070_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _27105_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _27107_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _27109_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _27111_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _28021_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _28023_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _28025_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _27113_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _28027_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _28029_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _28031_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _28033_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _28035_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _28037_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _28039_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _27115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _28041_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _28043_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _28045_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _28047_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _28049_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _28051_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _28053_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _27117_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _26462_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _26464_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _26466_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _26468_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _26469_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _26471_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _26473_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _19326_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _26474_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _26476_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _26478_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _26480_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _26482_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _26483_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _26485_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _19349_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _26487_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _26489_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _26490_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _26492_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _26494_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _26496_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _26497_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _19372_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _26499_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _26501_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _26503_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _26504_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _26506_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _26508_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _26510_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _19395_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _06362_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _06373_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _06384_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _06394_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _06405_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _06416_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _01583_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _26240_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _26249_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _26257_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _26266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _26274_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _26283_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _26291_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _25196_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _25177_);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in , ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in , ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], 1'b0);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], 1'b0);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.desAc , ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_sfr1.desOv , ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [8], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [9], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [10], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [11], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [12], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [13], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [14], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [15], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_data_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_comp1.des [0], ABINPUT[27]);
  buf(\oc8051_top_1.oc8051_comp1.des [1], ABINPUT[28]);
  buf(\oc8051_top_1.oc8051_comp1.des [2], ABINPUT[29]);
  buf(\oc8051_top_1.oc8051_comp1.des [3], ABINPUT[30]);
  buf(\oc8051_top_1.oc8051_comp1.des [4], ABINPUT[31]);
  buf(\oc8051_top_1.oc8051_comp1.des [5], ABINPUT[32]);
  buf(\oc8051_top_1.oc8051_comp1.des [6], ABINPUT[33]);
  buf(\oc8051_top_1.oc8051_comp1.des [7], ABINPUT[34]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.PSW_next [0], ABINPUT008[0]);
  buf(\oc8051_golden_model_1.PSW_next [1], ABINPUT008[1]);
  buf(\oc8051_golden_model_1.PSW_next [2], ABINPUT008[2]);
  buf(\oc8051_golden_model_1.PSW_next [3], ABINPUT008[3]);
  buf(\oc8051_golden_model_1.PSW_next [4], ABINPUT008[4]);
  buf(\oc8051_golden_model_1.PSW_next [5], ABINPUT008[5]);
  buf(\oc8051_golden_model_1.PSW_next [6], ABINPUT008[6]);
  buf(\oc8051_golden_model_1.PSW_next [7], ABINPUT008[7]);
  buf(\oc8051_golden_model_1.ABINPUT007 [0], ABINPUT008[0]);
  buf(\oc8051_golden_model_1.ABINPUT007 [1], ABINPUT008[1]);
  buf(\oc8051_golden_model_1.ABINPUT007 [2], ABINPUT008[2]);
  buf(\oc8051_golden_model_1.ABINPUT007 [3], ABINPUT008[3]);
  buf(\oc8051_golden_model_1.ABINPUT007 [4], ABINPUT008[4]);
  buf(\oc8051_golden_model_1.ABINPUT007 [5], ABINPUT008[5]);
  buf(\oc8051_golden_model_1.ABINPUT007 [6], ABINPUT008[6]);
  buf(\oc8051_golden_model_1.ABINPUT007 [7], ABINPUT008[7]);
  buf(\oc8051_golden_model_1.P2_next [0], ABINPUT006[0]);
  buf(\oc8051_golden_model_1.P2_next [1], ABINPUT006[1]);
  buf(\oc8051_golden_model_1.P2_next [2], ABINPUT006[2]);
  buf(\oc8051_golden_model_1.P2_next [3], ABINPUT006[3]);
  buf(\oc8051_golden_model_1.P2_next [4], ABINPUT006[4]);
  buf(\oc8051_golden_model_1.P2_next [5], ABINPUT006[5]);
  buf(\oc8051_golden_model_1.P2_next [6], ABINPUT006[6]);
  buf(\oc8051_golden_model_1.P2_next [7], ABINPUT006[7]);
  buf(\oc8051_golden_model_1.ABINPUT005 [0], ABINPUT006[0]);
  buf(\oc8051_golden_model_1.ABINPUT005 [1], ABINPUT006[1]);
  buf(\oc8051_golden_model_1.ABINPUT005 [2], ABINPUT006[2]);
  buf(\oc8051_golden_model_1.ABINPUT005 [3], ABINPUT006[3]);
  buf(\oc8051_golden_model_1.ABINPUT005 [4], ABINPUT006[4]);
  buf(\oc8051_golden_model_1.ABINPUT005 [5], ABINPUT006[5]);
  buf(\oc8051_golden_model_1.ABINPUT005 [6], ABINPUT006[6]);
  buf(\oc8051_golden_model_1.ABINPUT005 [7], ABINPUT006[7]);
  buf(\oc8051_golden_model_1.P0_next [0], ABINPUT004[0]);
  buf(\oc8051_golden_model_1.P0_next [1], ABINPUT004[1]);
  buf(\oc8051_golden_model_1.P0_next [2], ABINPUT004[2]);
  buf(\oc8051_golden_model_1.P0_next [3], ABINPUT004[3]);
  buf(\oc8051_golden_model_1.P0_next [4], ABINPUT004[4]);
  buf(\oc8051_golden_model_1.P0_next [5], ABINPUT004[5]);
  buf(\oc8051_golden_model_1.P0_next [6], ABINPUT004[6]);
  buf(\oc8051_golden_model_1.P0_next [7], ABINPUT004[7]);
  buf(\oc8051_golden_model_1.ABINPUT003 [0], ABINPUT004[0]);
  buf(\oc8051_golden_model_1.ABINPUT003 [1], ABINPUT004[1]);
  buf(\oc8051_golden_model_1.ABINPUT003 [2], ABINPUT004[2]);
  buf(\oc8051_golden_model_1.ABINPUT003 [3], ABINPUT004[3]);
  buf(\oc8051_golden_model_1.ABINPUT003 [4], ABINPUT004[4]);
  buf(\oc8051_golden_model_1.ABINPUT003 [5], ABINPUT004[5]);
  buf(\oc8051_golden_model_1.ABINPUT003 [6], ABINPUT004[6]);
  buf(\oc8051_golden_model_1.ABINPUT003 [7], ABINPUT004[7]);
  buf(\oc8051_golden_model_1.DPL_next [0], ABINPUT002[0]);
  buf(\oc8051_golden_model_1.DPL_next [1], ABINPUT002[1]);
  buf(\oc8051_golden_model_1.DPL_next [2], ABINPUT002[2]);
  buf(\oc8051_golden_model_1.DPL_next [3], ABINPUT002[3]);
  buf(\oc8051_golden_model_1.DPL_next [4], ABINPUT002[4]);
  buf(\oc8051_golden_model_1.DPL_next [5], ABINPUT002[5]);
  buf(\oc8051_golden_model_1.DPL_next [6], ABINPUT002[6]);
  buf(\oc8051_golden_model_1.DPL_next [7], ABINPUT002[7]);
  buf(\oc8051_golden_model_1.ABINPUT001 [0], ABINPUT002[0]);
  buf(\oc8051_golden_model_1.ABINPUT001 [1], ABINPUT002[1]);
  buf(\oc8051_golden_model_1.ABINPUT001 [2], ABINPUT002[2]);
  buf(\oc8051_golden_model_1.ABINPUT001 [3], ABINPUT002[3]);
  buf(\oc8051_golden_model_1.ABINPUT001 [4], ABINPUT002[4]);
  buf(\oc8051_golden_model_1.ABINPUT001 [5], ABINPUT002[5]);
  buf(\oc8051_golden_model_1.ABINPUT001 [6], ABINPUT002[6]);
  buf(\oc8051_golden_model_1.ABINPUT001 [7], ABINPUT002[7]);
  buf(\oc8051_golden_model_1.ACC_next [0], ABINPUT000[0]);
  buf(\oc8051_golden_model_1.ACC_next [1], ABINPUT000[1]);
  buf(\oc8051_golden_model_1.ACC_next [2], ABINPUT000[2]);
  buf(\oc8051_golden_model_1.ACC_next [3], ABINPUT000[3]);
  buf(\oc8051_golden_model_1.ACC_next [4], ABINPUT000[4]);
  buf(\oc8051_golden_model_1.ACC_next [5], ABINPUT000[5]);
  buf(\oc8051_golden_model_1.ACC_next [6], ABINPUT000[6]);
  buf(\oc8051_golden_model_1.ACC_next [7], ABINPUT000[7]);
  buf(\oc8051_golden_model_1.ABINPUT [0], ABINPUT000[0]);
  buf(\oc8051_golden_model_1.ABINPUT [1], ABINPUT000[1]);
  buf(\oc8051_golden_model_1.ABINPUT [2], ABINPUT000[2]);
  buf(\oc8051_golden_model_1.ABINPUT [3], ABINPUT000[3]);
  buf(\oc8051_golden_model_1.ABINPUT [4], ABINPUT000[4]);
  buf(\oc8051_golden_model_1.ABINPUT [5], ABINPUT000[5]);
  buf(\oc8051_golden_model_1.ABINPUT [6], ABINPUT000[6]);
  buf(\oc8051_golden_model_1.ABINPUT [7], ABINPUT000[7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e6 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.ACC_e6 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.ACC_e6 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.ACC_e6 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.ACC_e6 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.ACC_e6 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.ACC_e6 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.ACC_e6 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.ACC_e7 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.ACC_e7 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.ACC_e7 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.ACC_e7 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.ACC_e7 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.ACC_e7 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.ACC_e7 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.ACC_e7 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n2854 [0], \oc8051_golden_model_1.PSW_d4 [0]);
  buf(\oc8051_golden_model_1.n2854 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2854 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2854 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2854 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2854 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2854 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2854 [7], \oc8051_golden_model_1.PSW_d4 [7]);
  buf(\oc8051_golden_model_1.n2858 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n2858 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n2858 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n2858 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n2858 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2858 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2858 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2858 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2859 [0], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n2859 [1], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n2859 [2], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n2859 [3], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n2860 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2860 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2860 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2860 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2860 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n2860 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n2860 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n2860 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n2861 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2862 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2863 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2864 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2865 , \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n2866 , \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n2441 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2441 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2867 , \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n2868 , \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.IRAM_full [0], ABINPUT009[0]);
  buf(\oc8051_golden_model_1.IRAM_full [1], ABINPUT009[1]);
  buf(\oc8051_golden_model_1.IRAM_full [2], ABINPUT009[2]);
  buf(\oc8051_golden_model_1.IRAM_full [3], ABINPUT009[3]);
  buf(\oc8051_golden_model_1.IRAM_full [4], ABINPUT009[4]);
  buf(\oc8051_golden_model_1.IRAM_full [5], ABINPUT009[5]);
  buf(\oc8051_golden_model_1.IRAM_full [6], ABINPUT009[6]);
  buf(\oc8051_golden_model_1.IRAM_full [7], ABINPUT009[7]);
  buf(\oc8051_golden_model_1.IRAM_full [8], ABINPUT009[8]);
  buf(\oc8051_golden_model_1.IRAM_full [9], ABINPUT009[9]);
  buf(\oc8051_golden_model_1.IRAM_full [10], ABINPUT009[10]);
  buf(\oc8051_golden_model_1.IRAM_full [11], ABINPUT009[11]);
  buf(\oc8051_golden_model_1.IRAM_full [12], ABINPUT009[12]);
  buf(\oc8051_golden_model_1.IRAM_full [13], ABINPUT009[13]);
  buf(\oc8051_golden_model_1.IRAM_full [14], ABINPUT009[14]);
  buf(\oc8051_golden_model_1.IRAM_full [15], ABINPUT009[15]);
  buf(\oc8051_golden_model_1.IRAM_full [16], ABINPUT009[16]);
  buf(\oc8051_golden_model_1.IRAM_full [17], ABINPUT009[17]);
  buf(\oc8051_golden_model_1.IRAM_full [18], ABINPUT009[18]);
  buf(\oc8051_golden_model_1.IRAM_full [19], ABINPUT009[19]);
  buf(\oc8051_golden_model_1.IRAM_full [20], ABINPUT009[20]);
  buf(\oc8051_golden_model_1.IRAM_full [21], ABINPUT009[21]);
  buf(\oc8051_golden_model_1.IRAM_full [22], ABINPUT009[22]);
  buf(\oc8051_golden_model_1.IRAM_full [23], ABINPUT009[23]);
  buf(\oc8051_golden_model_1.IRAM_full [24], ABINPUT009[24]);
  buf(\oc8051_golden_model_1.IRAM_full [25], ABINPUT009[25]);
  buf(\oc8051_golden_model_1.IRAM_full [26], ABINPUT009[26]);
  buf(\oc8051_golden_model_1.IRAM_full [27], ABINPUT009[27]);
  buf(\oc8051_golden_model_1.IRAM_full [28], ABINPUT009[28]);
  buf(\oc8051_golden_model_1.IRAM_full [29], ABINPUT009[29]);
  buf(\oc8051_golden_model_1.IRAM_full [30], ABINPUT009[30]);
  buf(\oc8051_golden_model_1.IRAM_full [31], ABINPUT009[31]);
  buf(\oc8051_golden_model_1.IRAM_full [32], ABINPUT009[32]);
  buf(\oc8051_golden_model_1.IRAM_full [33], ABINPUT009[33]);
  buf(\oc8051_golden_model_1.IRAM_full [34], ABINPUT009[34]);
  buf(\oc8051_golden_model_1.IRAM_full [35], ABINPUT009[35]);
  buf(\oc8051_golden_model_1.IRAM_full [36], ABINPUT009[36]);
  buf(\oc8051_golden_model_1.IRAM_full [37], ABINPUT009[37]);
  buf(\oc8051_golden_model_1.IRAM_full [38], ABINPUT009[38]);
  buf(\oc8051_golden_model_1.IRAM_full [39], ABINPUT009[39]);
  buf(\oc8051_golden_model_1.IRAM_full [40], ABINPUT009[40]);
  buf(\oc8051_golden_model_1.IRAM_full [41], ABINPUT009[41]);
  buf(\oc8051_golden_model_1.IRAM_full [42], ABINPUT009[42]);
  buf(\oc8051_golden_model_1.IRAM_full [43], ABINPUT009[43]);
  buf(\oc8051_golden_model_1.IRAM_full [44], ABINPUT009[44]);
  buf(\oc8051_golden_model_1.IRAM_full [45], ABINPUT009[45]);
  buf(\oc8051_golden_model_1.IRAM_full [46], ABINPUT009[46]);
  buf(\oc8051_golden_model_1.IRAM_full [47], ABINPUT009[47]);
  buf(\oc8051_golden_model_1.IRAM_full [48], ABINPUT009[48]);
  buf(\oc8051_golden_model_1.IRAM_full [49], ABINPUT009[49]);
  buf(\oc8051_golden_model_1.IRAM_full [50], ABINPUT009[50]);
  buf(\oc8051_golden_model_1.IRAM_full [51], ABINPUT009[51]);
  buf(\oc8051_golden_model_1.IRAM_full [52], ABINPUT009[52]);
  buf(\oc8051_golden_model_1.IRAM_full [53], ABINPUT009[53]);
  buf(\oc8051_golden_model_1.IRAM_full [54], ABINPUT009[54]);
  buf(\oc8051_golden_model_1.IRAM_full [55], ABINPUT009[55]);
  buf(\oc8051_golden_model_1.IRAM_full [56], ABINPUT009[56]);
  buf(\oc8051_golden_model_1.IRAM_full [57], ABINPUT009[57]);
  buf(\oc8051_golden_model_1.IRAM_full [58], ABINPUT009[58]);
  buf(\oc8051_golden_model_1.IRAM_full [59], ABINPUT009[59]);
  buf(\oc8051_golden_model_1.IRAM_full [60], ABINPUT009[60]);
  buf(\oc8051_golden_model_1.IRAM_full [61], ABINPUT009[61]);
  buf(\oc8051_golden_model_1.IRAM_full [62], ABINPUT009[62]);
  buf(\oc8051_golden_model_1.IRAM_full [63], ABINPUT009[63]);
  buf(\oc8051_golden_model_1.IRAM_full [64], ABINPUT009[64]);
  buf(\oc8051_golden_model_1.IRAM_full [65], ABINPUT009[65]);
  buf(\oc8051_golden_model_1.IRAM_full [66], ABINPUT009[66]);
  buf(\oc8051_golden_model_1.IRAM_full [67], ABINPUT009[67]);
  buf(\oc8051_golden_model_1.IRAM_full [68], ABINPUT009[68]);
  buf(\oc8051_golden_model_1.IRAM_full [69], ABINPUT009[69]);
  buf(\oc8051_golden_model_1.IRAM_full [70], ABINPUT009[70]);
  buf(\oc8051_golden_model_1.IRAM_full [71], ABINPUT009[71]);
  buf(\oc8051_golden_model_1.IRAM_full [72], ABINPUT009[72]);
  buf(\oc8051_golden_model_1.IRAM_full [73], ABINPUT009[73]);
  buf(\oc8051_golden_model_1.IRAM_full [74], ABINPUT009[74]);
  buf(\oc8051_golden_model_1.IRAM_full [75], ABINPUT009[75]);
  buf(\oc8051_golden_model_1.IRAM_full [76], ABINPUT009[76]);
  buf(\oc8051_golden_model_1.IRAM_full [77], ABINPUT009[77]);
  buf(\oc8051_golden_model_1.IRAM_full [78], ABINPUT009[78]);
  buf(\oc8051_golden_model_1.IRAM_full [79], ABINPUT009[79]);
  buf(\oc8051_golden_model_1.IRAM_full [80], ABINPUT009[80]);
  buf(\oc8051_golden_model_1.IRAM_full [81], ABINPUT009[81]);
  buf(\oc8051_golden_model_1.IRAM_full [82], ABINPUT009[82]);
  buf(\oc8051_golden_model_1.IRAM_full [83], ABINPUT009[83]);
  buf(\oc8051_golden_model_1.IRAM_full [84], ABINPUT009[84]);
  buf(\oc8051_golden_model_1.IRAM_full [85], ABINPUT009[85]);
  buf(\oc8051_golden_model_1.IRAM_full [86], ABINPUT009[86]);
  buf(\oc8051_golden_model_1.IRAM_full [87], ABINPUT009[87]);
  buf(\oc8051_golden_model_1.IRAM_full [88], ABINPUT009[88]);
  buf(\oc8051_golden_model_1.IRAM_full [89], ABINPUT009[89]);
  buf(\oc8051_golden_model_1.IRAM_full [90], ABINPUT009[90]);
  buf(\oc8051_golden_model_1.IRAM_full [91], ABINPUT009[91]);
  buf(\oc8051_golden_model_1.IRAM_full [92], ABINPUT009[92]);
  buf(\oc8051_golden_model_1.IRAM_full [93], ABINPUT009[93]);
  buf(\oc8051_golden_model_1.IRAM_full [94], ABINPUT009[94]);
  buf(\oc8051_golden_model_1.IRAM_full [95], ABINPUT009[95]);
  buf(\oc8051_golden_model_1.IRAM_full [96], ABINPUT009[96]);
  buf(\oc8051_golden_model_1.IRAM_full [97], ABINPUT009[97]);
  buf(\oc8051_golden_model_1.IRAM_full [98], ABINPUT009[98]);
  buf(\oc8051_golden_model_1.IRAM_full [99], ABINPUT009[99]);
  buf(\oc8051_golden_model_1.IRAM_full [100], ABINPUT009[100]);
  buf(\oc8051_golden_model_1.IRAM_full [101], ABINPUT009[101]);
  buf(\oc8051_golden_model_1.IRAM_full [102], ABINPUT009[102]);
  buf(\oc8051_golden_model_1.IRAM_full [103], ABINPUT009[103]);
  buf(\oc8051_golden_model_1.IRAM_full [104], ABINPUT009[104]);
  buf(\oc8051_golden_model_1.IRAM_full [105], ABINPUT009[105]);
  buf(\oc8051_golden_model_1.IRAM_full [106], ABINPUT009[106]);
  buf(\oc8051_golden_model_1.IRAM_full [107], ABINPUT009[107]);
  buf(\oc8051_golden_model_1.IRAM_full [108], ABINPUT009[108]);
  buf(\oc8051_golden_model_1.IRAM_full [109], ABINPUT009[109]);
  buf(\oc8051_golden_model_1.IRAM_full [110], ABINPUT009[110]);
  buf(\oc8051_golden_model_1.IRAM_full [111], ABINPUT009[111]);
  buf(\oc8051_golden_model_1.IRAM_full [112], ABINPUT009[112]);
  buf(\oc8051_golden_model_1.IRAM_full [113], ABINPUT009[113]);
  buf(\oc8051_golden_model_1.IRAM_full [114], ABINPUT009[114]);
  buf(\oc8051_golden_model_1.IRAM_full [115], ABINPUT009[115]);
  buf(\oc8051_golden_model_1.IRAM_full [116], ABINPUT009[116]);
  buf(\oc8051_golden_model_1.IRAM_full [117], ABINPUT009[117]);
  buf(\oc8051_golden_model_1.IRAM_full [118], ABINPUT009[118]);
  buf(\oc8051_golden_model_1.IRAM_full [119], ABINPUT009[119]);
  buf(\oc8051_golden_model_1.IRAM_full [120], ABINPUT009[120]);
  buf(\oc8051_golden_model_1.IRAM_full [121], ABINPUT009[121]);
  buf(\oc8051_golden_model_1.IRAM_full [122], ABINPUT009[122]);
  buf(\oc8051_golden_model_1.IRAM_full [123], ABINPUT009[123]);
  buf(\oc8051_golden_model_1.IRAM_full [124], ABINPUT009[124]);
  buf(\oc8051_golden_model_1.IRAM_full [125], ABINPUT009[125]);
  buf(\oc8051_golden_model_1.IRAM_full [126], ABINPUT009[126]);
  buf(\oc8051_golden_model_1.IRAM_full [127], ABINPUT009[127]);
  buf(\oc8051_golden_model_1.ABINPUT008 [0], ABINPUT009[0]);
  buf(\oc8051_golden_model_1.ABINPUT008 [1], ABINPUT009[1]);
  buf(\oc8051_golden_model_1.ABINPUT008 [2], ABINPUT009[2]);
  buf(\oc8051_golden_model_1.ABINPUT008 [3], ABINPUT009[3]);
  buf(\oc8051_golden_model_1.ABINPUT008 [4], ABINPUT009[4]);
  buf(\oc8051_golden_model_1.ABINPUT008 [5], ABINPUT009[5]);
  buf(\oc8051_golden_model_1.ABINPUT008 [6], ABINPUT009[6]);
  buf(\oc8051_golden_model_1.ABINPUT008 [7], ABINPUT009[7]);
  buf(\oc8051_golden_model_1.ABINPUT008 [8], ABINPUT009[8]);
  buf(\oc8051_golden_model_1.ABINPUT008 [9], ABINPUT009[9]);
  buf(\oc8051_golden_model_1.ABINPUT008 [10], ABINPUT009[10]);
  buf(\oc8051_golden_model_1.ABINPUT008 [11], ABINPUT009[11]);
  buf(\oc8051_golden_model_1.ABINPUT008 [12], ABINPUT009[12]);
  buf(\oc8051_golden_model_1.ABINPUT008 [13], ABINPUT009[13]);
  buf(\oc8051_golden_model_1.ABINPUT008 [14], ABINPUT009[14]);
  buf(\oc8051_golden_model_1.ABINPUT008 [15], ABINPUT009[15]);
  buf(\oc8051_golden_model_1.ABINPUT008 [16], ABINPUT009[16]);
  buf(\oc8051_golden_model_1.ABINPUT008 [17], ABINPUT009[17]);
  buf(\oc8051_golden_model_1.ABINPUT008 [18], ABINPUT009[18]);
  buf(\oc8051_golden_model_1.ABINPUT008 [19], ABINPUT009[19]);
  buf(\oc8051_golden_model_1.ABINPUT008 [20], ABINPUT009[20]);
  buf(\oc8051_golden_model_1.ABINPUT008 [21], ABINPUT009[21]);
  buf(\oc8051_golden_model_1.ABINPUT008 [22], ABINPUT009[22]);
  buf(\oc8051_golden_model_1.ABINPUT008 [23], ABINPUT009[23]);
  buf(\oc8051_golden_model_1.ABINPUT008 [24], ABINPUT009[24]);
  buf(\oc8051_golden_model_1.ABINPUT008 [25], ABINPUT009[25]);
  buf(\oc8051_golden_model_1.ABINPUT008 [26], ABINPUT009[26]);
  buf(\oc8051_golden_model_1.ABINPUT008 [27], ABINPUT009[27]);
  buf(\oc8051_golden_model_1.ABINPUT008 [28], ABINPUT009[28]);
  buf(\oc8051_golden_model_1.ABINPUT008 [29], ABINPUT009[29]);
  buf(\oc8051_golden_model_1.ABINPUT008 [30], ABINPUT009[30]);
  buf(\oc8051_golden_model_1.ABINPUT008 [31], ABINPUT009[31]);
  buf(\oc8051_golden_model_1.ABINPUT008 [32], ABINPUT009[32]);
  buf(\oc8051_golden_model_1.ABINPUT008 [33], ABINPUT009[33]);
  buf(\oc8051_golden_model_1.ABINPUT008 [34], ABINPUT009[34]);
  buf(\oc8051_golden_model_1.ABINPUT008 [35], ABINPUT009[35]);
  buf(\oc8051_golden_model_1.ABINPUT008 [36], ABINPUT009[36]);
  buf(\oc8051_golden_model_1.ABINPUT008 [37], ABINPUT009[37]);
  buf(\oc8051_golden_model_1.ABINPUT008 [38], ABINPUT009[38]);
  buf(\oc8051_golden_model_1.ABINPUT008 [39], ABINPUT009[39]);
  buf(\oc8051_golden_model_1.ABINPUT008 [40], ABINPUT009[40]);
  buf(\oc8051_golden_model_1.ABINPUT008 [41], ABINPUT009[41]);
  buf(\oc8051_golden_model_1.ABINPUT008 [42], ABINPUT009[42]);
  buf(\oc8051_golden_model_1.ABINPUT008 [43], ABINPUT009[43]);
  buf(\oc8051_golden_model_1.ABINPUT008 [44], ABINPUT009[44]);
  buf(\oc8051_golden_model_1.ABINPUT008 [45], ABINPUT009[45]);
  buf(\oc8051_golden_model_1.ABINPUT008 [46], ABINPUT009[46]);
  buf(\oc8051_golden_model_1.ABINPUT008 [47], ABINPUT009[47]);
  buf(\oc8051_golden_model_1.ABINPUT008 [48], ABINPUT009[48]);
  buf(\oc8051_golden_model_1.ABINPUT008 [49], ABINPUT009[49]);
  buf(\oc8051_golden_model_1.ABINPUT008 [50], ABINPUT009[50]);
  buf(\oc8051_golden_model_1.ABINPUT008 [51], ABINPUT009[51]);
  buf(\oc8051_golden_model_1.ABINPUT008 [52], ABINPUT009[52]);
  buf(\oc8051_golden_model_1.ABINPUT008 [53], ABINPUT009[53]);
  buf(\oc8051_golden_model_1.ABINPUT008 [54], ABINPUT009[54]);
  buf(\oc8051_golden_model_1.ABINPUT008 [55], ABINPUT009[55]);
  buf(\oc8051_golden_model_1.ABINPUT008 [56], ABINPUT009[56]);
  buf(\oc8051_golden_model_1.ABINPUT008 [57], ABINPUT009[57]);
  buf(\oc8051_golden_model_1.ABINPUT008 [58], ABINPUT009[58]);
  buf(\oc8051_golden_model_1.ABINPUT008 [59], ABINPUT009[59]);
  buf(\oc8051_golden_model_1.ABINPUT008 [60], ABINPUT009[60]);
  buf(\oc8051_golden_model_1.ABINPUT008 [61], ABINPUT009[61]);
  buf(\oc8051_golden_model_1.ABINPUT008 [62], ABINPUT009[62]);
  buf(\oc8051_golden_model_1.ABINPUT008 [63], ABINPUT009[63]);
  buf(\oc8051_golden_model_1.ABINPUT008 [64], ABINPUT009[64]);
  buf(\oc8051_golden_model_1.ABINPUT008 [65], ABINPUT009[65]);
  buf(\oc8051_golden_model_1.ABINPUT008 [66], ABINPUT009[66]);
  buf(\oc8051_golden_model_1.ABINPUT008 [67], ABINPUT009[67]);
  buf(\oc8051_golden_model_1.ABINPUT008 [68], ABINPUT009[68]);
  buf(\oc8051_golden_model_1.ABINPUT008 [69], ABINPUT009[69]);
  buf(\oc8051_golden_model_1.ABINPUT008 [70], ABINPUT009[70]);
  buf(\oc8051_golden_model_1.ABINPUT008 [71], ABINPUT009[71]);
  buf(\oc8051_golden_model_1.ABINPUT008 [72], ABINPUT009[72]);
  buf(\oc8051_golden_model_1.ABINPUT008 [73], ABINPUT009[73]);
  buf(\oc8051_golden_model_1.ABINPUT008 [74], ABINPUT009[74]);
  buf(\oc8051_golden_model_1.ABINPUT008 [75], ABINPUT009[75]);
  buf(\oc8051_golden_model_1.ABINPUT008 [76], ABINPUT009[76]);
  buf(\oc8051_golden_model_1.ABINPUT008 [77], ABINPUT009[77]);
  buf(\oc8051_golden_model_1.ABINPUT008 [78], ABINPUT009[78]);
  buf(\oc8051_golden_model_1.ABINPUT008 [79], ABINPUT009[79]);
  buf(\oc8051_golden_model_1.ABINPUT008 [80], ABINPUT009[80]);
  buf(\oc8051_golden_model_1.ABINPUT008 [81], ABINPUT009[81]);
  buf(\oc8051_golden_model_1.ABINPUT008 [82], ABINPUT009[82]);
  buf(\oc8051_golden_model_1.ABINPUT008 [83], ABINPUT009[83]);
  buf(\oc8051_golden_model_1.ABINPUT008 [84], ABINPUT009[84]);
  buf(\oc8051_golden_model_1.ABINPUT008 [85], ABINPUT009[85]);
  buf(\oc8051_golden_model_1.ABINPUT008 [86], ABINPUT009[86]);
  buf(\oc8051_golden_model_1.ABINPUT008 [87], ABINPUT009[87]);
  buf(\oc8051_golden_model_1.ABINPUT008 [88], ABINPUT009[88]);
  buf(\oc8051_golden_model_1.ABINPUT008 [89], ABINPUT009[89]);
  buf(\oc8051_golden_model_1.ABINPUT008 [90], ABINPUT009[90]);
  buf(\oc8051_golden_model_1.ABINPUT008 [91], ABINPUT009[91]);
  buf(\oc8051_golden_model_1.ABINPUT008 [92], ABINPUT009[92]);
  buf(\oc8051_golden_model_1.ABINPUT008 [93], ABINPUT009[93]);
  buf(\oc8051_golden_model_1.ABINPUT008 [94], ABINPUT009[94]);
  buf(\oc8051_golden_model_1.ABINPUT008 [95], ABINPUT009[95]);
  buf(\oc8051_golden_model_1.ABINPUT008 [96], ABINPUT009[96]);
  buf(\oc8051_golden_model_1.ABINPUT008 [97], ABINPUT009[97]);
  buf(\oc8051_golden_model_1.ABINPUT008 [98], ABINPUT009[98]);
  buf(\oc8051_golden_model_1.ABINPUT008 [99], ABINPUT009[99]);
  buf(\oc8051_golden_model_1.ABINPUT008 [100], ABINPUT009[100]);
  buf(\oc8051_golden_model_1.ABINPUT008 [101], ABINPUT009[101]);
  buf(\oc8051_golden_model_1.ABINPUT008 [102], ABINPUT009[102]);
  buf(\oc8051_golden_model_1.ABINPUT008 [103], ABINPUT009[103]);
  buf(\oc8051_golden_model_1.ABINPUT008 [104], ABINPUT009[104]);
  buf(\oc8051_golden_model_1.ABINPUT008 [105], ABINPUT009[105]);
  buf(\oc8051_golden_model_1.ABINPUT008 [106], ABINPUT009[106]);
  buf(\oc8051_golden_model_1.ABINPUT008 [107], ABINPUT009[107]);
  buf(\oc8051_golden_model_1.ABINPUT008 [108], ABINPUT009[108]);
  buf(\oc8051_golden_model_1.ABINPUT008 [109], ABINPUT009[109]);
  buf(\oc8051_golden_model_1.ABINPUT008 [110], ABINPUT009[110]);
  buf(\oc8051_golden_model_1.ABINPUT008 [111], ABINPUT009[111]);
  buf(\oc8051_golden_model_1.ABINPUT008 [112], ABINPUT009[112]);
  buf(\oc8051_golden_model_1.ABINPUT008 [113], ABINPUT009[113]);
  buf(\oc8051_golden_model_1.ABINPUT008 [114], ABINPUT009[114]);
  buf(\oc8051_golden_model_1.ABINPUT008 [115], ABINPUT009[115]);
  buf(\oc8051_golden_model_1.ABINPUT008 [116], ABINPUT009[116]);
  buf(\oc8051_golden_model_1.ABINPUT008 [117], ABINPUT009[117]);
  buf(\oc8051_golden_model_1.ABINPUT008 [118], ABINPUT009[118]);
  buf(\oc8051_golden_model_1.ABINPUT008 [119], ABINPUT009[119]);
  buf(\oc8051_golden_model_1.ABINPUT008 [120], ABINPUT009[120]);
  buf(\oc8051_golden_model_1.ABINPUT008 [121], ABINPUT009[121]);
  buf(\oc8051_golden_model_1.ABINPUT008 [122], ABINPUT009[122]);
  buf(\oc8051_golden_model_1.ABINPUT008 [123], ABINPUT009[123]);
  buf(\oc8051_golden_model_1.ABINPUT008 [124], ABINPUT009[124]);
  buf(\oc8051_golden_model_1.ABINPUT008 [125], ABINPUT009[125]);
  buf(\oc8051_golden_model_1.ABINPUT008 [126], ABINPUT009[126]);
  buf(\oc8051_golden_model_1.ABINPUT008 [127], ABINPUT009[127]);
  buf(\oc8051_golden_model_1.P3_next [0], ABINPUT007[0]);
  buf(\oc8051_golden_model_1.P3_next [1], ABINPUT007[1]);
  buf(\oc8051_golden_model_1.P3_next [2], ABINPUT007[2]);
  buf(\oc8051_golden_model_1.P3_next [3], ABINPUT007[3]);
  buf(\oc8051_golden_model_1.P3_next [4], ABINPUT007[4]);
  buf(\oc8051_golden_model_1.P3_next [5], ABINPUT007[5]);
  buf(\oc8051_golden_model_1.P3_next [6], ABINPUT007[6]);
  buf(\oc8051_golden_model_1.P3_next [7], ABINPUT007[7]);
  buf(\oc8051_golden_model_1.ABINPUT006 [0], ABINPUT007[0]);
  buf(\oc8051_golden_model_1.ABINPUT006 [1], ABINPUT007[1]);
  buf(\oc8051_golden_model_1.ABINPUT006 [2], ABINPUT007[2]);
  buf(\oc8051_golden_model_1.ABINPUT006 [3], ABINPUT007[3]);
  buf(\oc8051_golden_model_1.ABINPUT006 [4], ABINPUT007[4]);
  buf(\oc8051_golden_model_1.ABINPUT006 [5], ABINPUT007[5]);
  buf(\oc8051_golden_model_1.ABINPUT006 [6], ABINPUT007[6]);
  buf(\oc8051_golden_model_1.ABINPUT006 [7], ABINPUT007[7]);
  buf(\oc8051_golden_model_1.P1_next [0], ABINPUT005[0]);
  buf(\oc8051_golden_model_1.P1_next [1], ABINPUT005[1]);
  buf(\oc8051_golden_model_1.P1_next [2], ABINPUT005[2]);
  buf(\oc8051_golden_model_1.P1_next [3], ABINPUT005[3]);
  buf(\oc8051_golden_model_1.P1_next [4], ABINPUT005[4]);
  buf(\oc8051_golden_model_1.P1_next [5], ABINPUT005[5]);
  buf(\oc8051_golden_model_1.P1_next [6], ABINPUT005[6]);
  buf(\oc8051_golden_model_1.P1_next [7], ABINPUT005[7]);
  buf(\oc8051_golden_model_1.ABINPUT004 [0], ABINPUT005[0]);
  buf(\oc8051_golden_model_1.ABINPUT004 [1], ABINPUT005[1]);
  buf(\oc8051_golden_model_1.ABINPUT004 [2], ABINPUT005[2]);
  buf(\oc8051_golden_model_1.ABINPUT004 [3], ABINPUT005[3]);
  buf(\oc8051_golden_model_1.ABINPUT004 [4], ABINPUT005[4]);
  buf(\oc8051_golden_model_1.ABINPUT004 [5], ABINPUT005[5]);
  buf(\oc8051_golden_model_1.ABINPUT004 [6], ABINPUT005[6]);
  buf(\oc8051_golden_model_1.ABINPUT004 [7], ABINPUT005[7]);
  buf(\oc8051_golden_model_1.DPH_next [0], ABINPUT003[0]);
  buf(\oc8051_golden_model_1.DPH_next [1], ABINPUT003[1]);
  buf(\oc8051_golden_model_1.DPH_next [2], ABINPUT003[2]);
  buf(\oc8051_golden_model_1.DPH_next [3], ABINPUT003[3]);
  buf(\oc8051_golden_model_1.DPH_next [4], ABINPUT003[4]);
  buf(\oc8051_golden_model_1.DPH_next [5], ABINPUT003[5]);
  buf(\oc8051_golden_model_1.DPH_next [6], ABINPUT003[6]);
  buf(\oc8051_golden_model_1.DPH_next [7], ABINPUT003[7]);
  buf(\oc8051_golden_model_1.ABINPUT002 [0], ABINPUT003[0]);
  buf(\oc8051_golden_model_1.ABINPUT002 [1], ABINPUT003[1]);
  buf(\oc8051_golden_model_1.ABINPUT002 [2], ABINPUT003[2]);
  buf(\oc8051_golden_model_1.ABINPUT002 [3], ABINPUT003[3]);
  buf(\oc8051_golden_model_1.ABINPUT002 [4], ABINPUT003[4]);
  buf(\oc8051_golden_model_1.ABINPUT002 [5], ABINPUT003[5]);
  buf(\oc8051_golden_model_1.ABINPUT002 [6], ABINPUT003[6]);
  buf(\oc8051_golden_model_1.ABINPUT002 [7], ABINPUT003[7]);
  buf(\oc8051_golden_model_1.B_next [0], ABINPUT001[0]);
  buf(\oc8051_golden_model_1.B_next [1], ABINPUT001[1]);
  buf(\oc8051_golden_model_1.B_next [2], ABINPUT001[2]);
  buf(\oc8051_golden_model_1.B_next [3], ABINPUT001[3]);
  buf(\oc8051_golden_model_1.B_next [4], ABINPUT001[4]);
  buf(\oc8051_golden_model_1.B_next [5], ABINPUT001[5]);
  buf(\oc8051_golden_model_1.B_next [6], ABINPUT001[6]);
  buf(\oc8051_golden_model_1.B_next [7], ABINPUT001[7]);
  buf(\oc8051_golden_model_1.ABINPUT000 [0], ABINPUT001[0]);
  buf(\oc8051_golden_model_1.ABINPUT000 [1], ABINPUT001[1]);
  buf(\oc8051_golden_model_1.ABINPUT000 [2], ABINPUT001[2]);
  buf(\oc8051_golden_model_1.ABINPUT000 [3], ABINPUT001[3]);
  buf(\oc8051_golden_model_1.ABINPUT000 [4], ABINPUT001[4]);
  buf(\oc8051_golden_model_1.ABINPUT000 [5], ABINPUT001[5]);
  buf(\oc8051_golden_model_1.ABINPUT000 [6], ABINPUT001[6]);
  buf(\oc8051_golden_model_1.ABINPUT000 [7], ABINPUT001[7]);
  buf(\oc8051_golden_model_1.n2453 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2453 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2453 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2453 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2453 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2453 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2453 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2453 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2454 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2454 [1], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.n2454 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2454 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2454 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2454 [5], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.n2454 [6], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.n2876 [0], \oc8051_golden_model_1.PSW_d6 [0]);
  buf(\oc8051_golden_model_1.n2876 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2876 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2876 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2876 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2876 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2876 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2876 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.PSW_26 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.PSW_26 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.PSW_29 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.PSW_29 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.PSW_29 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.PSW_29 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.PSW_2c [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.PSW_2a [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.PSW_2c [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.PSW_2a [6]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.PSW_29 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.PSW_29 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.PSW_2c [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.PSW_2c [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.PSW_2c [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.PSW_2c [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.PSW_36 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.PSW_36 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.PSW_36 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.PSW_36 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.PSW_3b [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.PSW_3b [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.PSW_3b [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.PSW_3b [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.PSW_3b [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.PSW_3b [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.PSW_3b [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.PSW_3b [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.PSW_3b [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.PSW_3b [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.PSW_3b [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.PSW_3b [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.PSW_3b [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.PSW_3b [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1805 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1822 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.PSW_47 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.PSW_57 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.PSW_67 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.PSW_68 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.PSW_68 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.PSW_68 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.PSW_68 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.PSW_68 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.PSW_68 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.PSW_68 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.PSW_74 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.PSW_74 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2470 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2470 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2470 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2484 [1]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2484 [5]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2484 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.PSW_97 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.PSW_97 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.PSW_97 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.PSW_97 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.PSW_98 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.PSW_98 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.PSW_98 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.PSW_98 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.PSW_98 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.PSW_98 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.PSW_98 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.PSW_98 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.PSW_98 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.PSW_98 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.PSW_98 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.PSW_98 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.PSW_98 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.PSW_98 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.PSW_98 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.PSW_98 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.PSW_98 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.PSW_98 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.PSW_98 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.PSW_98 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.PSW_98 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.PSW_98 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.PSW_98 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.PSW_98 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.PSW_98 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.PSW_98 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.PSW_98 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.PSW_98 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.PSW_d6 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2896 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fa [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_fa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fb [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_fb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fc [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_fc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fd [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_fd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fe [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_fe [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fe [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fe [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fe [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fe [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fe [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fe [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ff [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.PSW_ff [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ff [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ff [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ff [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ff [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ff [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ff [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0573 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n0573 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n0573 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n0573 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n0573 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n0573 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n0573 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n0573 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n0606 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n0606 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n0606 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n0606 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n0606 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n0606 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n0606 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n0606 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n0713 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0713 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0713 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0713 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0713 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0713 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0713 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0713 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0713 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0745 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0745 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0745 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0745 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0745 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0745 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0745 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0745 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0745 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0745 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0745 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0745 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0745 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0745 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0745 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0745 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n1004 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1004 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1004 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1004 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1004 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1004 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1004 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1004 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1004 [8], \oc8051_golden_model_1.P2 [0]);
  buf(\oc8051_golden_model_1.n1004 [9], \oc8051_golden_model_1.P2 [1]);
  buf(\oc8051_golden_model_1.n1004 [10], \oc8051_golden_model_1.P2 [2]);
  buf(\oc8051_golden_model_1.n1004 [11], \oc8051_golden_model_1.P2 [3]);
  buf(\oc8051_golden_model_1.n1004 [12], \oc8051_golden_model_1.P2 [4]);
  buf(\oc8051_golden_model_1.n1004 [13], \oc8051_golden_model_1.P2 [5]);
  buf(\oc8051_golden_model_1.n1004 [14], \oc8051_golden_model_1.P2 [6]);
  buf(\oc8051_golden_model_1.n1004 [15], \oc8051_golden_model_1.P2 [7]);
  buf(\oc8051_golden_model_1.n1008 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1008 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1008 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1008 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1008 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1008 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1008 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1009 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1010 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1011 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1012 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1013 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1014 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1015 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1016 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1023 , \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n1024 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n1024 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1024 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1024 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1024 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1024 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1024 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1024 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1031 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1031 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1031 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1031 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1031 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1031 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1031 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1031 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1032 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1033 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1034 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1035 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1036 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1037 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1038 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1039 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1047 [0], \oc8051_golden_model_1.PSW_03 [0]);
  buf(\oc8051_golden_model_1.n1047 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1047 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1047 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1047 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1047 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1047 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1047 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1064 [0], \oc8051_golden_model_1.PSW_04 [0]);
  buf(\oc8051_golden_model_1.n1064 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1064 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1064 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1064 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1064 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1064 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1064 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2469 , \oc8051_golden_model_1.n2470 [0]);
  buf(\oc8051_golden_model_1.n2470 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2470 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2470 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2470 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2474 , \oc8051_golden_model_1.n2484 [6]);
  buf(\oc8051_golden_model_1.n2476 , \oc8051_golden_model_1.n2484 [5]);
  buf(\oc8051_golden_model_1.n2482 , \oc8051_golden_model_1.n2484 [1]);
  buf(\oc8051_golden_model_1.n2483 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2483 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2483 [2], \oc8051_golden_model_1.n2484 [1]);
  buf(\oc8051_golden_model_1.n2483 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2483 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2483 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2483 [6], \oc8051_golden_model_1.n2484 [5]);
  buf(\oc8051_golden_model_1.n2483 [7], \oc8051_golden_model_1.n2484 [6]);
  buf(\oc8051_golden_model_1.n2484 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2484 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2484 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2484 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1157 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1157 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1157 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1157 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1159 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1159 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1161 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1161 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1162 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1162 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1162 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1163 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1163 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1163 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1164 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1164 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1164 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1165 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1165 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1165 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1166 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1166 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1166 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1167 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1167 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2499 , \oc8051_golden_model_1.n2500 [0]);
  buf(\oc8051_golden_model_1.n2500 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2500 [2], \oc8051_golden_model_1.n2484 [1]);
  buf(\oc8051_golden_model_1.n2500 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2500 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2500 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2500 [6], \oc8051_golden_model_1.n2484 [5]);
  buf(\oc8051_golden_model_1.n2500 [7], \oc8051_golden_model_1.n2484 [6]);
  buf(\oc8051_golden_model_1.n2504 , \oc8051_golden_model_1.PSW_97 [7]);
  buf(\oc8051_golden_model_1.n2506 , \oc8051_golden_model_1.PSW_97 [6]);
  buf(\oc8051_golden_model_1.n2512 , \oc8051_golden_model_1.PSW_97 [2]);
  buf(\oc8051_golden_model_1.n2513 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2513 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2513 [2], \oc8051_golden_model_1.PSW_97 [2]);
  buf(\oc8051_golden_model_1.n2513 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2513 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2513 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2513 [6], \oc8051_golden_model_1.PSW_97 [6]);
  buf(\oc8051_golden_model_1.n2513 [7], \oc8051_golden_model_1.PSW_97 [7]);
  buf(\oc8051_golden_model_1.n2514 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2514 [1], \oc8051_golden_model_1.PSW_97 [2]);
  buf(\oc8051_golden_model_1.n2514 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2514 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2514 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2514 [5], \oc8051_golden_model_1.PSW_97 [6]);
  buf(\oc8051_golden_model_1.n2514 [6], \oc8051_golden_model_1.PSW_97 [7]);
  buf(\oc8051_golden_model_1.n1259 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1260 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1261 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1261 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1261 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1261 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1261 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1261 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1261 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1261 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1262 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1262 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1262 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1262 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1262 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1262 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1262 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1262 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1265 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1266 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1266 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1267 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1267 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1267 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1267 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1267 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1267 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1267 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1268 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1268 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1268 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1268 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1268 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1268 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1268 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1269 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1270 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1271 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1272 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1273 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1274 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1276 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1284 [0], \oc8051_golden_model_1.PSW_13 [0]);
  buf(\oc8051_golden_model_1.n1284 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1284 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1284 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1284 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1284 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1284 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1284 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2529 , \oc8051_golden_model_1.PSW_97 [0]);
  buf(\oc8051_golden_model_1.n2530 [0], \oc8051_golden_model_1.PSW_97 [0]);
  buf(\oc8051_golden_model_1.n2530 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2530 [2], \oc8051_golden_model_1.PSW_97 [2]);
  buf(\oc8051_golden_model_1.n2530 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2530 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2530 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2530 [6], \oc8051_golden_model_1.PSW_97 [6]);
  buf(\oc8051_golden_model_1.n2530 [7], \oc8051_golden_model_1.PSW_97 [7]);
  buf(\oc8051_golden_model_1.n2534 , \oc8051_golden_model_1.PSW_98 [7]);
  buf(\oc8051_golden_model_1.n2536 , \oc8051_golden_model_1.PSW_98 [6]);
  buf(\oc8051_golden_model_1.n1301 [0], \oc8051_golden_model_1.PSW_14 [0]);
  buf(\oc8051_golden_model_1.n1301 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1301 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1301 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1301 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1301 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1301 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1301 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2542 , \oc8051_golden_model_1.PSW_98 [2]);
  buf(\oc8051_golden_model_1.n2543 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2543 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2543 [2], \oc8051_golden_model_1.PSW_98 [2]);
  buf(\oc8051_golden_model_1.n2543 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2543 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2543 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2543 [6], \oc8051_golden_model_1.PSW_98 [6]);
  buf(\oc8051_golden_model_1.n2543 [7], \oc8051_golden_model_1.PSW_98 [7]);
  buf(\oc8051_golden_model_1.n2544 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2544 [1], \oc8051_golden_model_1.PSW_98 [2]);
  buf(\oc8051_golden_model_1.n2544 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2544 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2544 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2544 [5], \oc8051_golden_model_1.PSW_98 [6]);
  buf(\oc8051_golden_model_1.n2544 [6], \oc8051_golden_model_1.PSW_98 [7]);
  buf(\oc8051_golden_model_1.n2559 , \oc8051_golden_model_1.PSW_98 [0]);
  buf(\oc8051_golden_model_1.n2560 [0], \oc8051_golden_model_1.PSW_98 [0]);
  buf(\oc8051_golden_model_1.n2560 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2560 [2], \oc8051_golden_model_1.PSW_98 [2]);
  buf(\oc8051_golden_model_1.n2560 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2560 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2560 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2560 [6], \oc8051_golden_model_1.PSW_98 [6]);
  buf(\oc8051_golden_model_1.n2560 [7], \oc8051_golden_model_1.PSW_98 [7]);
  buf(\oc8051_golden_model_1.n2563 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2563 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2563 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2563 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2563 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2563 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2563 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2563 [7], \oc8051_golden_model_1.PSW_a0 [7]);
  buf(\oc8051_golden_model_1.n2564 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2564 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2564 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2564 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2564 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2564 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2564 [6], \oc8051_golden_model_1.PSW_a0 [7]);
  buf(\oc8051_golden_model_1.n2565 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2565 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2565 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2565 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2565 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2565 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2565 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2565 [7], \oc8051_golden_model_1.PSW_a0 [7]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1343 [8], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1343 [9], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1343 [10], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1343 [11], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1343 [12], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1343 [13], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1343 [14], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1343 [15], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1345 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1345 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1345 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1345 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1345 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1345 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1345 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1345 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1346 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1347 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1348 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1350 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1351 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1352 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1353 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2566 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2566 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2566 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2566 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2566 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2566 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2566 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2566 [7], \oc8051_golden_model_1.PSW_a2 [7]);
  buf(\oc8051_golden_model_1.n2567 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2567 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2567 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2567 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2567 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2567 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2567 [6], \oc8051_golden_model_1.PSW_a2 [7]);
  buf(\oc8051_golden_model_1.n2568 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2568 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2568 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2568 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2568 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2568 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2568 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2568 [7], \oc8051_golden_model_1.PSW_a2 [7]);
  buf(\oc8051_golden_model_1.n1361 [0], \oc8051_golden_model_1.PSW_23 [0]);
  buf(\oc8051_golden_model_1.n1361 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1361 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1361 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1361 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1361 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1361 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1361 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2572 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2572 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2572 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2572 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2572 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2572 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2572 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2572 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2572 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2572 [15], 1'b0);
  buf(\oc8051_golden_model_1.n1363 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1363 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1363 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1363 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1363 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1363 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1363 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1363 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1363 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1369 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1369 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1369 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1369 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1370 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1370 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1370 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1370 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1376 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1376 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1376 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1376 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1376 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1376 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1376 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1376 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1376 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2578 , \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2579 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2579 [2], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2579 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2579 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2579 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2579 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2579 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2580 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2580 [1], \oc8051_golden_model_1.n2596 [2]);
  buf(\oc8051_golden_model_1.n2580 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2580 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2580 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2580 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2580 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1385 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1385 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1385 [2], \oc8051_golden_model_1.PSW_24 [2]);
  buf(\oc8051_golden_model_1.n1385 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1385 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1385 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1385 [6], \oc8051_golden_model_1.PSW_24 [6]);
  buf(\oc8051_golden_model_1.n1385 [7], \oc8051_golden_model_1.PSW_24 [7]);
  buf(\oc8051_golden_model_1.n1386 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1386 [1], \oc8051_golden_model_1.PSW_24 [2]);
  buf(\oc8051_golden_model_1.n1386 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1386 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1386 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1386 [5], \oc8051_golden_model_1.PSW_24 [6]);
  buf(\oc8051_golden_model_1.n1386 [6], \oc8051_golden_model_1.PSW_24 [7]);
  buf(\oc8051_golden_model_1.n2595 , \oc8051_golden_model_1.n2596 [0]);
  buf(\oc8051_golden_model_1.n2596 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2596 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2596 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2596 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2596 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2596 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1402 [0], \oc8051_golden_model_1.PSW_24 [0]);
  buf(\oc8051_golden_model_1.n1402 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1402 [2], \oc8051_golden_model_1.PSW_24 [2]);
  buf(\oc8051_golden_model_1.n1402 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1402 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1402 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1402 [6], \oc8051_golden_model_1.PSW_24 [6]);
  buf(\oc8051_golden_model_1.n1402 [7], \oc8051_golden_model_1.PSW_24 [7]);
  buf(\oc8051_golden_model_1.n2599 , \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2600 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2600 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2600 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2600 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2600 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2600 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2600 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2600 [7], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2601 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2601 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2601 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2601 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2601 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2601 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2601 [6], \oc8051_golden_model_1.n2602 [7]);
  buf(\oc8051_golden_model_1.n2602 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2602 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2602 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2602 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2602 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2602 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2602 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1440 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1440 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1440 [2], \oc8051_golden_model_1.PSW_25 [2]);
  buf(\oc8051_golden_model_1.n1440 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1440 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1440 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1440 [6], \oc8051_golden_model_1.PSW_25 [6]);
  buf(\oc8051_golden_model_1.n1440 [7], \oc8051_golden_model_1.PSW_25 [7]);
  buf(\oc8051_golden_model_1.n1441 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1441 [1], \oc8051_golden_model_1.PSW_25 [2]);
  buf(\oc8051_golden_model_1.n1441 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1441 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1441 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1441 [5], \oc8051_golden_model_1.PSW_25 [6]);
  buf(\oc8051_golden_model_1.n1441 [6], \oc8051_golden_model_1.PSW_25 [7]);
  buf(\oc8051_golden_model_1.n1457 [0], \oc8051_golden_model_1.PSW_25 [0]);
  buf(\oc8051_golden_model_1.n1457 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1457 [2], \oc8051_golden_model_1.PSW_25 [2]);
  buf(\oc8051_golden_model_1.n1457 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1457 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1457 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1457 [6], \oc8051_golden_model_1.PSW_25 [6]);
  buf(\oc8051_golden_model_1.n1457 [7], \oc8051_golden_model_1.PSW_25 [7]);
  buf(\oc8051_golden_model_1.n1459 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n1459 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n1459 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n1459 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n1459 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1459 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1459 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1459 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1459 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1463 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n1463 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n1463 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n1463 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n1464 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n1464 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n1464 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n1464 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n1464 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1466 [4], \oc8051_golden_model_1.PSW_26 [6]);
  buf(\oc8051_golden_model_1.n1467 , \oc8051_golden_model_1.PSW_26 [6]);
  buf(\oc8051_golden_model_1.n1468 [0], \oc8051_golden_model_1.n2759 );
  buf(\oc8051_golden_model_1.n1468 [1], \oc8051_golden_model_1.n2758 );
  buf(\oc8051_golden_model_1.n1468 [2], \oc8051_golden_model_1.n2757 );
  buf(\oc8051_golden_model_1.n1468 [3], \oc8051_golden_model_1.n2756 );
  buf(\oc8051_golden_model_1.n1468 [4], \oc8051_golden_model_1.n2755 );
  buf(\oc8051_golden_model_1.n1468 [5], \oc8051_golden_model_1.n2754 );
  buf(\oc8051_golden_model_1.n1468 [6], \oc8051_golden_model_1.n2753 );
  buf(\oc8051_golden_model_1.n1468 [7], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1468 [8], \oc8051_golden_model_1.n2752 );
  buf(\oc8051_golden_model_1.n1476 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1476 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1476 [2], \oc8051_golden_model_1.PSW_26 [2]);
  buf(\oc8051_golden_model_1.n1476 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1476 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1476 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1476 [6], \oc8051_golden_model_1.PSW_26 [6]);
  buf(\oc8051_golden_model_1.n1476 [7], \oc8051_golden_model_1.PSW_26 [7]);
  buf(\oc8051_golden_model_1.n1477 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1477 [1], \oc8051_golden_model_1.PSW_26 [2]);
  buf(\oc8051_golden_model_1.n1477 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1477 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1477 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1477 [5], \oc8051_golden_model_1.PSW_26 [6]);
  buf(\oc8051_golden_model_1.n1477 [6], \oc8051_golden_model_1.PSW_26 [7]);
  buf(\oc8051_golden_model_1.n2634 , \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2635 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2635 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2635 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2635 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2635 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2635 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2635 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2635 [7], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2636 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2636 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2636 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2636 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2636 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2636 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2636 [6], \oc8051_golden_model_1.n2637 [7]);
  buf(\oc8051_golden_model_1.n2637 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2637 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2637 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2637 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2637 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2637 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2637 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2642 , \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2643 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2643 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2643 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2643 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2643 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2643 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2643 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2643 [7], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n1492 , \oc8051_golden_model_1.PSW_26 [0]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.PSW_26 [0]);
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1493 [2], \oc8051_golden_model_1.PSW_26 [2]);
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1493 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1493 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1493 [6], \oc8051_golden_model_1.PSW_26 [6]);
  buf(\oc8051_golden_model_1.n1493 [7], \oc8051_golden_model_1.PSW_26 [7]);
  buf(\oc8051_golden_model_1.n2644 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2644 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2644 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2644 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2644 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2644 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2644 [6], \oc8051_golden_model_1.n2645 [7]);
  buf(\oc8051_golden_model_1.n2645 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2645 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2645 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2645 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2645 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2645 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2645 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2650 , \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n2651 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2651 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2651 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2651 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2651 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2651 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2651 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2651 [7], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n1505 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1505 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1505 [2], \oc8051_golden_model_1.PSW_27 [2]);
  buf(\oc8051_golden_model_1.n1505 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1505 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1505 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1505 [6], \oc8051_golden_model_1.PSW_26 [6]);
  buf(\oc8051_golden_model_1.n1505 [7], \oc8051_golden_model_1.PSW_27 [7]);
  buf(\oc8051_golden_model_1.n1506 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1506 [1], \oc8051_golden_model_1.PSW_27 [2]);
  buf(\oc8051_golden_model_1.n1506 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1506 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1506 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1506 [5], \oc8051_golden_model_1.PSW_26 [6]);
  buf(\oc8051_golden_model_1.n1506 [6], \oc8051_golden_model_1.PSW_27 [7]);
  buf(\oc8051_golden_model_1.n1507 [0], \oc8051_golden_model_1.PSW_26 [0]);
  buf(\oc8051_golden_model_1.n1507 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1507 [2], \oc8051_golden_model_1.PSW_27 [2]);
  buf(\oc8051_golden_model_1.n1507 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1507 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1507 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1507 [6], \oc8051_golden_model_1.PSW_26 [6]);
  buf(\oc8051_golden_model_1.n1507 [7], \oc8051_golden_model_1.PSW_27 [7]);
  buf(\oc8051_golden_model_1.n2652 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2652 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2652 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2652 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2652 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2652 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2652 [6], \oc8051_golden_model_1.n2653 [7]);
  buf(\oc8051_golden_model_1.n1509 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1509 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1509 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1509 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1509 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1509 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1509 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1509 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1509 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2653 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2653 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2653 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2653 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2653 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2653 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2653 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1511 [8], \oc8051_golden_model_1.PSW_29 [7]);
  buf(\oc8051_golden_model_1.n1512 , \oc8051_golden_model_1.PSW_29 [7]);
  buf(\oc8051_golden_model_1.n1513 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1513 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1513 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1513 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1513 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1515 [4], \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.n1516 , \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.n1517 [0], \oc8051_golden_model_1.n2775 );
  buf(\oc8051_golden_model_1.n1517 [1], \oc8051_golden_model_1.n2774 );
  buf(\oc8051_golden_model_1.n1517 [2], \oc8051_golden_model_1.n2773 );
  buf(\oc8051_golden_model_1.n1517 [3], \oc8051_golden_model_1.n2772 );
  buf(\oc8051_golden_model_1.n1517 [4], \oc8051_golden_model_1.n2771 );
  buf(\oc8051_golden_model_1.n1517 [5], \oc8051_golden_model_1.n2770 );
  buf(\oc8051_golden_model_1.n1517 [6], \oc8051_golden_model_1.n2769 );
  buf(\oc8051_golden_model_1.n1517 [7], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n1517 [8], \oc8051_golden_model_1.n2768 );
  buf(\oc8051_golden_model_1.n2658 , \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2659 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2659 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2659 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2659 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2659 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2659 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2659 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2659 [7], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n2660 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2660 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2660 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2660 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2660 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2660 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2660 [6], \oc8051_golden_model_1.n2661 [7]);
  buf(\oc8051_golden_model_1.n1524 , \oc8051_golden_model_1.PSW_29 [2]);
  buf(\oc8051_golden_model_1.n1525 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1525 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1525 [2], \oc8051_golden_model_1.PSW_29 [2]);
  buf(\oc8051_golden_model_1.n1525 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1525 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1525 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1525 [6], \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.n1525 [7], \oc8051_golden_model_1.PSW_29 [7]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.PSW_29 [2]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.PSW_29 [7]);
  buf(\oc8051_golden_model_1.n2661 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2661 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2661 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2661 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2661 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2661 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2661 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2666 , \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2667 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2667 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2667 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2667 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2667 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2667 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2667 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2667 [7], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2668 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2668 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2668 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2668 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2668 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2668 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2668 [6], \oc8051_golden_model_1.n2669 [7]);
  buf(\oc8051_golden_model_1.n2669 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2669 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2669 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1541 , \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.n1542 [0], \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.n1542 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1542 [2], \oc8051_golden_model_1.PSW_29 [2]);
  buf(\oc8051_golden_model_1.n1542 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1542 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1542 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1542 [6], \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.n1542 [7], \oc8051_golden_model_1.PSW_29 [7]);
  buf(\oc8051_golden_model_1.n1544 [4], \oc8051_golden_model_1.PSW_2a [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.PSW_2a [6]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.PSW_29 [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.PSW_2a [6]);
  buf(\oc8051_golden_model_1.n1546 [7], \oc8051_golden_model_1.PSW_29 [7]);
  buf(\oc8051_golden_model_1.n1547 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1547 [1], \oc8051_golden_model_1.PSW_29 [2]);
  buf(\oc8051_golden_model_1.n1547 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1547 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1547 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1547 [5], \oc8051_golden_model_1.PSW_2a [6]);
  buf(\oc8051_golden_model_1.n1547 [6], \oc8051_golden_model_1.PSW_29 [7]);
  buf(\oc8051_golden_model_1.n1548 [0], \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.n1548 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1548 [2], \oc8051_golden_model_1.PSW_29 [2]);
  buf(\oc8051_golden_model_1.n1548 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1548 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1548 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1548 [6], \oc8051_golden_model_1.PSW_2a [6]);
  buf(\oc8051_golden_model_1.n1548 [7], \oc8051_golden_model_1.PSW_29 [7]);
  buf(\oc8051_golden_model_1.n1550 [8], \oc8051_golden_model_1.PSW_2c [7]);
  buf(\oc8051_golden_model_1.n1551 , \oc8051_golden_model_1.PSW_2c [7]);
  buf(\oc8051_golden_model_1.n2894 , \oc8051_golden_model_1.n2895 [0]);
  buf(\oc8051_golden_model_1.n2895 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2895 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2895 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2895 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2895 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2895 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2895 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2896 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2896 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2896 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2896 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2896 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2896 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2896 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.PSW_2c [2]);
  buf(\oc8051_golden_model_1.n1559 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1559 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1559 [2], \oc8051_golden_model_1.PSW_2c [2]);
  buf(\oc8051_golden_model_1.n1559 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1559 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1559 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1559 [6], \oc8051_golden_model_1.PSW_2a [6]);
  buf(\oc8051_golden_model_1.n1559 [7], \oc8051_golden_model_1.PSW_2c [7]);
  buf(\oc8051_golden_model_1.n1560 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1560 [1], \oc8051_golden_model_1.PSW_2c [2]);
  buf(\oc8051_golden_model_1.n1560 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1560 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1560 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1560 [5], \oc8051_golden_model_1.PSW_2a [6]);
  buf(\oc8051_golden_model_1.n1560 [6], \oc8051_golden_model_1.PSW_2c [7]);
  buf(\oc8051_golden_model_1.n1561 [0], \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.n1561 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1561 [2], \oc8051_golden_model_1.PSW_2c [2]);
  buf(\oc8051_golden_model_1.n1561 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1561 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1561 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1561 [6], \oc8051_golden_model_1.PSW_2a [6]);
  buf(\oc8051_golden_model_1.n1561 [7], \oc8051_golden_model_1.PSW_2c [7]);
  buf(\oc8051_golden_model_1.n1562 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1562 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1562 [2], \oc8051_golden_model_1.PSW_2c [2]);
  buf(\oc8051_golden_model_1.n1562 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1562 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1562 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1562 [6], \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.n1562 [7], \oc8051_golden_model_1.PSW_2c [7]);
  buf(\oc8051_golden_model_1.n1563 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1563 [1], \oc8051_golden_model_1.PSW_2c [2]);
  buf(\oc8051_golden_model_1.n1563 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1563 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1563 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1563 [5], \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.n1563 [6], \oc8051_golden_model_1.PSW_2c [7]);
  buf(\oc8051_golden_model_1.n1564 [0], \oc8051_golden_model_1.PSW_29 [0]);
  buf(\oc8051_golden_model_1.n1564 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1564 [2], \oc8051_golden_model_1.PSW_2c [2]);
  buf(\oc8051_golden_model_1.n1564 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1564 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1564 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1564 [6], \oc8051_golden_model_1.PSW_29 [6]);
  buf(\oc8051_golden_model_1.n1564 [7], \oc8051_golden_model_1.PSW_2c [7]);
  buf(\oc8051_golden_model_1.n1567 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1567 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1567 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1567 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1567 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1567 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1567 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1567 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1567 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1568 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1568 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1568 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1568 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1568 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1568 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1568 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1568 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1569 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1569 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1569 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1569 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1569 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1569 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1569 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1569 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1570 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1570 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1570 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1570 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1570 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1570 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1570 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1570 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1571 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1571 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1571 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1571 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1571 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1571 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1572 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1573 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1574 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1575 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1576 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1577 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1578 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1579 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1587 [0], \oc8051_golden_model_1.PSW_33 [0]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1587 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1587 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1588 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1588 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1588 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1591 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1591 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1595 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1595 [4], 1'b0);
  buf(\oc8051_golden_model_1.n2694 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2694 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2694 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2694 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2694 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2694 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2694 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2694 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2695 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2695 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2695 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2695 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2695 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2695 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2695 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2696 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2696 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2696 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2696 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2696 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2696 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2696 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2696 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2697 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2697 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2697 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2697 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2698 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2698 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2698 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2698 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2698 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2698 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2698 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1606 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1606 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1606 [2], \oc8051_golden_model_1.PSW_34 [2]);
  buf(\oc8051_golden_model_1.n1606 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1606 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1606 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1606 [6], \oc8051_golden_model_1.PSW_34 [6]);
  buf(\oc8051_golden_model_1.n1606 [7], \oc8051_golden_model_1.PSW_34 [7]);
  buf(\oc8051_golden_model_1.n1607 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1607 [1], \oc8051_golden_model_1.PSW_34 [2]);
  buf(\oc8051_golden_model_1.n1607 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1607 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1607 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1607 [5], \oc8051_golden_model_1.PSW_34 [6]);
  buf(\oc8051_golden_model_1.n1607 [6], \oc8051_golden_model_1.PSW_34 [7]);
  buf(\oc8051_golden_model_1.n2699 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2700 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2701 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2702 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2703 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2704 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2705 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2706 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2912 , \oc8051_golden_model_1.n2913 [0]);
  buf(\oc8051_golden_model_1.n2913 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2913 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2913 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2913 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2913 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2913 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2913 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1623 [0], \oc8051_golden_model_1.PSW_34 [0]);
  buf(\oc8051_golden_model_1.n1623 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1623 [2], \oc8051_golden_model_1.PSW_34 [2]);
  buf(\oc8051_golden_model_1.n1623 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1623 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1623 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1623 [6], \oc8051_golden_model_1.PSW_34 [6]);
  buf(\oc8051_golden_model_1.n1623 [7], \oc8051_golden_model_1.PSW_34 [7]);
  buf(\oc8051_golden_model_1.n2713 , \oc8051_golden_model_1.n2714 [0]);
  buf(\oc8051_golden_model_1.n2714 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2714 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2714 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2714 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2714 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2714 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2714 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1639 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1639 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1639 [2], \oc8051_golden_model_1.PSW_35 [2]);
  buf(\oc8051_golden_model_1.n1639 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1639 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1639 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1639 [6], \oc8051_golden_model_1.PSW_35 [6]);
  buf(\oc8051_golden_model_1.n1639 [7], \oc8051_golden_model_1.PSW_35 [7]);
  buf(\oc8051_golden_model_1.n1640 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1640 [1], \oc8051_golden_model_1.PSW_35 [2]);
  buf(\oc8051_golden_model_1.n1640 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1640 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1640 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1640 [5], \oc8051_golden_model_1.PSW_35 [6]);
  buf(\oc8051_golden_model_1.n1640 [6], \oc8051_golden_model_1.PSW_35 [7]);
  buf(\oc8051_golden_model_1.n1656 [0], \oc8051_golden_model_1.PSW_35 [0]);
  buf(\oc8051_golden_model_1.n1656 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1656 [2], \oc8051_golden_model_1.PSW_35 [2]);
  buf(\oc8051_golden_model_1.n1656 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1656 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1656 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1656 [6], \oc8051_golden_model_1.PSW_35 [6]);
  buf(\oc8051_golden_model_1.n1656 [7], \oc8051_golden_model_1.PSW_35 [7]);
  buf(\oc8051_golden_model_1.n1660 [8], \oc8051_golden_model_1.PSW_36 [7]);
  buf(\oc8051_golden_model_1.n1661 , \oc8051_golden_model_1.PSW_36 [7]);
  buf(\oc8051_golden_model_1.n1663 [4], \oc8051_golden_model_1.PSW_36 [6]);
  buf(\oc8051_golden_model_1.n1664 , \oc8051_golden_model_1.PSW_36 [6]);
  buf(\oc8051_golden_model_1.n1671 , \oc8051_golden_model_1.PSW_36 [2]);
  buf(\oc8051_golden_model_1.n1672 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1672 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1672 [2], \oc8051_golden_model_1.PSW_36 [2]);
  buf(\oc8051_golden_model_1.n1672 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1672 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1672 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1672 [6], \oc8051_golden_model_1.PSW_36 [6]);
  buf(\oc8051_golden_model_1.n1672 [7], \oc8051_golden_model_1.PSW_36 [7]);
  buf(\oc8051_golden_model_1.n1673 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1673 [1], \oc8051_golden_model_1.PSW_36 [2]);
  buf(\oc8051_golden_model_1.n1673 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1673 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1673 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1673 [5], \oc8051_golden_model_1.PSW_36 [6]);
  buf(\oc8051_golden_model_1.n1673 [6], \oc8051_golden_model_1.PSW_36 [7]);
  buf(\oc8051_golden_model_1.n1688 , \oc8051_golden_model_1.PSW_36 [0]);
  buf(\oc8051_golden_model_1.n1689 [0], \oc8051_golden_model_1.PSW_36 [0]);
  buf(\oc8051_golden_model_1.n1689 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1689 [2], \oc8051_golden_model_1.PSW_36 [2]);
  buf(\oc8051_golden_model_1.n1689 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1689 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1689 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1689 [6], \oc8051_golden_model_1.PSW_36 [6]);
  buf(\oc8051_golden_model_1.n1689 [7], \oc8051_golden_model_1.PSW_36 [7]);
  buf(\oc8051_golden_model_1.n1693 [8], \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.n1694 , \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.n1696 [4], \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.n1697 , \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.PSW_3b [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [2], \oc8051_golden_model_1.PSW_3b [2]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1705 [6], \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.n1705 [7], \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.n1706 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1706 [1], \oc8051_golden_model_1.PSW_3b [2]);
  buf(\oc8051_golden_model_1.n1706 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1706 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1706 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1706 [5], \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.n1706 [6], \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.n1721 , \oc8051_golden_model_1.PSW_3b [0]);
  buf(\oc8051_golden_model_1.n1722 [0], \oc8051_golden_model_1.PSW_3b [0]);
  buf(\oc8051_golden_model_1.n1722 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1722 [2], \oc8051_golden_model_1.PSW_3b [2]);
  buf(\oc8051_golden_model_1.n1722 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1722 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1722 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1722 [6], \oc8051_golden_model_1.PSW_3b [6]);
  buf(\oc8051_golden_model_1.n1722 [7], \oc8051_golden_model_1.PSW_3b [7]);
  buf(\oc8051_golden_model_1.n1749 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n1749 [1], \oc8051_golden_model_1.PSW_42 [1]);
  buf(\oc8051_golden_model_1.n1749 [2], \oc8051_golden_model_1.PSW_42 [2]);
  buf(\oc8051_golden_model_1.n1749 [3], \oc8051_golden_model_1.PSW_42 [3]);
  buf(\oc8051_golden_model_1.n1749 [4], \oc8051_golden_model_1.PSW_42 [4]);
  buf(\oc8051_golden_model_1.n1749 [5], \oc8051_golden_model_1.PSW_42 [5]);
  buf(\oc8051_golden_model_1.n1749 [6], \oc8051_golden_model_1.PSW_42 [6]);
  buf(\oc8051_golden_model_1.n1749 [7], \oc8051_golden_model_1.PSW_42 [7]);
  buf(\oc8051_golden_model_1.n1804 , \oc8051_golden_model_1.n1805 [0]);
  buf(\oc8051_golden_model_1.n1805 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1805 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1805 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1805 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1805 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1805 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1805 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1821 , \oc8051_golden_model_1.n1822 [0]);
  buf(\oc8051_golden_model_1.n1822 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1822 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1822 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1822 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1822 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1822 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1822 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1838 , \oc8051_golden_model_1.PSW_47 [0]);
  buf(\oc8051_golden_model_1.n1839 [0], \oc8051_golden_model_1.PSW_47 [0]);
  buf(\oc8051_golden_model_1.n1839 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1839 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1839 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1839 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1839 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1839 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1839 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1855 , \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.n1856 [0], \oc8051_golden_model_1.PSW_48 [0]);
  buf(\oc8051_golden_model_1.n1856 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1856 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1856 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1856 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1856 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1856 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1856 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1881 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n1881 [1], \oc8051_golden_model_1.PSW_52 [1]);
  buf(\oc8051_golden_model_1.n1881 [2], \oc8051_golden_model_1.PSW_52 [2]);
  buf(\oc8051_golden_model_1.n1881 [3], \oc8051_golden_model_1.PSW_52 [3]);
  buf(\oc8051_golden_model_1.n1881 [4], \oc8051_golden_model_1.PSW_52 [4]);
  buf(\oc8051_golden_model_1.n1881 [5], \oc8051_golden_model_1.PSW_52 [5]);
  buf(\oc8051_golden_model_1.n1881 [6], \oc8051_golden_model_1.PSW_52 [6]);
  buf(\oc8051_golden_model_1.n1881 [7], \oc8051_golden_model_1.PSW_52 [7]);
  buf(\oc8051_golden_model_1.n2766 , \oc8051_golden_model_1.n2767 [0]);
  buf(\oc8051_golden_model_1.n2767 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2767 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2767 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2767 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2767 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2767 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2767 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2782 , \oc8051_golden_model_1.n2783 [0]);
  buf(\oc8051_golden_model_1.n2783 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2783 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2783 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2783 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2783 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2783 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2783 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1937 [0], \oc8051_golden_model_1.PSW_54 [0]);
  buf(\oc8051_golden_model_1.n1937 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1937 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1937 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1937 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1937 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1937 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1937 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1954 [0], \oc8051_golden_model_1.PSW_55 [0]);
  buf(\oc8051_golden_model_1.n1954 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1954 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1954 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1954 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1954 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1954 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1954 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1970 , \oc8051_golden_model_1.PSW_57 [0]);
  buf(\oc8051_golden_model_1.n1971 [0], \oc8051_golden_model_1.PSW_57 [0]);
  buf(\oc8051_golden_model_1.n1971 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1971 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1971 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1971 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1971 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1971 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1971 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2815 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2815 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2815 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2815 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2815 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2815 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2815 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2815 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2816 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2816 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2816 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2816 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2816 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2816 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2816 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2817 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2817 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2817 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2817 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2817 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2817 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2817 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2817 [7], 1'b1);
  buf(\oc8051_golden_model_1.n1987 , \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.n1988 [0], \oc8051_golden_model_1.PSW_58 [0]);
  buf(\oc8051_golden_model_1.n1988 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1988 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1988 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1988 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1988 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1988 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1988 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2836 , \oc8051_golden_model_1.PSW_d4 [7]);
  buf(\oc8051_golden_model_1.n2837 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2837 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2837 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2837 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2837 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2837 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2837 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2837 [7], \oc8051_golden_model_1.PSW_d4 [7]);
  buf(\oc8051_golden_model_1.n2838 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2838 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2838 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2838 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2838 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2838 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2838 [6], \oc8051_golden_model_1.PSW_d4 [7]);
  buf(\oc8051_golden_model_1.n2086 [0], \oc8051_golden_model_1.PSW_64 [0]);
  buf(\oc8051_golden_model_1.n2086 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2086 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2086 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2086 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2086 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2086 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2086 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2103 [0], \oc8051_golden_model_1.PSW_65 [0]);
  buf(\oc8051_golden_model_1.n2103 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2103 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2103 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2103 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2103 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2103 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2103 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2119 , \oc8051_golden_model_1.PSW_67 [0]);
  buf(\oc8051_golden_model_1.n2120 [0], \oc8051_golden_model_1.PSW_67 [0]);
  buf(\oc8051_golden_model_1.n2120 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2120 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2120 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2120 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2120 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2120 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2120 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2136 , \oc8051_golden_model_1.PSW_68 [0]);
  buf(\oc8051_golden_model_1.n2137 [0], \oc8051_golden_model_1.PSW_68 [0]);
  buf(\oc8051_golden_model_1.n2137 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2137 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2137 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2137 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2137 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2137 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2137 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2142 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2142 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2142 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2142 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2142 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2142 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2142 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2143 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2143 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2143 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2143 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2143 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2143 [7], \oc8051_golden_model_1.PSW_72 [7]);
  buf(\oc8051_golden_model_1.n2144 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2144 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2144 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2144 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2144 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2144 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2144 [6], \oc8051_golden_model_1.PSW_72 [7]);
  buf(\oc8051_golden_model_1.n2145 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2145 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2145 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2145 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2145 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2145 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2145 [7], \oc8051_golden_model_1.PSW_72 [7]);
  buf(\oc8051_golden_model_1.n2160 , \oc8051_golden_model_1.PSW_74 [0]);
  buf(\oc8051_golden_model_1.n2161 [0], \oc8051_golden_model_1.PSW_74 [0]);
  buf(\oc8051_golden_model_1.n2161 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2161 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2161 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2161 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2161 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2161 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2161 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2200 , \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2201 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2201 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2201 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2201 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2201 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2201 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2201 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2201 [7], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2202 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2202 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2202 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2202 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2202 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2202 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2202 [6], \oc8051_golden_model_1.n2203 [7]);
  buf(\oc8051_golden_model_1.n2203 [0], \oc8051_golden_model_1.PSW_0a [0]);
  buf(\oc8051_golden_model_1.n2203 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2203 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2203 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2203 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2203 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2203 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2210 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2210 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2210 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2210 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2211 , \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2212 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2212 [2], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2212 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2212 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2212 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2212 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2212 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2213 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2213 [1], \oc8051_golden_model_1.n2229 [2]);
  buf(\oc8051_golden_model_1.n2213 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2213 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2213 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2213 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2213 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2228 , \oc8051_golden_model_1.n2229 [0]);
  buf(\oc8051_golden_model_1.n2229 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2229 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2229 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2229 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2229 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2229 [7], 1'b0);
  buf(\oc8051_top_1.sub_result [0], ABINPUT[27]);
  buf(\oc8051_top_1.sub_result [1], ABINPUT[28]);
  buf(\oc8051_top_1.sub_result [2], ABINPUT[29]);
  buf(\oc8051_top_1.sub_result [3], ABINPUT[30]);
  buf(\oc8051_top_1.sub_result [4], ABINPUT[31]);
  buf(\oc8051_top_1.sub_result [5], ABINPUT[32]);
  buf(\oc8051_top_1.sub_result [6], ABINPUT[33]);
  buf(\oc8051_top_1.sub_result [7], ABINPUT[34]);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.ABINPUT [9], ABINPUT[9]);
  buf(\oc8051_top_1.ABINPUT [10], ABINPUT[10]);
  buf(\oc8051_top_1.ABINPUT [11], ABINPUT[11]);
  buf(\oc8051_top_1.ABINPUT [12], ABINPUT[12]);
  buf(\oc8051_top_1.ABINPUT [13], ABINPUT[13]);
  buf(\oc8051_top_1.ABINPUT [14], ABINPUT[14]);
  buf(\oc8051_top_1.ABINPUT [15], ABINPUT[15]);
  buf(\oc8051_top_1.ABINPUT [16], ABINPUT[16]);
  buf(\oc8051_top_1.ABINPUT [17], ABINPUT[17]);
  buf(\oc8051_top_1.ABINPUT [18], ABINPUT[18]);
  buf(\oc8051_top_1.ABINPUT [19], ABINPUT[19]);
  buf(\oc8051_top_1.ABINPUT [20], ABINPUT[20]);
  buf(\oc8051_top_1.ABINPUT [21], ABINPUT[21]);
  buf(\oc8051_top_1.ABINPUT [22], ABINPUT[22]);
  buf(\oc8051_top_1.ABINPUT [23], ABINPUT[23]);
  buf(\oc8051_top_1.ABINPUT [24], ABINPUT[24]);
  buf(\oc8051_top_1.ABINPUT [25], ABINPUT[25]);
  buf(\oc8051_top_1.ABINPUT [26], ABINPUT[26]);
  buf(\oc8051_top_1.ABINPUT [27], ABINPUT[27]);
  buf(\oc8051_top_1.ABINPUT [28], ABINPUT[28]);
  buf(\oc8051_top_1.ABINPUT [29], ABINPUT[29]);
  buf(\oc8051_top_1.ABINPUT [30], ABINPUT[30]);
  buf(\oc8051_top_1.ABINPUT [31], ABINPUT[31]);
  buf(\oc8051_top_1.ABINPUT [32], ABINPUT[32]);
  buf(\oc8051_top_1.ABINPUT [33], ABINPUT[33]);
  buf(\oc8051_top_1.ABINPUT [34], ABINPUT[34]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.desOv , ABINPUT[2]);
  buf(\oc8051_top_1.desAc , ABINPUT[1]);
  buf(\oc8051_top_1.desCy , ABINPUT[0]);
  buf(\oc8051_top_1.des2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.des2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.des2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.des2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.des2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.des2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.des2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.des2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.des1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.des1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.des1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.des1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.des1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.des1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.des1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.des1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.wr_dat [0], ABINPUT[3]);
  buf(\oc8051_top_1.wr_dat [1], ABINPUT[4]);
  buf(\oc8051_top_1.wr_dat [2], ABINPUT[5]);
  buf(\oc8051_top_1.wr_dat [3], ABINPUT[6]);
  buf(\oc8051_top_1.wr_dat [4], ABINPUT[7]);
  buf(\oc8051_top_1.wr_dat [5], ABINPUT[8]);
  buf(\oc8051_top_1.wr_dat [6], ABINPUT[9]);
  buf(\oc8051_top_1.wr_dat [7], ABINPUT[10]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(IRAM_gm[0], ABINPUT009[0]);
  buf(IRAM_gm[1], ABINPUT009[1]);
  buf(IRAM_gm[2], ABINPUT009[2]);
  buf(IRAM_gm[3], ABINPUT009[3]);
  buf(IRAM_gm[4], ABINPUT009[4]);
  buf(IRAM_gm[5], ABINPUT009[5]);
  buf(IRAM_gm[6], ABINPUT009[6]);
  buf(IRAM_gm[7], ABINPUT009[7]);
  buf(IRAM_gm[8], ABINPUT009[8]);
  buf(IRAM_gm[9], ABINPUT009[9]);
  buf(IRAM_gm[10], ABINPUT009[10]);
  buf(IRAM_gm[11], ABINPUT009[11]);
  buf(IRAM_gm[12], ABINPUT009[12]);
  buf(IRAM_gm[13], ABINPUT009[13]);
  buf(IRAM_gm[14], ABINPUT009[14]);
  buf(IRAM_gm[15], ABINPUT009[15]);
  buf(IRAM_gm[16], ABINPUT009[16]);
  buf(IRAM_gm[17], ABINPUT009[17]);
  buf(IRAM_gm[18], ABINPUT009[18]);
  buf(IRAM_gm[19], ABINPUT009[19]);
  buf(IRAM_gm[20], ABINPUT009[20]);
  buf(IRAM_gm[21], ABINPUT009[21]);
  buf(IRAM_gm[22], ABINPUT009[22]);
  buf(IRAM_gm[23], ABINPUT009[23]);
  buf(IRAM_gm[24], ABINPUT009[24]);
  buf(IRAM_gm[25], ABINPUT009[25]);
  buf(IRAM_gm[26], ABINPUT009[26]);
  buf(IRAM_gm[27], ABINPUT009[27]);
  buf(IRAM_gm[28], ABINPUT009[28]);
  buf(IRAM_gm[29], ABINPUT009[29]);
  buf(IRAM_gm[30], ABINPUT009[30]);
  buf(IRAM_gm[31], ABINPUT009[31]);
  buf(IRAM_gm[32], ABINPUT009[32]);
  buf(IRAM_gm[33], ABINPUT009[33]);
  buf(IRAM_gm[34], ABINPUT009[34]);
  buf(IRAM_gm[35], ABINPUT009[35]);
  buf(IRAM_gm[36], ABINPUT009[36]);
  buf(IRAM_gm[37], ABINPUT009[37]);
  buf(IRAM_gm[38], ABINPUT009[38]);
  buf(IRAM_gm[39], ABINPUT009[39]);
  buf(IRAM_gm[40], ABINPUT009[40]);
  buf(IRAM_gm[41], ABINPUT009[41]);
  buf(IRAM_gm[42], ABINPUT009[42]);
  buf(IRAM_gm[43], ABINPUT009[43]);
  buf(IRAM_gm[44], ABINPUT009[44]);
  buf(IRAM_gm[45], ABINPUT009[45]);
  buf(IRAM_gm[46], ABINPUT009[46]);
  buf(IRAM_gm[47], ABINPUT009[47]);
  buf(IRAM_gm[48], ABINPUT009[48]);
  buf(IRAM_gm[49], ABINPUT009[49]);
  buf(IRAM_gm[50], ABINPUT009[50]);
  buf(IRAM_gm[51], ABINPUT009[51]);
  buf(IRAM_gm[52], ABINPUT009[52]);
  buf(IRAM_gm[53], ABINPUT009[53]);
  buf(IRAM_gm[54], ABINPUT009[54]);
  buf(IRAM_gm[55], ABINPUT009[55]);
  buf(IRAM_gm[56], ABINPUT009[56]);
  buf(IRAM_gm[57], ABINPUT009[57]);
  buf(IRAM_gm[58], ABINPUT009[58]);
  buf(IRAM_gm[59], ABINPUT009[59]);
  buf(IRAM_gm[60], ABINPUT009[60]);
  buf(IRAM_gm[61], ABINPUT009[61]);
  buf(IRAM_gm[62], ABINPUT009[62]);
  buf(IRAM_gm[63], ABINPUT009[63]);
  buf(IRAM_gm[64], ABINPUT009[64]);
  buf(IRAM_gm[65], ABINPUT009[65]);
  buf(IRAM_gm[66], ABINPUT009[66]);
  buf(IRAM_gm[67], ABINPUT009[67]);
  buf(IRAM_gm[68], ABINPUT009[68]);
  buf(IRAM_gm[69], ABINPUT009[69]);
  buf(IRAM_gm[70], ABINPUT009[70]);
  buf(IRAM_gm[71], ABINPUT009[71]);
  buf(IRAM_gm[72], ABINPUT009[72]);
  buf(IRAM_gm[73], ABINPUT009[73]);
  buf(IRAM_gm[74], ABINPUT009[74]);
  buf(IRAM_gm[75], ABINPUT009[75]);
  buf(IRAM_gm[76], ABINPUT009[76]);
  buf(IRAM_gm[77], ABINPUT009[77]);
  buf(IRAM_gm[78], ABINPUT009[78]);
  buf(IRAM_gm[79], ABINPUT009[79]);
  buf(IRAM_gm[80], ABINPUT009[80]);
  buf(IRAM_gm[81], ABINPUT009[81]);
  buf(IRAM_gm[82], ABINPUT009[82]);
  buf(IRAM_gm[83], ABINPUT009[83]);
  buf(IRAM_gm[84], ABINPUT009[84]);
  buf(IRAM_gm[85], ABINPUT009[85]);
  buf(IRAM_gm[86], ABINPUT009[86]);
  buf(IRAM_gm[87], ABINPUT009[87]);
  buf(IRAM_gm[88], ABINPUT009[88]);
  buf(IRAM_gm[89], ABINPUT009[89]);
  buf(IRAM_gm[90], ABINPUT009[90]);
  buf(IRAM_gm[91], ABINPUT009[91]);
  buf(IRAM_gm[92], ABINPUT009[92]);
  buf(IRAM_gm[93], ABINPUT009[93]);
  buf(IRAM_gm[94], ABINPUT009[94]);
  buf(IRAM_gm[95], ABINPUT009[95]);
  buf(IRAM_gm[96], ABINPUT009[96]);
  buf(IRAM_gm[97], ABINPUT009[97]);
  buf(IRAM_gm[98], ABINPUT009[98]);
  buf(IRAM_gm[99], ABINPUT009[99]);
  buf(IRAM_gm[100], ABINPUT009[100]);
  buf(IRAM_gm[101], ABINPUT009[101]);
  buf(IRAM_gm[102], ABINPUT009[102]);
  buf(IRAM_gm[103], ABINPUT009[103]);
  buf(IRAM_gm[104], ABINPUT009[104]);
  buf(IRAM_gm[105], ABINPUT009[105]);
  buf(IRAM_gm[106], ABINPUT009[106]);
  buf(IRAM_gm[107], ABINPUT009[107]);
  buf(IRAM_gm[108], ABINPUT009[108]);
  buf(IRAM_gm[109], ABINPUT009[109]);
  buf(IRAM_gm[110], ABINPUT009[110]);
  buf(IRAM_gm[111], ABINPUT009[111]);
  buf(IRAM_gm[112], ABINPUT009[112]);
  buf(IRAM_gm[113], ABINPUT009[113]);
  buf(IRAM_gm[114], ABINPUT009[114]);
  buf(IRAM_gm[115], ABINPUT009[115]);
  buf(IRAM_gm[116], ABINPUT009[116]);
  buf(IRAM_gm[117], ABINPUT009[117]);
  buf(IRAM_gm[118], ABINPUT009[118]);
  buf(IRAM_gm[119], ABINPUT009[119]);
  buf(IRAM_gm[120], ABINPUT009[120]);
  buf(IRAM_gm[121], ABINPUT009[121]);
  buf(IRAM_gm[122], ABINPUT009[122]);
  buf(IRAM_gm[123], ABINPUT009[123]);
  buf(IRAM_gm[124], ABINPUT009[124]);
  buf(IRAM_gm[125], ABINPUT009[125]);
  buf(IRAM_gm[126], ABINPUT009[126]);
  buf(IRAM_gm[127], ABINPUT009[127]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm_next[0], ABINPUT008[0]);
  buf(PSW_gm_next[1], ABINPUT008[1]);
  buf(PSW_gm_next[2], ABINPUT008[2]);
  buf(PSW_gm_next[3], ABINPUT008[3]);
  buf(PSW_gm_next[4], ABINPUT008[4]);
  buf(PSW_gm_next[5], ABINPUT008[5]);
  buf(PSW_gm_next[6], ABINPUT008[6]);
  buf(PSW_gm_next[7], ABINPUT008[7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
