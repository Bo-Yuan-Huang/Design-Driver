module oc8051_symbolic_cxrom(
    clk,
    rst,
    word_in,
    cxrom_addr,
    pc1,
    pc2,
    cxrom_data_out,
    op_valid,
    op_out
);
    input clk, rst;
    input [31:0] word_in;
    input [15:0] cxrom_addr;
    input [15:0] pc1;
    input [15:0] pc2;

    output [31:0] cxrom_data_out;
    output op_valid;
    output [7:0] op_out;

    reg [7:0] regarray [15:0];
    reg [15:0] regvalid;

    wire [15:0] regvalid_ormask;

    wire [3:0] addr0 = cxrom_addr[3:0];
    wire [3:0] addr1 = cxrom_addr[3:0] + 1;
    wire [3:0] addr2 = cxrom_addr[3:0] + 2;
    wire [3:0] addr3 = cxrom_addr[3:0] + 3;

    assign regvalid_ormask = 
        addr0 == 0  ? 16'b0000000000001111 : 
        addr0 == 1  ? 16'b0000000000011110 : 
        addr0 == 2  ? 16'b0000000000111100 : 
        addr0 == 3  ? 16'b0000000001111000 : 
        addr0 == 4  ? 16'b0000000011110000 : 
        addr0 == 5  ? 16'b0000000111100000 : 
        addr0 == 6  ? 16'b0000001111000000 : 
        addr0 == 7  ? 16'b0000011110000000 : 
        addr0 == 8  ? 16'b0000111100000000 : 
        addr0 == 9  ? 16'b0001111000000000 : 
        addr0 == 10 ? 16'b0011110000000000 : 
        addr0 == 11 ? 16'b0111100000000000 : 
        addr0 == 12 ? 16'b1111000000000000 : 
        addr0 == 13 ? 16'b1110000000000001 : 
        addr0 == 14 ? 16'b1100000000000011 : 16'b1000000000000111;

    wire [15:0] regvalid_next;
    wire [7:0] bytein0 = word_in[7:0];
    wire [7:0] bytein1 = word_in[15:8];
    wire [7:0] bytein2 = word_in[23:16];
    wire [7:0] bytein3 = word_in[31:24];

    always @(posedge clk) begin
        if (rst) begin
            regvalid <= 16'b0;
        end
        else begin
            regvalid <= regvalid | regvalid_ormask;
            if (!regvalid[addr0])
                regarray[addr0] <= bytein0;
            if (!regvalid[addr1])
                regarray[addr1] <= bytein1;
            if (!regvalid[addr2])
                regarray[addr2] <= bytein2;
            if (!regvalid[addr3])
                regarray[addr3] <= bytein3;
        end
    end

    wire [7:0] byteout0 = regvalid[addr0] ? regarray[addr0] : bytein0;
    wire [7:0] byteout1 = regvalid[addr1] ? regarray[addr1] : bytein1;
    wire [7:0] byteout2 = regvalid[addr2] ? regarray[addr2] : bytein2;
    wire [7:0] byteout3 = regvalid[addr3] ? regarray[addr3] : bytein3;

    assign cxrom_data_out = { byteout3, byteout2, byteout1, byteout0 };
    
    wire [3:0] pc10 = pc1[3:0];
    wire [3:0] pc11 = pc1[3:0] + 1;
    wire [3:0] pc12 = pc1[3:0] + 2;
    wire [3:0] pc13 = pc1[3:0] + 3;
    wire pc1_valid = regvalid[pc10] && regvalid[pc11] && regvalid[pc12] && regvalid[pc13];

    wire [3:0] pc20 = pc2[3:0];
    wire [3:0] pc21 = pc2[3:0] + 1;
    wire [3:0] pc22 = pc2[3:0] + 2;
    wire [3:0] pc23 = pc2[3:0] + 3;
    wire pc2_valid = regvalid[pc20] && regvalid[pc21] && regvalid[pc22] && regvalid[pc23];

    assign op_valid = pc1_valid && pc2_valid;
    assign op_out = pc10 ? regarray[pc10] : 8'b0;
endmodule
