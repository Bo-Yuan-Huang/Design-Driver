
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire [15:0] _26822_;
  wire [7:0] _26823_;
  wire [7:0] _26824_;
  wire [7:0] _26825_;
  wire [7:0] _26826_;
  wire [7:0] _26827_;
  wire [7:0] _26828_;
  wire [7:0] _26829_;
  wire [7:0] _26830_;
  wire [7:0] _26831_;
  wire [7:0] _26832_;
  wire [7:0] _26833_;
  wire [7:0] _26834_;
  wire [7:0] _26835_;
  wire [7:0] _26836_;
  wire [7:0] _26837_;
  wire [7:0] _26838_;
  wire _26839_;
  wire [7:0] _26840_;
  wire [2:0] _26841_;
  wire [2:0] _26842_;
  wire [1:0] _26843_;
  wire [7:0] _26844_;
  wire _26845_;
  wire [1:0] _26846_;
  wire [1:0] _26847_;
  wire [2:0] _26848_;
  wire [2:0] _26849_;
  wire [1:0] _26850_;
  wire [3:0] _26851_;
  wire [1:0] _26852_;
  wire _26853_;
  wire [7:0] _26854_;
  wire [7:0] _26855_;
  wire [7:0] _26856_;
  wire [7:0] _26857_;
  wire [7:0] _26858_;
  wire [7:0] _26859_;
  wire [7:0] _26860_;
  wire [7:0] _26861_;
  wire [15:0] _26862_;
  wire [15:0] _26863_;
  wire _26864_;
  wire [4:0] _26865_;
  wire [7:0] _26866_;
  wire [7:0] _26867_;
  wire _26868_;
  wire _26869_;
  wire [15:0] _26870_;
  wire [15:0] _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire [7:0] _26875_;
  wire [2:0] _26876_;
  wire [7:0] _26877_;
  wire _26878_;
  wire [7:0] _26879_;
  wire _26880_;
  wire _26881_;
  wire [3:0] _26882_;
  wire [31:0] _26883_;
  wire [31:0] _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire [15:0] _26888_;
  wire _26889_;
  wire _26890_;
  wire [7:0] _26891_;
  wire _26892_;
  wire [2:0] _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire [7:0] _27313_;
  wire _27314_;
  wire [3:0] _27315_;
  wire _27316_;
  wire _27317_;
  wire [7:0] _27318_;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not (_22731_, rst);
  not (_22732_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  nor (_22733_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_22734_, _22733_, _22732_);
  not (_22735_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_22736_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_22737_, _22736_, _22735_);
  and (_22738_, _22737_, _22734_);
  and (_22740_, _22738_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_22741_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_22742_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_22744_, _22740_, _22742_);
  or (_22745_, _22744_, _22741_);
  and (_26863_[0], _22745_, _22731_);
  and (_22746_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_22747_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_22749_, _22740_, _22747_);
  or (_22750_, _22749_, _22746_);
  and (_26863_[1], _22750_, _22731_);
  and (_22751_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_22752_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_22753_, _22740_, _22752_);
  or (_22755_, _22753_, _22751_);
  and (_26863_[2], _22755_, _22731_);
  and (_22757_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_22758_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_22759_, _22740_, _22758_);
  or (_22760_, _22759_, _22757_);
  and (_26863_[3], _22760_, _22731_);
  or (_22761_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  not (_22762_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_22763_, _22740_, _22762_);
  and (_22764_, _22763_, _22731_);
  and (_26863_[4], _22764_, _22761_);
  or (_22766_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  not (_22767_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_22768_, _22740_, _22767_);
  and (_22769_, _22768_, _22731_);
  and (_26863_[5], _22769_, _22766_);
  or (_22771_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not (_22772_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_22773_, _22740_, _22772_);
  and (_22774_, _22773_, _22731_);
  and (_26863_[6], _22774_, _22771_);
  and (_22775_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_22776_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_22777_, _22740_, _22776_);
  or (_22778_, _22777_, _22775_);
  and (_26863_[7], _22778_, _22731_);
  or (_22779_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  not (_22780_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_22781_, _22740_, _22780_);
  and (_22782_, _22781_, _22731_);
  and (_26863_[8], _22782_, _22779_);
  and (_22783_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  not (_22784_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_22785_, _22740_, _22784_);
  or (_22786_, _22785_, _22783_);
  and (_26863_[9], _22786_, _22731_);
  or (_22788_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  not (_22789_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_22790_, _22740_, _22789_);
  and (_22791_, _22790_, _22731_);
  and (_26863_[10], _22791_, _22788_);
  or (_22792_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  not (_22793_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_22794_, _22740_, _22793_);
  and (_22795_, _22794_, _22731_);
  and (_26863_[11], _22795_, _22792_);
  or (_22796_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not (_22797_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_22799_, _22740_, _22797_);
  and (_22800_, _22799_, _22731_);
  and (_26863_[12], _22800_, _22796_);
  and (_22801_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not (_22802_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_22803_, _22740_, _22802_);
  or (_22804_, _22803_, _22801_);
  and (_26863_[13], _22804_, _22731_);
  or (_22805_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not (_22806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_22808_, _22740_, _22806_);
  and (_22809_, _22808_, _22731_);
  and (_26863_[14], _22809_, _22805_);
  and (_22810_, \oc8051_top_1.oc8051_decoder1.wr , _22735_);
  not (_22811_, _22810_);
  not (_22812_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22813_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _22735_);
  and (_22814_, _22813_, _22812_);
  and (_22815_, _22814_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_22816_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_22817_, _22816_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_22818_, _22817_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_22820_, _22818_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_22821_, _22820_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_22822_, _22821_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_22823_, _22822_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_22824_, _22822_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_22825_, _22824_, _22823_);
  and (_22826_, _22825_, _22815_);
  not (_22827_, _22826_);
  and (_22828_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_22829_, _22828_, _22813_);
  not (_22830_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_22831_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _22735_);
  and (_22832_, _22831_, _22830_);
  and (_22833_, _22832_, _22812_);
  and (_22834_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_22835_, _22834_, _22829_);
  nor (_22836_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_22837_, _22836_, _22813_);
  and (_22838_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_22839_, _22832_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_22840_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_22841_, _22840_, _22838_);
  and (_22843_, _22841_, _22835_);
  nand (_22844_, _22843_, _22827_);
  not (_22845_, _22844_);
  nor (_22846_, _22845_, _22814_);
  nor (_22847_, _22846_, _22811_);
  not (_22849_, _22847_);
  and (_22850_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_22851_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_22852_, _22851_, _22850_);
  not (_22853_, _22818_);
  not (_22854_, _22815_);
  nor (_22855_, _22817_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_22856_, _22855_, _22854_);
  and (_22857_, _22856_, _22853_);
  and (_22858_, _22836_, _22830_);
  nor (_22859_, _22858_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_22861_, _22859_);
  and (_22862_, _22861_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_22863_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_22864_, _22863_, _22862_);
  not (_22865_, _22864_);
  nor (_22866_, _22865_, _22857_);
  and (_22867_, _22866_, _22852_);
  not (_22868_, _22867_);
  not (_22869_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_22871_, _22844_, _22869_);
  and (_22872_, _22871_, _22868_);
  not (_22874_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_22875_, _22815_, _22874_);
  and (_22876_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_22877_, _22876_, _22875_);
  and (_22878_, _22861_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  not (_22880_, _22878_);
  and (_22881_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_22882_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_22884_, _22882_, _22881_);
  and (_22885_, _22884_, _22880_);
  and (_22886_, _22885_, _22877_);
  nor (_22887_, _22886_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_22888_, _22887_, _22872_);
  nor (_22890_, _22888_, _22849_);
  nor (_22891_, _22818_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_22893_, _22891_);
  nor (_22894_, _22854_, _22820_);
  and (_22896_, _22894_, _22893_);
  and (_22897_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor (_22898_, _22897_, _22896_);
  and (_22899_, _22861_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_22900_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_22901_, _22900_, _22899_);
  and (_22902_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_22903_, _22902_, _22829_);
  and (_22904_, _22903_, _22901_);
  and (_22905_, _22904_, _22898_);
  not (_22906_, _22905_);
  and (_22907_, _22906_, _22871_);
  and (_22908_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  nor (_22909_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_22910_, _22909_, _22816_);
  and (_22911_, _22910_, _22815_);
  nor (_22912_, _22911_, _22908_);
  and (_22913_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and (_22914_, _22861_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_22916_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_22917_, _22916_, _22914_);
  nor (_22918_, _22917_, _22913_);
  and (_22919_, _22918_, _22912_);
  nor (_22920_, _22919_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_22921_, _22920_, _22907_);
  nor (_22922_, _22921_, _22849_);
  nor (_22923_, _22922_, _22890_);
  nor (_22924_, _22820_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_22925_, _22924_);
  nor (_22926_, _22854_, _22821_);
  and (_22927_, _22926_, _22925_);
  not (_22928_, _22927_);
  and (_22930_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  nor (_22931_, _22930_, _22829_);
  and (_22932_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_22933_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_22934_, _22933_, _22932_);
  and (_22935_, _22934_, _22931_);
  and (_22936_, _22935_, _22928_);
  not (_22937_, _22936_);
  and (_22938_, _22937_, _22871_);
  nor (_22940_, _22816_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_22941_, _22940_, _22817_);
  and (_22942_, _22941_, _22815_);
  and (_22943_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_22945_, _22943_, _22942_);
  and (_22946_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_22947_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and (_22948_, _22861_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_22949_, _22948_, _22947_);
  nor (_22950_, _22949_, _22946_);
  and (_22951_, _22950_, _22945_);
  nor (_22952_, _22951_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_22953_, _22952_, _22938_);
  nor (_22954_, _22953_, _22849_);
  nor (_22956_, _22821_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_22957_, _22956_);
  nor (_22958_, _22854_, _22822_);
  and (_22960_, _22958_, _22957_);
  not (_22961_, _22960_);
  and (_22962_, _22837_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  nor (_22963_, _22962_, _22829_);
  and (_22964_, _22839_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and (_22965_, _22833_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_22966_, _22965_, _22964_);
  and (_22967_, _22966_, _22963_);
  and (_22968_, _22967_, _22961_);
  not (_22969_, _22968_);
  and (_22970_, _22969_, _22871_);
  nor (_22971_, _22871_, _22867_);
  nor (_22972_, _22971_, _22970_);
  and (_22973_, _22972_, _22954_);
  and (_22974_, _22973_, _22923_);
  nor (_22975_, _22905_, _22871_);
  and (_22976_, _22975_, _22847_);
  and (_22977_, _22976_, _22936_);
  and (_22978_, _22810_, _22869_);
  not (_22979_, _22978_);
  or (_22980_, _22979_, _22968_);
  nor (_22981_, _22980_, _22844_);
  and (_22982_, _22981_, _22977_);
  and (_22983_, _22982_, _22974_);
  not (_22984_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  nor (_22985_, _22984_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  not (_22986_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_22987_, _22986_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_22988_, _22987_, _22985_);
  and (_22989_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _22735_);
  and (_22990_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _22735_);
  nor (_22991_, _22990_, _22989_);
  not (_22992_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_22993_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _22735_);
  and (_22994_, _22993_, _22992_);
  and (_22995_, _22994_, _22991_);
  not (_22996_, _22995_);
  not (_22997_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_22998_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  not (_22999_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_23000_, _22999_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_23001_, _23000_, _22998_);
  or (_23002_, _23001_, _22997_);
  not (_23003_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_23004_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  nand (_23005_, _23004_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_23006_, _23005_, _23003_);
  and (_23007_, _23006_, _23002_);
  not (_23008_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  or (_23009_, _23000_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_23010_, _23009_, _23008_);
  not (_23011_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  or (_23012_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_23013_, _23012_, _22999_);
  or (_23015_, _23013_, _23011_);
  and (_23016_, _23015_, _23010_);
  and (_23017_, _23016_, _23007_);
  or (_23018_, _23012_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or (_23019_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  not (_23020_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23022_, _23020_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  and (_23023_, _23022_, _23019_);
  not (_23024_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_23025_, _23024_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or (_23026_, _23025_, _23023_);
  nand (_23027_, _23024_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or (_23028_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_23029_, _23028_, _23026_);
  or (_23030_, _23029_, _23018_);
  and (_23031_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_23032_, _23031_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_23033_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  not (_23034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand (_23035_, _23031_, _22998_);
  or (_23036_, _23035_, _23034_);
  and (_23037_, _23036_, _23033_);
  and (_23038_, _23037_, _23030_);
  and (_23039_, _23038_, _23017_);
  or (_23040_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_23041_, _23040_, _23029_);
  and (_23042_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_23043_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not (_23044_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_23045_, _23044_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  nor (_23047_, _23045_, _23034_);
  nor (_23048_, _23047_, _23043_);
  and (_23049_, _23048_, _23041_);
  not (_23050_, _23049_);
  and (_23051_, _23050_, _23039_);
  nor (_23052_, _23049_, _23039_);
  and (_23053_, _23049_, _23039_);
  nor (_23054_, _23053_, _23052_);
  not (_23055_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_23056_, _23001_, _23055_);
  not (_23057_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_23058_, _23005_, _23057_);
  and (_23059_, _23058_, _23056_);
  not (_23060_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or (_23061_, _23013_, _23060_);
  not (_23062_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or (_23063_, _23009_, _23062_);
  and (_23064_, _23063_, _23061_);
  and (_23065_, _23064_, _23059_);
  or (_23066_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23067_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _23020_);
  and (_23068_, _23067_, _23066_);
  or (_23069_, _23068_, _23025_);
  or (_23070_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_23071_, _23070_, _23069_);
  or (_23072_, _23071_, _23018_);
  nand (_23073_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  not (_23074_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_23075_, _23035_, _23074_);
  and (_23076_, _23075_, _23073_);
  and (_23078_, _23076_, _23072_);
  and (_23079_, _23078_, _23065_);
  or (_23080_, _23071_, _23040_);
  nand (_23081_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or (_23082_, _23045_, _23074_);
  and (_23083_, _23082_, _23081_);
  nand (_23084_, _23083_, _23080_);
  nor (_23085_, _23084_, _23079_);
  not (_23086_, _23084_);
  nor (_23087_, _23086_, _23079_);
  and (_23088_, _23086_, _23079_);
  nor (_23089_, _23088_, _23087_);
  not (_23090_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_23091_, _23001_, _23090_);
  not (_23092_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_23093_, _23005_, _23092_);
  and (_23094_, _23093_, _23091_);
  not (_23095_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  or (_23096_, _23013_, _23095_);
  not (_23097_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or (_23098_, _23009_, _23097_);
  and (_23099_, _23098_, _23096_);
  and (_23100_, _23099_, _23094_);
  or (_23101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23103_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _23020_);
  and (_23104_, _23103_, _23101_);
  or (_23105_, _23104_, _23025_);
  or (_23106_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_23107_, _23106_, _23105_);
  or (_23108_, _23107_, _23018_);
  not (_23109_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_23111_, _23035_, _23109_);
  nand (_23112_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_23113_, _23112_, _23111_);
  and (_23114_, _23113_, _23108_);
  nand (_23115_, _23114_, _23100_);
  or (_23116_, _23107_, _23040_);
  nand (_23117_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  or (_23118_, _23045_, _23109_);
  and (_23119_, _23118_, _23117_);
  and (_23120_, _23119_, _23116_);
  and (_23121_, _23120_, _23115_);
  nand (_23122_, _23119_, _23116_);
  and (_23123_, _23122_, _23115_);
  nor (_23124_, _23122_, _23115_);
  nor (_23125_, _23124_, _23123_);
  not (_23126_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_23127_, _23001_, _23126_);
  not (_23128_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_23129_, _23005_, _23128_);
  and (_23130_, _23129_, _23127_);
  not (_23131_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  or (_23132_, _23013_, _23131_);
  not (_23133_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or (_23134_, _23009_, _23133_);
  and (_23136_, _23134_, _23132_);
  and (_23137_, _23136_, _23130_);
  or (_23138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23139_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _23020_);
  and (_23140_, _23139_, _23138_);
  or (_23141_, _23140_, _23025_);
  or (_23142_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_23143_, _23142_, _23141_);
  or (_23144_, _23143_, _23018_);
  not (_23145_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_23146_, _23035_, _23145_);
  nand (_23147_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and (_23148_, _23147_, _23146_);
  and (_23149_, _23148_, _23144_);
  and (_23150_, _23149_, _23137_);
  or (_23151_, _23143_, _23040_);
  nand (_23152_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  or (_23154_, _23045_, _23145_);
  and (_23155_, _23154_, _23152_);
  nand (_23156_, _23155_, _23151_);
  and (_23157_, _23156_, _23150_);
  nor (_23158_, _23157_, _23125_);
  nor (_23159_, _23158_, _23121_);
  nor (_23160_, _23159_, _23089_);
  nor (_23161_, _23160_, _23085_);
  and (_23162_, _23159_, _23089_);
  nor (_23163_, _23162_, _23160_);
  not (_23164_, _23163_);
  and (_23166_, _23157_, _23125_);
  nor (_23167_, _23166_, _23158_);
  not (_23168_, _23167_);
  and (_23169_, _23155_, _23151_);
  nor (_23170_, _23169_, _23150_);
  and (_23172_, _23169_, _23150_);
  nor (_23173_, _23172_, _23170_);
  not (_23174_, _23173_);
  not (_23175_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  or (_23176_, _23001_, _23175_);
  not (_23177_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_23178_, _23005_, _23177_);
  and (_23179_, _23178_, _23176_);
  not (_23181_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or (_23182_, _23013_, _23181_);
  not (_23183_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or (_23184_, _23009_, _23183_);
  and (_23185_, _23184_, _23182_);
  and (_23186_, _23185_, _23179_);
  or (_23187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23188_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _23020_);
  and (_23189_, _23188_, _23187_);
  or (_23190_, _23189_, _23025_);
  or (_23191_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_23192_, _23191_, _23190_);
  or (_23193_, _23192_, _23018_);
  nand (_23194_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  not (_23195_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_23196_, _23035_, _23195_);
  and (_23197_, _23196_, _23194_);
  and (_23198_, _23197_, _23193_);
  and (_23199_, _23198_, _23186_);
  or (_23201_, _23192_, _23040_);
  nand (_23202_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  or (_23203_, _23045_, _23195_);
  and (_23204_, _23203_, _23202_);
  and (_23205_, _23204_, _23201_);
  and (_23206_, _23205_, _23199_);
  nor (_23207_, _23205_, _23199_);
  nor (_23208_, _23207_, _23206_);
  nand (_23209_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  not (_23210_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_23211_, _23035_, _23210_);
  and (_23212_, _23211_, _23209_);
  not (_23213_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_23214_, _23001_, _23213_);
  not (_23215_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_23216_, _23005_, _23215_);
  and (_23217_, _23216_, _23214_);
  and (_23218_, _23217_, _23212_);
  or (_23219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23220_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _23020_);
  and (_23221_, _23220_, _23219_);
  or (_23222_, _23221_, _23025_);
  or (_23223_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_23224_, _23223_, _23222_);
  or (_23225_, _23224_, _23018_);
  not (_23226_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_23227_, _23009_, _23226_);
  not (_23228_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  or (_23229_, _23013_, _23228_);
  and (_23230_, _23229_, _23227_);
  and (_23231_, _23230_, _23225_);
  nand (_23232_, _23231_, _23218_);
  or (_23233_, _23224_, _23040_);
  nand (_23234_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_23235_, _23045_, _23210_);
  and (_23236_, _23235_, _23234_);
  nand (_23237_, _23236_, _23233_);
  and (_23238_, _23237_, _23232_);
  nor (_23239_, _23237_, _23232_);
  nor (_23240_, _23239_, _23238_);
  not (_23241_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_23242_, _23001_, _23241_);
  not (_23243_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_23244_, _23005_, _23243_);
  and (_23245_, _23244_, _23242_);
  not (_23246_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  or (_23247_, _23013_, _23246_);
  not (_23248_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_23249_, _23009_, _23248_);
  and (_23250_, _23249_, _23247_);
  and (_23251_, _23250_, _23245_);
  or (_23252_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23253_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _23020_);
  and (_23254_, _23253_, _23252_);
  or (_23255_, _23254_, _23025_);
  or (_23256_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_23257_, _23256_, _23255_);
  or (_23258_, _23257_, _23018_);
  nand (_23259_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  not (_23260_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_23261_, _23035_, _23260_);
  and (_23262_, _23261_, _23259_);
  and (_23263_, _23262_, _23258_);
  nand (_23264_, _23263_, _23251_);
  or (_23265_, _23257_, _23040_);
  nand (_23266_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_23267_, _23045_, _23260_);
  and (_23268_, _23267_, _23266_);
  nand (_23269_, _23268_, _23265_);
  nor (_23270_, _23269_, _23264_);
  and (_23271_, _23269_, _23264_);
  nor (_23272_, _23271_, _23270_);
  not (_23273_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_23274_, _23001_, _23273_);
  not (_23275_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_23276_, _23005_, _23275_);
  nor (_23277_, _23276_, _23274_);
  not (_23278_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor (_23279_, _23013_, _23278_);
  not (_23280_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor (_23281_, _23009_, _23280_);
  nor (_23282_, _23281_, _23279_);
  and (_23283_, _23282_, _23277_);
  or (_23284_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  or (_23285_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _23020_);
  and (_23286_, _23285_, _23284_);
  or (_23287_, _23286_, _23025_);
  or (_23288_, _23027_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_23289_, _23288_, _23287_);
  or (_23290_, _23289_, _23018_);
  not (_23291_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_23292_, _23035_, _23291_);
  and (_23293_, _23032_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_23294_, _23293_, _23292_);
  and (_23295_, _23294_, _23290_);
  and (_23296_, _23295_, _23283_);
  or (_23297_, _23289_, _23040_);
  nand (_23298_, _23042_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  or (_23299_, _23045_, _23291_);
  and (_23300_, _23299_, _23298_);
  nand (_23301_, _23300_, _23297_);
  and (_23302_, _23301_, _23296_);
  nor (_23304_, _23302_, _23272_);
  not (_23305_, _23269_);
  and (_23306_, _23305_, _23264_);
  nor (_23308_, _23306_, _23304_);
  nor (_23309_, _23308_, _23240_);
  and (_23310_, _23236_, _23233_);
  and (_23311_, _23310_, _23232_);
  nor (_23312_, _23311_, _23309_);
  nor (_23313_, _23312_, _23208_);
  and (_23314_, _23312_, _23208_);
  nor (_23316_, _23314_, _23313_);
  and (_23317_, _23308_, _23240_);
  nor (_23318_, _23317_, _23309_);
  not (_23319_, _23318_);
  and (_23320_, _23302_, _23272_);
  nor (_23321_, _23320_, _23304_);
  not (_23322_, _23321_);
  not (_23323_, _23301_);
  nor (_23324_, _23323_, _23296_);
  and (_23325_, _23323_, _23296_);
  nor (_23327_, _23325_, _23324_);
  and (_23328_, _22984_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nand (_23329_, _23068_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23330_, _23221_, _22986_);
  nand (_23331_, _23330_, _23329_);
  nand (_23333_, _23331_, _23328_);
  and (_23334_, _22985_, _22986_);
  nand (_23335_, _23334_, _23254_);
  and (_23336_, _22985_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23337_, _23336_, _23104_);
  and (_23338_, _23337_, _23335_);
  and (_23340_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_23341_, _23340_, _22986_);
  nand (_23342_, _23341_, _23189_);
  and (_23343_, _23340_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23344_, _23343_, _23023_);
  and (_23345_, _23344_, _23342_);
  nor (_23346_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_23347_, _23346_, _22986_);
  nand (_23348_, _23347_, _23286_);
  and (_23349_, _23346_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand (_23350_, _23349_, _23140_);
  and (_23351_, _23350_, _23348_);
  and (_23352_, _23351_, _23345_);
  and (_23353_, _23352_, _23338_);
  nand (_23354_, _23353_, _23333_);
  nand (_23355_, _23354_, _23027_);
  and (_23356_, _23025_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not (_23357_, _23356_);
  and (_23358_, _23357_, _23355_);
  and (_23359_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_23360_, _23359_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nor (_23361_, _23360_, _23358_);
  not (_23362_, _23360_);
  and (_23363_, _23362_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_23364_, _23363_, _23361_);
  nor (_23366_, _23364_, _23327_);
  and (_23367_, _23366_, _23322_);
  and (_23368_, _23367_, _23319_);
  not (_23369_, _23368_);
  nor (_23370_, _23369_, _23316_);
  nand (_23371_, _23204_, _23201_);
  or (_23372_, _23371_, _23199_);
  and (_23373_, _23371_, _23199_);
  or (_23374_, _23312_, _23373_);
  and (_23375_, _23374_, _23372_);
  or (_23376_, _23375_, _23370_);
  and (_23377_, _23376_, _23174_);
  and (_23378_, _23377_, _23168_);
  and (_23379_, _23378_, _23164_);
  nor (_23380_, _23379_, _23161_);
  nor (_23381_, _23380_, _23054_);
  nor (_23382_, _23381_, _23051_);
  nor (_23383_, _23382_, _22996_);
  not (_23385_, _23383_);
  not (_23386_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_23387_, _22735_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_23388_, _23387_, _23386_);
  and (_23390_, _23388_, _22991_);
  not (_23391_, _23390_);
  not (_23392_, _23052_);
  not (_23393_, _23054_);
  not (_23395_, _23240_);
  and (_23396_, _23324_, _23272_);
  nor (_23397_, _23396_, _23271_);
  nor (_23398_, _23397_, _23395_);
  nor (_23399_, _23398_, _23238_);
  nor (_23400_, _23399_, _23208_);
  and (_23401_, _23399_, _23208_);
  nor (_23402_, _23401_, _23400_);
  not (_23403_, _23327_);
  nor (_23404_, _23364_, _23403_);
  and (_23405_, _23404_, _23272_);
  and (_23406_, _23397_, _23395_);
  nor (_23407_, _23406_, _23398_);
  and (_23408_, _23407_, _23405_);
  not (_23409_, _23408_);
  nor (_23410_, _23409_, _23402_);
  nor (_23411_, _23399_, _23206_);
  or (_23412_, _23411_, _23207_);
  or (_23413_, _23412_, _23410_);
  and (_23414_, _23413_, _23173_);
  and (_23415_, _23170_, _23125_);
  nor (_23416_, _23170_, _23125_);
  nor (_23417_, _23416_, _23415_);
  and (_23418_, _23417_, _23414_);
  not (_23419_, _23089_);
  nor (_23420_, _23415_, _23123_);
  nor (_23421_, _23420_, _23419_);
  and (_23422_, _23420_, _23419_);
  nor (_23423_, _23422_, _23421_);
  and (_23424_, _23423_, _23418_);
  not (_23425_, _23424_);
  nor (_23426_, _23421_, _23087_);
  and (_23427_, _23426_, _23425_);
  or (_23429_, _23427_, _23393_);
  and (_23430_, _23429_, _23392_);
  nor (_23432_, _23430_, _23391_);
  not (_23433_, _23363_);
  not (_23434_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_23436_, _22990_, _23434_);
  and (_23437_, _23436_, _22994_);
  and (_23438_, _23437_, _23433_);
  nor (_23439_, _23387_, _22993_);
  and (_23440_, _22989_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_23441_, _23440_, _23439_);
  and (_23442_, _23441_, _23363_);
  nor (_23443_, _23442_, _23438_);
  nor (_23444_, _23443_, _23361_);
  not (_23445_, _23444_);
  and (_23446_, _23433_, _23358_);
  not (_23447_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_23448_, _22989_, _23447_);
  and (_23449_, _23448_, _23388_);
  and (_23450_, _23439_, _23448_);
  not (_23451_, _23450_);
  nor (_23452_, _23451_, _23361_);
  nor (_23453_, _23452_, _23449_);
  nor (_23454_, _23453_, _23446_);
  not (_23455_, _23454_);
  not (_23456_, _23364_);
  not (_23457_, _23115_);
  and (_23458_, _23457_, _23079_);
  not (_23459_, _23458_);
  not (_23460_, _23150_);
  and (_23461_, _23436_, _23388_);
  nor (_23462_, _23264_, _23232_);
  nor (_23463_, _23462_, _23199_);
  and (_23464_, _23463_, _23461_);
  and (_23465_, _23464_, _23460_);
  nor (_23466_, _23465_, _23459_);
  nor (_23467_, _23466_, _23039_);
  nor (_23468_, _23467_, _23456_);
  not (_23469_, _23468_);
  not (_23470_, _23461_);
  not (_23471_, _23466_);
  nor (_23472_, _23364_, _23039_);
  and (_23473_, _23472_, _23471_);
  nor (_23474_, _23473_, _23470_);
  and (_23475_, _23474_, _23469_);
  nor (_23476_, _23362_, _23358_);
  and (_23477_, _23448_, _22994_);
  not (_23478_, _23358_);
  and (_23479_, _22993_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_23480_, _23479_, _23436_);
  and (_23481_, _23480_, _23478_);
  nor (_23482_, _23481_, _23477_);
  nor (_23483_, _23482_, _23476_);
  and (_23484_, _23439_, _22991_);
  and (_23485_, _23484_, _23456_);
  not (_23486_, _23485_);
  not (_23487_, _23039_);
  and (_23488_, _23479_, _23448_);
  and (_23489_, _23488_, _23487_);
  not (_23490_, _23489_);
  not (_23491_, _23296_);
  and (_23492_, _23440_, _23388_);
  and (_23493_, _23492_, _23491_);
  nor (_23494_, _23493_, _23464_);
  and (_23495_, _23494_, _23490_);
  nand (_23496_, _23495_, _23486_);
  or (_23497_, _23496_, _23483_);
  nor (_23498_, _23497_, _23475_);
  and (_23499_, _23498_, _23455_);
  and (_23500_, _23499_, _23445_);
  not (_23501_, _23500_);
  nor (_23503_, _23501_, _23432_);
  and (_23504_, _23503_, _23385_);
  nor (_23505_, _23504_, _22988_);
  and (_23506_, _23440_, _23479_);
  and (_23507_, _23506_, _23269_);
  and (_23508_, _23491_, _23264_);
  not (_23509_, _23264_);
  and (_23510_, _23296_, _23509_);
  nor (_23511_, _23510_, _23508_);
  not (_23512_, _23511_);
  nand (_23513_, _23512_, _23364_);
  and (_23514_, _23440_, _22994_);
  or (_23515_, _23512_, _23364_);
  and (_23516_, _23515_, _23514_);
  and (_23517_, _23516_, _23513_);
  nor (_23518_, _23517_, _23507_);
  and (_23519_, _23450_, _23272_);
  not (_23520_, _23449_);
  nor (_23521_, _23520_, _23270_);
  or (_23522_, _23521_, _23519_);
  not (_23523_, _23522_);
  and (_23524_, _23480_, _23271_);
  and (_23525_, _23437_, _23509_);
  nor (_23526_, _23525_, _23524_);
  and (_23527_, _23526_, _23523_);
  and (_23528_, _23439_, _23436_);
  not (_23529_, _23528_);
  and (_23530_, _23388_, _23434_);
  and (_23531_, _23479_, _22991_);
  nor (_23532_, _23531_, _23530_);
  and (_23533_, _23532_, _23529_);
  and (_23534_, _23440_, _23386_);
  and (_23535_, _23448_, _22993_);
  or (_23536_, _23535_, _23534_);
  nor (_23537_, _23536_, _23484_);
  and (_23538_, _23537_, _23533_);
  nor (_23539_, _23538_, _23509_);
  not (_23540_, _23539_);
  and (_23541_, _23540_, _23527_);
  and (_23542_, _23541_, _23518_);
  nor (_23543_, _23542_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23544_, _23334_, _22869_);
  and (_23545_, _23544_, _23254_);
  or (_23546_, _23545_, _23543_);
  or (_23547_, _23546_, _23505_);
  and (_23548_, _23547_, _22847_);
  and (_23549_, _23548_, _22983_);
  not (_23550_, _22983_);
  and (_23551_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  or (_03395_, _23551_, _23549_);
  nand (_23552_, _23340_, _22987_);
  nor (_23553_, _23552_, _23504_);
  and (_23554_, _23450_, _23208_);
  nor (_23555_, _23520_, _23206_);
  or (_23556_, _23555_, _23554_);
  and (_23557_, _23480_, _23207_);
  and (_23558_, _23437_, _23199_);
  nor (_23559_, _23558_, _23557_);
  not (_23560_, _23559_);
  nor (_23561_, _23560_, _23556_);
  nor (_23562_, _23538_, _23199_);
  not (_23563_, _23199_);
  nand (_23564_, _23508_, _23232_);
  or (_23565_, _23564_, _23456_);
  nand (_23566_, _23462_, _23296_);
  or (_23567_, _23566_, _23364_);
  nand (_23568_, _23567_, _23565_);
  nand (_23569_, _23568_, _23563_);
  or (_23570_, _23568_, _23563_);
  and (_23571_, _23570_, _23514_);
  nand (_23572_, _23571_, _23569_);
  and (_23573_, _23506_, _23371_);
  not (_23574_, _23573_);
  nand (_23575_, _23574_, _23572_);
  nor (_23576_, _23575_, _23562_);
  nand (_23577_, _23576_, _23561_);
  and (_23578_, _23577_, _22869_);
  nor (_23579_, _23341_, _22869_);
  and (_23580_, _23579_, _23189_);
  or (_23581_, _23580_, _23578_);
  or (_23582_, _23581_, _23553_);
  and (_23583_, _23582_, _22847_);
  and (_23584_, _23583_, _22983_);
  and (_23585_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  or (_04137_, _23585_, _23584_);
  and (_23586_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_23587_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_23588_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_23589_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_23590_, _23589_, _23588_);
  nand (_23591_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_23592_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_23593_, _23592_, _23588_);
  nand (_23594_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_23595_, _23594_, _23591_);
  nor (_23596_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_23597_, _23596_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nand (_23598_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  not (_23599_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_23600_, _23599_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_23601_, _23600_, _23588_);
  not (_23602_, _23601_);
  nand (_23603_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_23604_, _23603_, _23598_);
  nor (_23605_, _23589_, _23588_);
  nand (_23606_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_23607_, _23589_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_23608_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_23609_, _23608_, _23606_);
  and (_23610_, _23609_, _23604_);
  and (_23611_, _23610_, _23595_);
  or (_23612_, _23611_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_23613_, _23612_, _23587_);
  nor (_23614_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _23587_);
  or (_23615_, _23614_, _23613_);
  and (_23616_, _23615_, _22738_);
  not (_23617_, _23616_);
  not (_23618_, _22734_);
  nor (_23619_, _22737_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_23620_, _23619_, _23618_);
  nand (_23621_, _23620_, _23617_);
  not (_23622_, _22738_);
  not (_23623_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_23624_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and (_23625_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_23626_, _23625_, _23624_);
  nand (_23627_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand (_23628_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_23629_, _23628_, _23627_);
  nand (_23630_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nand (_23631_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_23632_, _23631_, _23630_);
  and (_23633_, _23632_, _23629_);
  nand (_23634_, _23633_, _23626_);
  nand (_23635_, _23634_, _23623_);
  nand (_23636_, _23635_, _23587_);
  nor (_23637_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _23587_);
  not (_23638_, _23637_);
  and (_23639_, _23638_, _23636_);
  or (_23640_, _23639_, _23622_);
  nor (_23641_, _22737_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_23642_, _23641_, _23618_);
  and (_23643_, _23642_, _23640_);
  and (_23644_, _23643_, _23621_);
  nand (_23645_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand (_23646_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nand (_23647_, _23646_, _23645_);
  and (_23648_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_23649_, _23648_, _23647_);
  nand (_23650_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_23651_, _23650_, _23623_);
  nand (_23652_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_23653_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_23654_, _23653_, _23652_);
  and (_23655_, _23654_, _23651_);
  nand (_23656_, _23655_, _23649_);
  or (_23657_, _23656_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_23658_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _23587_);
  not (_23659_, _23658_);
  and (_23660_, _23659_, _23657_);
  or (_23661_, _23660_, _23622_);
  nor (_23662_, _22737_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_23663_, _23662_, _23618_);
  and (_23664_, _23663_, _23661_);
  nand (_23665_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nand (_23666_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_23667_, _23666_, _23665_);
  nand (_23668_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_23669_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_23670_, _23669_, _23668_);
  nand (_23671_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nand (_23672_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_23673_, _23672_, _23671_);
  and (_23674_, _23673_, _23670_);
  and (_23675_, _23674_, _23667_);
  or (_23676_, _23675_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_23677_, _23676_, _23587_);
  nor (_23679_, _23587_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  not (_23680_, _23679_);
  and (_23681_, _23680_, _23677_);
  or (_23682_, _23681_, _23622_);
  nor (_23683_, _22737_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_23684_, _23683_, _23618_);
  and (_23685_, _23684_, _23682_);
  nor (_23686_, _23685_, _23664_);
  and (_23687_, _23686_, _23644_);
  and (_23688_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_23689_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_23690_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_23691_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_23692_, _23691_, _23690_);
  and (_23693_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_23694_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_23695_, _23694_, _23693_);
  nand (_23696_, _23695_, _23692_);
  or (_23697_, _23696_, _23689_);
  or (_23698_, _23697_, _23688_);
  or (_23699_, _23698_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_23700_, _23699_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_23701_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _23587_);
  not (_23702_, _23701_);
  and (_23703_, _23702_, _23700_);
  or (_23704_, _23703_, _23622_);
  nor (_23705_, _22737_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_23706_, _23705_, _23618_);
  and (_23707_, _23706_, _23704_);
  not (_23708_, _23707_);
  nand (_23709_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nand (_23710_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_23711_, _23710_, _23709_);
  nand (_23712_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_23713_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_23714_, _23713_, _23712_);
  nand (_23715_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_23716_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_23717_, _23716_, _23715_);
  and (_23718_, _23717_, _23714_);
  nand (_23719_, _23718_, _23711_);
  nand (_23720_, _23719_, _23623_);
  nand (_23721_, _23720_, _23587_);
  nor (_23722_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _23587_);
  not (_23723_, _23722_);
  and (_23724_, _23723_, _23721_);
  or (_23726_, _23724_, _23622_);
  nor (_23727_, _22737_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_23728_, _23727_, _23618_);
  and (_23729_, _23728_, _23726_);
  nand (_23730_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand (_23731_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_23732_, _23731_, _23730_);
  nand (_23733_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nand (_23734_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_23735_, _23734_, _23733_);
  and (_23736_, _23735_, _23732_);
  nand (_23737_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_23738_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_23739_, _23738_, _23737_);
  and (_23740_, _23739_, _23736_);
  or (_23741_, _23740_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_23742_, _23741_, _23587_);
  nor (_23743_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _23587_);
  not (_23744_, _23743_);
  and (_23745_, _23744_, _23742_);
  or (_23746_, _23745_, _23622_);
  nor (_23747_, _22737_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_23748_, _23747_, _23618_);
  nand (_23749_, _23748_, _23746_);
  nand (_23750_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nand (_23751_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_23752_, _23751_, _23750_);
  nand (_23753_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_23754_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_23755_, _23754_, _23753_);
  nand (_23756_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand (_23757_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_23758_, _23757_, _23756_);
  and (_23759_, _23758_, _23755_);
  nand (_23760_, _23759_, _23752_);
  and (_23761_, _23760_, _23623_);
  or (_23762_, _23761_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_23763_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _23587_);
  not (_23764_, _23763_);
  and (_23765_, _23764_, _23762_);
  or (_23766_, _23765_, _23622_);
  nor (_23767_, _22737_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_23768_, _23767_, _23618_);
  nand (_23769_, _23768_, _23766_);
  and (_23770_, _23769_, _23749_);
  and (_23771_, _23770_, _23729_);
  and (_23772_, _23771_, _23708_);
  and (_23773_, _23772_, _23687_);
  and (_23774_, _23773_, _22735_);
  or (_23775_, _23774_, _23586_);
  and (_23776_, _23775_, _22731_);
  not (_23777_, _23643_);
  and (_23778_, _23777_, _23621_);
  and (_23779_, _23778_, _23664_);
  and (_23780_, _23779_, _23685_);
  and (_23781_, _23768_, _23766_);
  and (_23782_, _23781_, _23729_);
  and (_23783_, _23782_, _23749_);
  and (_23784_, _23783_, _23707_);
  and (_23785_, _23784_, _23780_);
  and (_23786_, _23748_, _23746_);
  and (_23788_, _23782_, _23786_);
  and (_23789_, _23788_, _23707_);
  and (_23790_, _23789_, _23687_);
  not (_23791_, _23685_);
  and (_23792_, _23779_, _23791_);
  and (_23793_, _23792_, _23784_);
  or (_23794_, _23793_, _23790_);
  or (_23795_, _23794_, _23785_);
  not (_23796_, _23664_);
  and (_23797_, _23796_, _23644_);
  not (_23798_, _23729_);
  and (_23799_, _23749_, _23798_);
  and (_23800_, _23799_, _23769_);
  and (_23801_, _23800_, _23708_);
  and (_23802_, _23685_, _23796_);
  and (_23803_, _23802_, _23644_);
  and (_23804_, _23769_, _23786_);
  and (_23805_, _23804_, _23729_);
  and (_23806_, _23805_, _23707_);
  and (_23807_, _23806_, _23803_);
  or (_23808_, _23807_, _23801_);
  and (_23809_, _23808_, _23797_);
  and (_23810_, _23786_, _23798_);
  and (_23811_, _23810_, _23769_);
  and (_23812_, _23811_, _23707_);
  and (_23813_, _23664_, _23643_);
  and (_23814_, _23813_, _23621_);
  and (_23815_, _23814_, _23812_);
  and (_23816_, _23778_, _23686_);
  and (_23817_, _23816_, _23784_);
  and (_23818_, _23800_, _23707_);
  and (_23819_, _23818_, _23797_);
  or (_23820_, _23819_, _23817_);
  or (_23821_, _23820_, _23815_);
  or (_23822_, _23821_, _23809_);
  or (_23823_, _23822_, _23795_);
  not (_23824_, _23621_);
  and (_23825_, _23707_, _23824_);
  and (_23826_, _23825_, _23811_);
  or (_23827_, _23806_, _23800_);
  and (_23828_, _23827_, _23824_);
  nor (_23829_, _23828_, _23826_);
  and (_23830_, _23812_, _23779_);
  and (_23831_, _23792_, _23772_);
  or (_23832_, _23831_, _23830_);
  and (_23833_, _23812_, _23797_);
  nor (_23834_, _23833_, _23832_);
  nand (_23835_, _23834_, _23829_);
  and (_23836_, _23799_, _23780_);
  and (_23837_, _23836_, _23769_);
  nor (_23838_, _23707_, _23621_);
  and (_23839_, _23838_, _23805_);
  and (_23840_, _23814_, _23800_);
  and (_23841_, _23814_, _23805_);
  or (_23842_, _23841_, _23840_);
  or (_23843_, _23842_, _23839_);
  and (_23844_, _23805_, _23708_);
  and (_23845_, _23844_, _23803_);
  and (_23846_, _23806_, _23687_);
  or (_23847_, _23846_, _23845_);
  or (_23848_, _23847_, _23843_);
  or (_23850_, _23848_, _23837_);
  or (_23851_, _23850_, _23835_);
  or (_23853_, _23851_, _23823_);
  nor (_23854_, \oc8051_top_1.oc8051_sfr1.wait_data , rst);
  and (_23855_, _23854_, _22736_);
  and (_23856_, _23855_, _23853_);
  or (_26851_[2], _23856_, _23776_);
  nand (_23857_, _23328_, _22987_);
  nor (_23858_, _23857_, _23504_);
  and (_23859_, _23506_, _23237_);
  or (_23860_, _23510_, _23364_);
  or (_23861_, _23508_, _23456_);
  and (_23862_, _23861_, _23860_);
  nand (_23863_, _23862_, _23232_);
  or (_23864_, _23862_, _23232_);
  and (_23865_, _23864_, _23514_);
  and (_23867_, _23865_, _23863_);
  nor (_23868_, _23867_, _23859_);
  and (_23869_, _23450_, _23240_);
  and (_23870_, _23480_, _23238_);
  nor (_23871_, _23520_, _23239_);
  not (_23872_, _23232_);
  and (_23873_, _23437_, _23872_);
  or (_23874_, _23873_, _23871_);
  or (_23875_, _23874_, _23870_);
  nor (_23876_, _23875_, _23869_);
  nor (_23877_, _23538_, _23872_);
  not (_23878_, _23877_);
  and (_23879_, _23878_, _23876_);
  nand (_23880_, _23879_, _23868_);
  and (_23881_, _23880_, _22869_);
  nand (_23882_, _23328_, _22986_);
  and (_23883_, _23221_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_23884_, _23883_, _23882_);
  or (_23885_, _23884_, _23881_);
  or (_23886_, _23885_, _23858_);
  and (_23887_, _23886_, _22847_);
  and (_23888_, _23887_, _22983_);
  and (_23889_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  or (_06732_, _23889_, _23888_);
  and (_23890_, \oc8051_top_1.oc8051_sfr1.wait_data , _22731_);
  and (_23891_, _23890_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  and (_23892_, _23783_, _23708_);
  and (_23893_, _23892_, _23792_);
  and (_23894_, _23844_, _23780_);
  or (_23895_, _23894_, _23893_);
  or (_23896_, _23813_, _23824_);
  and (_23897_, _23896_, _23784_);
  and (_23898_, _23797_, _23784_);
  or (_23899_, _23898_, _23897_);
  or (_23900_, _23899_, _23895_);
  or (_23901_, _23846_, _23785_);
  nor (_23902_, _23831_, _23817_);
  and (_23903_, _23799_, _23781_);
  and (_23904_, _23903_, _23780_);
  nand (_23905_, _23904_, _23707_);
  nand (_23906_, _23905_, _23902_);
  or (_23907_, _23906_, _23901_);
  or (_23908_, _23907_, _23900_);
  and (_23909_, _23814_, _23707_);
  and (_23910_, _23909_, _23771_);
  and (_23911_, _23771_, _23707_);
  and (_23912_, _23911_, _23797_);
  or (_23913_, _23912_, _23910_);
  and (_23914_, _23903_, _23814_);
  and (_23915_, _23825_, _23770_);
  and (_23916_, _23915_, _23729_);
  or (_23917_, _23916_, _23914_);
  and (_23918_, _23903_, _23824_);
  and (_23919_, _23903_, _23797_);
  or (_23920_, _23919_, _23918_);
  or (_23921_, _23920_, _23917_);
  or (_23922_, _23921_, _23913_);
  and (_23923_, _23806_, _23779_);
  and (_23924_, _23923_, _23685_);
  and (_23925_, _23818_, _23780_);
  and (_23926_, _23810_, _23781_);
  and (_23927_, _23926_, _23707_);
  and (_23928_, _23927_, _23792_);
  and (_23929_, _23816_, _23783_);
  and (_23930_, _23929_, _23708_);
  nor (_23931_, _23930_, _23928_);
  not (_23932_, _23931_);
  or (_23933_, _23932_, _23925_);
  or (_23934_, _23933_, _23924_);
  or (_23935_, _23934_, _23922_);
  or (_23936_, _23935_, _23908_);
  and (_23937_, _23936_, _23855_);
  or (_26852_[0], _23937_, _23891_);
  and (_23938_, _22922_, _22888_);
  nor (_23939_, _22972_, _22849_);
  and (_23940_, _23939_, _22953_);
  and (_23941_, _23940_, _23938_);
  and (_23943_, _22976_, _22937_);
  and (_23944_, _22968_, _22844_);
  and (_23945_, _23944_, _23943_);
  and (_23946_, _23945_, _23941_);
  and (_23947_, \oc8051_top_1.oc8051_ram_top1.bit_select [2], \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_23948_, _23947_, _23340_);
  nor (_23950_, _23948_, _23504_);
  nor (_23951_, _23538_, _23039_);
  not (_23952_, _23951_);
  not (_23953_, _23514_);
  nor (_23954_, _23566_, _23563_);
  and (_23955_, _23954_, _23150_);
  and (_23957_, _23955_, _23458_);
  nor (_23958_, _23957_, _23364_);
  not (_23959_, _23079_);
  nor (_23960_, _23564_, _23199_);
  and (_23962_, _23960_, _23460_);
  and (_23963_, _23962_, _23115_);
  and (_23964_, _23963_, _23959_);
  nor (_23965_, _23964_, _23456_);
  or (_23966_, _23965_, _23958_);
  nor (_23967_, _23966_, _23487_);
  and (_23968_, _23966_, _23487_);
  nor (_23969_, _23968_, _23967_);
  nor (_23970_, _23969_, _23953_);
  nor (_23971_, _23364_, _23050_);
  not (_23973_, _23971_);
  not (_23974_, _23506_);
  and (_23975_, _23364_, _23039_);
  nor (_23976_, _23975_, _23974_);
  and (_23977_, _23976_, _23973_);
  and (_23978_, _23450_, _23054_);
  and (_23979_, _23480_, _23052_);
  nor (_23980_, _23520_, _23053_);
  and (_23981_, _23437_, _23039_);
  or (_23982_, _23981_, _23980_);
  or (_23983_, _23982_, _23979_);
  nor (_23984_, _23983_, _23978_);
  not (_23985_, _23984_);
  nor (_23986_, _23985_, _23977_);
  not (_23987_, _23986_);
  nor (_23988_, _23987_, _23970_);
  and (_23989_, _23988_, _23952_);
  nor (_23990_, _23989_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_23991_, _23343_, _22869_);
  and (_23992_, _23991_, _23023_);
  or (_23994_, _23992_, _23990_);
  or (_23995_, _23994_, _23950_);
  and (_23996_, _23995_, _22847_);
  and (_23997_, _23996_, _23946_);
  not (_23998_, _23946_);
  and (_23999_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  or (_09147_, _23999_, _23997_);
  nor (_24000_, _22937_, _22871_);
  not (_24001_, _24000_);
  and (_24002_, _24001_, _22847_);
  nor (_24003_, _24002_, _22976_);
  and (_24004_, _22969_, _22844_);
  and (_24005_, _24004_, _22847_);
  and (_24006_, _24005_, _24003_);
  and (_24008_, _24006_, _23941_);
  and (_24009_, _24008_, _23996_);
  not (_24011_, _24008_);
  and (_24013_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or (_13109_, _24013_, _24009_);
  and (_24014_, _22921_, _22890_);
  and (_24015_, _23939_, _22954_);
  and (_24016_, _24015_, _24014_);
  and (_24017_, _24016_, _23945_);
  nand (_24018_, _23947_, _22985_);
  nor (_24019_, _24018_, _23504_);
  and (_24020_, _23364_, _23457_);
  not (_24021_, _24020_);
  nor (_24022_, _23364_, _23122_);
  nor (_24023_, _24022_, _23974_);
  and (_24024_, _24023_, _24021_);
  nor (_24025_, _23962_, _23456_);
  nor (_24026_, _23955_, _23364_);
  nor (_24027_, _24026_, _24025_);
  nor (_24028_, _24027_, _23115_);
  and (_24029_, _24027_, _23115_);
  or (_24030_, _24029_, _23953_);
  nor (_24031_, _24030_, _24028_);
  nor (_24032_, _24031_, _24024_);
  and (_24033_, _23450_, _23125_);
  and (_24034_, _23480_, _23123_);
  nor (_24035_, _23520_, _23124_);
  and (_24036_, _23437_, _23457_);
  or (_24037_, _24036_, _24035_);
  or (_24038_, _24037_, _24034_);
  nor (_24039_, _24038_, _24033_);
  nor (_24040_, _23538_, _23457_);
  not (_24041_, _24040_);
  and (_24042_, _24041_, _24039_);
  and (_24043_, _24042_, _24032_);
  nor (_24044_, _24043_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_24045_, _23336_, _22869_);
  and (_24047_, _24045_, _23104_);
  or (_24048_, _24047_, _24044_);
  or (_24050_, _24048_, _24019_);
  and (_24051_, _24050_, _22847_);
  and (_24052_, _24051_, _24017_);
  not (_24053_, _24017_);
  and (_24054_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  or (_18267_, _24054_, _24052_);
  and (_24055_, _22922_, _22890_);
  and (_24056_, _24055_, _22973_);
  and (_24057_, _24056_, _22982_);
  nand (_24058_, _23947_, _23346_);
  nor (_24059_, _24058_, _23504_);
  nand (_24060_, _23960_, _23364_);
  nand (_24061_, _23954_, _23456_);
  and (_24062_, _24061_, _24060_);
  or (_24063_, _24062_, _23150_);
  nand (_24064_, _24062_, _23150_);
  and (_24065_, _24064_, _24063_);
  nand (_24066_, _24065_, _23514_);
  and (_24067_, _23364_, _23150_);
  nor (_24068_, _23364_, _23156_);
  or (_24069_, _24068_, _23974_);
  nor (_24070_, _24069_, _24067_);
  not (_24071_, _24070_);
  and (_24072_, _24071_, _24066_);
  and (_24073_, _23480_, _23170_);
  and (_24074_, _23437_, _23150_);
  nor (_24075_, _24074_, _24073_);
  nor (_24076_, _23538_, _23150_);
  and (_24077_, _23450_, _23173_);
  nor (_24078_, _23520_, _23172_);
  or (_24079_, _24078_, _24077_);
  nor (_24080_, _24079_, _24076_);
  and (_24081_, _24080_, _24075_);
  and (_24082_, _24081_, _24072_);
  nor (_24083_, _24082_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_24085_, _23349_, _22869_);
  and (_24086_, _24085_, _23140_);
  or (_24087_, _24086_, _24083_);
  or (_24088_, _24087_, _24059_);
  and (_24089_, _24088_, _22847_);
  and (_24091_, _24089_, _24057_);
  not (_24092_, _24057_);
  and (_24093_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  or (_27284_, _24093_, _24091_);
  nor (_24094_, _23939_, _22954_);
  and (_24095_, _24094_, _24055_);
  not (_24096_, _22975_);
  and (_24097_, _24002_, _24096_);
  and (_24098_, _24097_, _22981_);
  and (_24099_, _24098_, _24095_);
  nand (_24100_, _23947_, _23328_);
  nor (_24101_, _24100_, _23504_);
  nor (_24102_, _23364_, _23086_);
  and (_24104_, _23364_, _23959_);
  nor (_24105_, _24104_, _24102_);
  nor (_24106_, _24105_, _23974_);
  or (_24107_, _23963_, _23959_);
  and (_24108_, _24107_, _23965_);
  and (_24109_, _23955_, _23457_);
  nor (_24110_, _24109_, _23079_);
  or (_24111_, _24110_, _23957_);
  and (_24112_, _24111_, _23456_);
  or (_24113_, _24112_, _24108_);
  and (_24114_, _24113_, _23514_);
  nor (_24115_, _24114_, _24106_);
  and (_24116_, _23450_, _23089_);
  and (_24117_, _23480_, _23087_);
  nor (_24118_, _23520_, _23088_);
  and (_24119_, _23437_, _23079_);
  or (_24120_, _24119_, _24118_);
  or (_24121_, _24120_, _24117_);
  nor (_24122_, _24121_, _24116_);
  nor (_24123_, _23538_, _23079_);
  not (_24124_, _24123_);
  and (_24125_, _24124_, _24122_);
  and (_24126_, _24125_, _24115_);
  nor (_24127_, _24126_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_24129_, _23328_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_24130_, _23068_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_24131_, _24130_, _24129_);
  or (_24132_, _24131_, _24127_);
  or (_24133_, _24132_, _24101_);
  and (_24134_, _24133_, _22847_);
  and (_24136_, _24134_, _24099_);
  not (_24137_, _24099_);
  and (_24139_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_27310_, _24139_, _24136_);
  and (_24140_, _24094_, _22923_);
  and (_24141_, _23943_, _22981_);
  and (_24142_, _24141_, _24140_);
  and (_24143_, _24142_, _23548_);
  not (_24144_, _24142_);
  and (_24145_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  or (_22611_, _24145_, _24143_);
  and (_24146_, _24094_, _24014_);
  and (_24147_, _24146_, _24141_);
  and (_24148_, _24147_, _23548_);
  not (_24149_, _24147_);
  and (_24150_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_22616_, _24150_, _24148_);
  and (_24151_, _24142_, _24134_);
  and (_24152_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  or (_22620_, _24152_, _24151_);
  and (_24153_, _24147_, _23887_);
  and (_24154_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_22688_, _24154_, _24153_);
  and (_24155_, _24095_, _22982_);
  and (_24156_, _24155_, _24051_);
  not (_24157_, _24155_);
  and (_24158_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  or (_22689_, _24158_, _24156_);
  and (_24159_, _24055_, _24015_);
  and (_24160_, _24159_, _24098_);
  and (_24161_, _24160_, _23887_);
  not (_24162_, _24160_);
  and (_24163_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  or (_23787_, _24163_, _24161_);
  and (_24164_, _24147_, _23996_);
  and (_24165_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_23949_, _24165_, _24164_);
  and (_24166_, _24147_, _24089_);
  and (_24167_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_23972_, _24167_, _24166_);
  and (_24169_, _23946_, _23548_);
  and (_24170_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  or (_23993_, _24170_, _24169_);
  and (_24171_, _24147_, _24051_);
  and (_24172_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_26923_, _24172_, _24171_);
  and (_24173_, _22936_, _22905_);
  and (_24174_, _24173_, _23944_);
  not (_24175_, _22886_);
  and (_24176_, _22951_, _22919_);
  and (_24177_, _24176_, _24175_);
  nor (_24178_, _22814_, _22811_);
  and (_24179_, _24178_, _22869_);
  not (_24180_, _24179_);
  nor (_24181_, _24180_, _22867_);
  and (_24182_, _24181_, _24177_);
  and (_24184_, _24182_, _24174_);
  or (_24185_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_24186_, _24185_, _22731_);
  and (_24187_, _24177_, _22868_);
  and (_24188_, _24174_, _24179_);
  and (_24189_, _24188_, _24187_);
  nand (_24190_, _24189_, _24126_);
  and (_24427_, _24190_, _24186_);
  nand (_24192_, _23346_, _22987_);
  nor (_24193_, _24192_, _23504_);
  nor (_24194_, _23451_, _23324_);
  nor (_24196_, _24194_, _23449_);
  or (_24197_, _24196_, _23325_);
  and (_24198_, _23480_, _23324_);
  and (_24200_, _23437_, _23296_);
  nor (_24201_, _24200_, _24198_);
  and (_24203_, _23506_, _23301_);
  and (_24204_, _23514_, _23296_);
  nor (_24206_, _24204_, _24203_);
  or (_24207_, _23538_, _23296_);
  and (_24208_, _24207_, _24206_);
  and (_24209_, _24208_, _24201_);
  and (_24210_, _24209_, _24197_);
  nor (_24212_, _24210_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nand (_24214_, _23286_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  nor (_24216_, _24214_, _23347_);
  or (_24217_, _24216_, _24212_);
  or (_24218_, _24217_, _24193_);
  and (_24219_, _24218_, _22847_);
  and (_24220_, _24219_, _23946_);
  and (_24221_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  or (_27056_, _24221_, _24220_);
  and (_24223_, _23938_, _22973_);
  and (_24224_, _24223_, _22982_);
  and (_24225_, _24224_, _23996_);
  not (_24226_, _24224_);
  and (_24228_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_24683_, _24228_, _24225_);
  and (_24229_, _24224_, _24134_);
  and (_24230_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_24796_, _24230_, _24229_);
  and (_24231_, _24224_, _24051_);
  and (_24232_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_24901_, _24232_, _24231_);
  and (_24233_, _24134_, _24008_);
  and (_24234_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_25095_, _24234_, _24233_);
  and (_24236_, _24015_, _22923_);
  and (_24237_, _24236_, _23945_);
  and (_24238_, _24237_, _24089_);
  not (_24239_, _24237_);
  and (_24240_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_25114_, _24240_, _24238_);
  and (_24243_, _23890_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_24244_, _23892_, _23687_);
  or (_24245_, _24244_, _23833_);
  and (_24246_, _23780_, _23771_);
  and (_24247_, _23903_, _23707_);
  and (_24248_, _24247_, _23797_);
  or (_24249_, _24248_, _24246_);
  or (_24250_, _24249_, _24245_);
  and (_24251_, _23927_, _23780_);
  and (_24253_, _23892_, _23780_);
  nor (_24254_, _24253_, _24251_);
  not (_24255_, _24254_);
  and (_24257_, _23811_, _23708_);
  and (_24258_, _24257_, _23687_);
  and (_24259_, _24257_, _23779_);
  nor (_24260_, _24259_, _23928_);
  not (_24261_, _24260_);
  or (_24262_, _24261_, _24258_);
  or (_24263_, _24262_, _24255_);
  or (_24264_, _24263_, _24250_);
  nor (_24265_, _23831_, _23830_);
  nand (_24266_, _23905_, _24265_);
  or (_24267_, _23918_, _23826_);
  and (_24268_, _23909_, _23811_);
  or (_24269_, _23914_, _24268_);
  or (_24270_, _24269_, _24267_);
  or (_24271_, _24270_, _24266_);
  and (_24272_, _23903_, _23708_);
  and (_24273_, _24272_, _23797_);
  and (_24274_, _24257_, _23803_);
  and (_24275_, _23844_, _23797_);
  or (_24276_, _24275_, _24274_);
  or (_24277_, _24276_, _24273_);
  or (_24278_, _22736_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_24279_, _24278_);
  and (_24281_, _23838_, _23804_);
  or (_24283_, _24281_, _24279_);
  or (_24284_, _24283_, _23841_);
  or (_24286_, _24284_, _23846_);
  and (_24287_, _24257_, _23814_);
  or (_24289_, _24287_, _23925_);
  or (_24290_, _24289_, _24286_);
  or (_24291_, _24290_, _24277_);
  or (_24292_, _24291_, _24271_);
  or (_24293_, _24292_, _24264_);
  or (_24294_, _24244_, _24278_);
  and (_24295_, _24294_, _23854_);
  and (_24296_, _24295_, _24293_);
  or (_26851_[0], _24296_, _24243_);
  and (_24297_, _24015_, _23938_);
  nor (_24298_, _22969_, _22844_);
  nor (_24299_, _24298_, _22871_);
  not (_24300_, _24299_);
  and (_24301_, _24300_, _23943_);
  and (_24302_, _24301_, _24297_);
  and (_24303_, _24302_, _23548_);
  not (_24304_, _24302_);
  and (_24305_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  or (_25352_, _24305_, _24303_);
  and (_24306_, _24057_, _23887_);
  and (_24307_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  or (_25419_, _24307_, _24306_);
  and (_24308_, _24057_, _23548_);
  and (_24309_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  or (_25474_, _24309_, _24308_);
  and (_24310_, _23946_, _23583_);
  and (_24311_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  or (_25595_, _24311_, _24310_);
  and (_24312_, _24219_, _24057_);
  and (_24313_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  or (_25624_, _24313_, _24312_);
  and (_24314_, _24237_, _24134_);
  and (_24315_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_27064_, _24315_, _24314_);
  and (_24317_, _23946_, _23887_);
  and (_24318_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  or (_25749_, _24318_, _24317_);
  and (_24319_, _24014_, _22973_);
  and (_24320_, _24319_, _22982_);
  and (_24321_, _24320_, _24134_);
  not (_24322_, _24320_);
  and (_24323_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_25824_, _24323_, _24321_);
  and (_24324_, _24224_, _24219_);
  and (_24325_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_25843_, _24325_, _24324_);
  and (_24327_, _24320_, _23996_);
  and (_24328_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_25943_, _24328_, _24327_);
  and (_24330_, _24223_, _23945_);
  and (_24331_, _24330_, _23548_);
  not (_24332_, _24330_);
  and (_24333_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_26134_, _24333_, _24331_);
  or (_24334_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_24336_, _24334_, _22731_);
  nand (_24337_, _24189_, _24082_);
  and (_26179_, _24337_, _24336_);
  and (_24339_, _24330_, _24219_);
  and (_24340_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_26270_, _24340_, _24339_);
  and (_24341_, _24224_, _23583_);
  and (_24342_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_27282_, _24342_, _24341_);
  and (_24343_, _24224_, _23887_);
  and (_24345_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_27281_, _24345_, _24343_);
  and (_24347_, _24224_, _23548_);
  and (_24348_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_27280_, _24348_, _24347_);
  and (_24349_, _24055_, _23940_);
  and (_24350_, _24349_, _23945_);
  and (_24351_, _24350_, _24051_);
  not (_24352_, _24350_);
  and (_24353_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_27061_, _24353_, _24351_);
  and (_24354_, _24330_, _24089_);
  and (_24355_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_27049_, _24355_, _24354_);
  and (_24357_, _24320_, _24089_);
  and (_24358_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_27278_, _24358_, _24357_);
  and (_24360_, _24330_, _23583_);
  and (_24361_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_27048_, _24361_, _24360_);
  and (_24362_, _24330_, _23887_);
  and (_24364_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_27047_, _24364_, _24362_);
  and (_24365_, _24300_, _24097_);
  and (_24367_, _24365_, _24349_);
  and (_24368_, _24367_, _23996_);
  not (_24369_, _24367_);
  and (_24371_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  or (_27202_, _24371_, _24368_);
  and (_24372_, _24094_, _23938_);
  and (_24373_, _24372_, _22982_);
  and (_24374_, _24373_, _23887_);
  not (_24375_, _24373_);
  and (_24376_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_27270_, _24376_, _24374_);
  and (_24377_, _24373_, _23548_);
  and (_24378_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_27269_, _24378_, _24377_);
  and (_24379_, _24373_, _24219_);
  and (_24380_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_27268_, _24380_, _24379_);
  and (_24381_, _24319_, _23945_);
  and (_24382_, _24381_, _23887_);
  not (_24383_, _24381_);
  and (_24384_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_27043_, _24384_, _24382_);
  and (_24385_, _24381_, _23583_);
  and (_24386_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_27044_, _24386_, _24385_);
  and (_24387_, _24373_, _24051_);
  and (_24388_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_27273_, _24388_, _24387_);
  and (_24389_, _24373_, _24089_);
  and (_24391_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_27272_, _24391_, _24389_);
  and (_24392_, _24373_, _23583_);
  and (_24393_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_27271_, _24393_, _24392_);
  and (_24394_, _24146_, _22982_);
  and (_24395_, _24394_, _24089_);
  not (_24396_, _24394_);
  and (_24397_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_27264_, _24397_, _24395_);
  and (_24398_, _24381_, _24134_);
  and (_24399_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_27046_, _24399_, _24398_);
  and (_24400_, _24394_, _23583_);
  and (_24401_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_27263_, _24401_, _24400_);
  and (_24402_, _24381_, _24051_);
  and (_24403_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_27045_, _24403_, _24402_);
  and (_24404_, _24394_, _23996_);
  and (_24405_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_27267_, _24405_, _24404_);
  and (_24406_, _24394_, _24134_);
  and (_24407_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_27266_, _24407_, _24406_);
  and (_24408_, _24097_, _24004_);
  and (_24409_, _24408_, _24319_);
  and (_24410_, _24409_, _24219_);
  not (_24411_, _24409_);
  and (_24412_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  or (_27118_, _24412_, _24410_);
  and (_24413_, _24394_, _24051_);
  and (_24414_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_27265_, _24414_, _24413_);
  and (_24415_, _23945_, _22974_);
  and (_24416_, _24415_, _24134_);
  not (_24417_, _24415_);
  and (_24418_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  or (_27041_, _24418_, _24416_);
  and (_24420_, _24415_, _24051_);
  and (_24421_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  or (_27040_, _24421_, _24420_);
  or (_24422_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_24424_, _24422_, _22731_);
  nand (_24425_, _24189_, _23989_);
  and (_02924_, _24425_, _24424_);
  and (_24426_, _24155_, _23548_);
  and (_24428_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  or (_27275_, _24428_, _24426_);
  and (_24430_, _24219_, _24155_);
  and (_24431_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  or (_27274_, _24431_, _24430_);
  and (_24433_, _24350_, _23583_);
  and (_24434_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_27059_, _24434_, _24433_);
  and (_03359_, t1_i, _22731_);
  and (_24436_, _24381_, _24219_);
  and (_24437_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_27042_, _24437_, _24436_);
  and (_24438_, _24155_, _23583_);
  and (_24439_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  or (_27277_, _24439_, _24438_);
  and (_24440_, _24155_, _23887_);
  and (_24441_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  or (_27276_, _24441_, _24440_);
  and (_24442_, _24146_, _24006_);
  and (_24443_, _24442_, _23887_);
  not (_24444_, _24442_);
  and (_24446_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  or (_27074_, _24446_, _24443_);
  and (_24447_, _24302_, _23996_);
  and (_24448_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  or (_04393_, _24448_, _24447_);
  and (_24449_, _24415_, _24219_);
  and (_24450_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  or (_27039_, _24450_, _24449_);
  and (_24451_, _24301_, _24146_);
  and (_24452_, _24451_, _24134_);
  not (_24453_, _24451_);
  and (_24454_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_04780_, _24454_, _24452_);
  nor (_24455_, _22737_, _23183_);
  and (_24457_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_24458_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_24459_, _24458_, _24457_);
  and (_24460_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_24461_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_24462_, _24461_, _24460_);
  and (_24464_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_24465_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_24467_, _24465_, _24464_);
  and (_24468_, _24467_, _24462_);
  and (_24469_, _24468_, _24459_);
  and (_24470_, _22737_, _23623_);
  not (_24471_, _24470_);
  nor (_24472_, _24471_, _24469_);
  nor (_24473_, _24472_, _24455_);
  nor (_26867_[3], _24473_, rst);
  and (_24474_, _23940_, _22923_);
  and (_24476_, _24300_, _22977_);
  and (_24478_, _24476_, _24474_);
  and (_24479_, _24478_, _23548_);
  not (_24480_, _24478_);
  and (_24481_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_27171_, _24481_, _24479_);
  and (_24482_, _24478_, _24219_);
  and (_24484_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_04945_, _24484_, _24482_);
  and (_24485_, _24095_, _23945_);
  and (_24486_, _24485_, _23996_);
  not (_24487_, _24485_);
  and (_24489_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  or (_05303_, _24489_, _24486_);
  and (_24490_, _24365_, _24095_);
  and (_24491_, _24490_, _24134_);
  not (_24492_, _24490_);
  and (_24493_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_05608_, _24493_, _24491_);
  and (_24494_, _24409_, _23887_);
  and (_24495_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  or (_05764_, _24495_, _24494_);
  and (_24496_, _24003_, _22981_);
  and (_24497_, _24496_, _24474_);
  and (_24499_, _24497_, _23548_);
  not (_24500_, _24497_);
  and (_24502_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  or (_05861_, _24502_, _24499_);
  and (_24503_, _24365_, _22974_);
  and (_24504_, _24503_, _23548_);
  not (_24505_, _24503_);
  and (_24507_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_05882_, _24507_, _24504_);
  and (_24508_, _24503_, _23887_);
  and (_24509_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_05940_, _24509_, _24508_);
  and (_24510_, _24365_, _24140_);
  and (_24511_, _24510_, _24089_);
  not (_24512_, _24510_);
  and (_24513_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_06025_, _24513_, _24511_);
  and (_24514_, _24415_, _23887_);
  and (_24515_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  or (_06056_, _24515_, _24514_);
  and (_24516_, _24510_, _24051_);
  and (_24517_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_06076_, _24517_, _24516_);
  and (_24518_, _24301_, _24056_);
  and (_24519_, _24518_, _23548_);
  not (_24520_, _24518_);
  and (_24521_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  or (_27219_, _24521_, _24519_);
  and (_24522_, _24510_, _23996_);
  and (_24523_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_06235_, _24523_, _24522_);
  and (_24525_, _24365_, _24146_);
  and (_24526_, _24525_, _24219_);
  not (_24527_, _24525_);
  and (_24528_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  or (_06304_, _24528_, _24526_);
  and (_24529_, _24525_, _23583_);
  and (_24530_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  or (_06382_, _24530_, _24529_);
  not (_24531_, _23504_);
  nor (_24532_, _22919_, _22886_);
  and (_24533_, _24532_, _22951_);
  and (_24534_, _24533_, _24531_);
  nand (_24535_, _22951_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor (_24536_, _24535_, _24532_);
  or (_24537_, _24536_, _24534_);
  and (_24538_, _22968_, _22937_);
  and (_24539_, _24178_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  not (_24540_, _24539_);
  nor (_24541_, _24540_, _22867_);
  and (_24542_, _24541_, _22906_);
  and (_24543_, _24542_, _22844_);
  and (_24544_, _24543_, _24538_);
  and (_24545_, _24544_, _24537_);
  nand (_24546_, _24544_, _22951_);
  and (_24547_, _24546_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor (_24548_, _22936_, _22905_);
  and (_24549_, _24548_, _23944_);
  not (_24550_, _22951_);
  and (_24551_, _24550_, _22867_);
  and (_24552_, _24532_, _24179_);
  and (_24553_, _24552_, _24551_);
  and (_24554_, _24553_, _24549_);
  or (_24555_, _24554_, _24547_);
  or (_24556_, _24555_, _24545_);
  not (_24557_, _24554_);
  or (_24558_, _24557_, _23577_);
  and (_24559_, _24558_, _22731_);
  and (_06442_, _24559_, _24556_);
  not (_24560_, _22919_);
  and (_24561_, _24560_, _22886_);
  and (_24562_, _24561_, _22951_);
  and (_24563_, _24544_, _24562_);
  or (_24564_, _24563_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_24565_, _24564_, _24557_);
  nand (_24566_, _24563_, _23504_);
  and (_24567_, _24566_, _24565_);
  and (_24568_, _24554_, _23880_);
  or (_24569_, _24568_, _24567_);
  and (_06510_, _24569_, _22731_);
  and (_24570_, _24544_, _24177_);
  and (_24571_, _24570_, _23504_);
  nor (_24572_, _24570_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_24573_, _24572_, _24571_);
  nand (_24574_, _24573_, _24557_);
  nand (_24575_, _24554_, _23542_);
  and (_24576_, _24575_, _22731_);
  and (_06536_, _24576_, _24574_);
  and (_24577_, _24176_, _22886_);
  and (_24578_, _24544_, _24577_);
  and (_24579_, _24578_, _23504_);
  nor (_24580_, _24578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_24581_, _24580_, _24579_);
  nand (_24582_, _24581_, _24557_);
  nand (_24583_, _24554_, _24210_);
  and (_24584_, _24583_, _22731_);
  and (_06560_, _24584_, _24582_);
  and (_24585_, _24415_, _23583_);
  and (_24586_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  or (_06601_, _24586_, _24585_);
  and (_24587_, _24525_, _24089_);
  and (_24588_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  or (_06622_, _24588_, _24587_);
  and (_24589_, _24525_, _24134_);
  and (_24590_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  or (_27194_, _24590_, _24589_);
  and (_24591_, _24525_, _23996_);
  and (_24592_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  or (_06722_, _24592_, _24591_);
  nor (_24593_, _22951_, _22919_);
  and (_24594_, _24593_, _22886_);
  and (_24595_, _24594_, _24544_);
  and (_24596_, _24595_, _23504_);
  nor (_24597_, _24595_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_24598_, _24597_, _24596_);
  nand (_24599_, _24598_, _24557_);
  nand (_24600_, _24554_, _24126_);
  and (_24601_, _24600_, _22731_);
  and (_06752_, _24601_, _24599_);
  and (_24602_, _24372_, _24365_);
  and (_24603_, _24602_, _23548_);
  not (_24604_, _24602_);
  and (_24605_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  or (_06772_, _24605_, _24603_);
  and (_24606_, _22919_, _24175_);
  and (_24607_, _24606_, _24550_);
  and (_24608_, _24607_, _24544_);
  nand (_24609_, _24608_, _23504_);
  or (_24610_, _24608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_24611_, _24610_, _24557_);
  and (_24612_, _24611_, _24609_);
  nor (_24613_, _24557_, _24043_);
  or (_24614_, _24613_, _24612_);
  and (_06793_, _24614_, _22731_);
  and (_24615_, _24602_, _23583_);
  and (_24616_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  or (_06814_, _24616_, _24615_);
  and (_24617_, _24602_, _24051_);
  and (_24618_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  or (_06894_, _24618_, _24617_);
  and (_24619_, _24541_, _22905_);
  and (_24620_, _24619_, _22844_);
  and (_24621_, _24620_, _24538_);
  and (_24622_, _24621_, _24177_);
  nand (_24623_, _24622_, _23504_);
  or (_24624_, _24622_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_24625_, _22937_, _22905_);
  and (_24626_, _24625_, _23944_);
  and (_24627_, _24577_, _22868_);
  and (_24628_, _24627_, _24179_);
  and (_24629_, _24628_, _24626_);
  not (_24630_, _24629_);
  and (_24631_, _24630_, _24624_);
  and (_24632_, _24631_, _24623_);
  nor (_24633_, _24630_, _23542_);
  or (_24634_, _24633_, _24632_);
  and (_06967_, _24634_, _22731_);
  and (_24635_, _22919_, _22886_);
  and (_24636_, _24635_, _24550_);
  and (_24637_, _24636_, _24531_);
  nor (_24638_, _24635_, _24550_);
  and (_24639_, _24638_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_24640_, _24639_, _24637_);
  and (_24641_, _24640_, _24621_);
  not (_24642_, _24621_);
  nor (_24643_, _24638_, _24636_);
  or (_24644_, _24643_, _24642_);
  and (_24645_, _24644_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_24646_, _24645_, _24629_);
  or (_24647_, _24646_, _24641_);
  nand (_24648_, _24629_, _24082_);
  and (_24649_, _24648_, _22731_);
  and (_07024_, _24649_, _24647_);
  and (_24650_, _24602_, _24134_);
  and (_24651_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  or (_07047_, _24651_, _24650_);
  and (_24652_, _24621_, _24533_);
  nand (_24653_, _24652_, _23504_);
  or (_24654_, _24652_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_24655_, _24654_, _24630_);
  and (_24656_, _24655_, _24653_);
  and (_24657_, _24629_, _23577_);
  or (_24658_, _24657_, _24656_);
  and (_07072_, _24658_, _22731_);
  and (_24659_, _24621_, _24562_);
  nand (_24660_, _24659_, _23504_);
  or (_24661_, _24659_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_24662_, _24661_, _24630_);
  and (_24663_, _24662_, _24660_);
  and (_24664_, _24629_, _23880_);
  or (_24665_, _24664_, _24663_);
  and (_07135_, _24665_, _22731_);
  and (_24666_, _24621_, _24577_);
  nand (_24667_, _24666_, _23504_);
  or (_24668_, _24666_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_24669_, _24668_, _24630_);
  and (_24670_, _24669_, _24667_);
  not (_24671_, _24210_);
  and (_24672_, _24629_, _24671_);
  or (_24673_, _24672_, _24670_);
  and (_07156_, _24673_, _22731_);
  and (_24674_, _24490_, _24219_);
  and (_24675_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_07199_, _24675_, _24674_);
  and (_24676_, _24490_, _23887_);
  and (_24677_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_07223_, _24677_, _24676_);
  and (_24678_, _24490_, _24089_);
  and (_24679_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_07276_, _24679_, _24678_);
  and (_24680_, _24490_, _24051_);
  and (_24681_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_07366_, _24681_, _24680_);
  and (_24682_, _24503_, _24051_);
  and (_24684_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_07386_, _24684_, _24682_);
  and (_24685_, _24621_, _24594_);
  nand (_24686_, _24685_, _23504_);
  or (_24687_, _24685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_24688_, _24687_, _24630_);
  and (_24689_, _24688_, _24686_);
  nor (_24690_, _24630_, _24126_);
  or (_24691_, _24690_, _24689_);
  and (_07479_, _24691_, _22731_);
  and (_24692_, _24503_, _24134_);
  and (_24693_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_07614_, _24693_, _24692_);
  and (_24694_, _24365_, _24319_);
  and (_24695_, _24694_, _24219_);
  not (_24696_, _24694_);
  and (_24697_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  or (_07645_, _24697_, _24695_);
  and (_24698_, _22968_, _22936_);
  and (_24699_, _24698_, _24620_);
  and (_24700_, _24699_, _24636_);
  nand (_24701_, _24700_, _23504_);
  or (_24702_, _24700_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_24703_, _24628_, _24174_);
  not (_24704_, _24703_);
  and (_24705_, _24704_, _24702_);
  and (_24706_, _24705_, _24701_);
  nor (_24707_, _24704_, _24082_);
  or (_24708_, _24707_, _24706_);
  and (_07703_, _24708_, _22731_);
  and (_24709_, _24699_, _24562_);
  nand (_24710_, _24709_, _23504_);
  or (_24711_, _24709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_24712_, _24711_, _24704_);
  and (_24713_, _24712_, _24710_);
  and (_24714_, _24703_, _23880_);
  or (_24715_, _24714_, _24713_);
  and (_07723_, _24715_, _22731_);
  and (_24716_, _24699_, _24577_);
  or (_24717_, _24716_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_24718_, _24717_, _24704_);
  nand (_24719_, _24716_, _23504_);
  and (_24720_, _24719_, _24718_);
  and (_24721_, _24703_, _24671_);
  or (_24722_, _24721_, _24720_);
  and (_07742_, _24722_, _22731_);
  and (_24723_, _24694_, _23548_);
  and (_24724_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  or (_07762_, _24724_, _24723_);
  and (_24725_, _24694_, _24089_);
  and (_24726_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  or (_07812_, _24726_, _24725_);
  and (_24727_, _24485_, _24219_);
  and (_24728_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  or (_07894_, _24728_, _24727_);
  and (_24729_, _24694_, _24051_);
  and (_24730_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  or (_07923_, _24730_, _24729_);
  and (_24731_, _24694_, _23996_);
  and (_24732_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  or (_07944_, _24732_, _24731_);
  and (_24733_, _24302_, _24134_);
  and (_24734_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  or (_08017_, _24734_, _24733_);
  and (_24735_, _24365_, _24223_);
  and (_24736_, _24735_, _24219_);
  not (_24737_, _24735_);
  and (_24738_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  or (_08087_, _24738_, _24736_);
  and (_24739_, _24485_, _23887_);
  and (_24740_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  or (_08103_, _24740_, _24739_);
  and (_24741_, _24735_, _23583_);
  and (_24742_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  or (_08123_, _24742_, _24741_);
  and (_24743_, _24735_, _24051_);
  and (_24744_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  or (_08142_, _24744_, _24743_);
  and (_24745_, _24735_, _23996_);
  and (_24746_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  or (_08169_, _24746_, _24745_);
  and (_24747_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_24748_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_24749_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_24750_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_24751_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _24750_);
  and (_24752_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_24753_, _24752_, _24751_);
  and (_24754_, _24753_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_24755_, _24754_, _24749_);
  and (_24756_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_24757_, _24756_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_24758_, _24757_);
  and (_24759_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_24760_, _24759_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24761_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_24762_, _24761_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_24763_, _24762_, _24760_);
  and (_24764_, _24763_, _24758_);
  nor (_24765_, _24764_, _24755_);
  not (_24766_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_24767_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_24768_, _24767_, _24766_);
  nand (_24769_, _24768_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_24770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_24771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_24772_, _24771_, _24770_);
  and (_24773_, _24772_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_24774_, _24773_);
  and (_24775_, _24774_, _24769_);
  and (_24776_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_24777_, _24776_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_24778_, _24777_);
  and (_24779_, _24778_, _24775_);
  nor (_24780_, _24779_, _24755_);
  nor (_24781_, _24780_, _24765_);
  and (_24782_, _24749_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not (_24783_, _24782_);
  not (_24784_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_24785_, _24768_, _24784_);
  not (_24786_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_24787_, _24772_, _24786_);
  nor (_24788_, _24787_, _24785_);
  not (_24789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_24790_, _24776_, _24789_);
  not (_24791_, _24790_);
  and (_24792_, _24791_, _24788_);
  nor (_24793_, _24792_, _24783_);
  not (_24794_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_24795_, _24756_, _24794_);
  not (_24797_, _24795_);
  not (_24798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_24799_, _24759_, _24798_);
  not (_24800_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_24801_, _24761_, _24800_);
  nor (_24802_, _24801_, _24799_);
  and (_24803_, _24802_, _24797_);
  nor (_24804_, _24803_, _24783_);
  nor (_24805_, _24804_, _24793_);
  not (_24806_, _24805_);
  and (_24807_, _24806_, _24781_);
  nand (_24808_, _24807_, _24748_);
  not (_24809_, _24781_);
  and (_24810_, _24809_, _24748_);
  or (_24811_, _24810_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and (_24812_, _24811_, _22731_);
  and (_08233_, _24812_, _24808_);
  and (_24813_, _24365_, _24056_);
  and (_24814_, _24813_, _24219_);
  not (_24815_, _24813_);
  and (_24816_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_08294_, _24816_, _24814_);
  and (_24817_, _24485_, _23548_);
  and (_24818_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  or (_08331_, _24818_, _24817_);
  and (_24819_, _24813_, _23887_);
  and (_24820_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_08378_, _24820_, _24819_);
  and (_24821_, _24813_, _24089_);
  and (_24822_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_08397_, _24822_, _24821_);
  and (_26840_[6], _23745_, _22731_);
  and (_24823_, _24813_, _24134_);
  and (_24824_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_08490_, _24824_, _24823_);
  and (_24825_, _24813_, _23996_);
  and (_24826_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_27196_, _24826_, _24825_);
  nor (_24827_, _24747_, _24750_);
  nand (_24828_, _24827_, _24807_);
  and (_24829_, _24827_, _24809_);
  or (_24830_, _24829_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and (_24831_, _24830_, _22731_);
  and (_08572_, _24831_, _24828_);
  and (_24832_, _24474_, _24365_);
  and (_24833_, _24832_, _23887_);
  not (_24834_, _24832_);
  and (_24835_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  or (_08606_, _24835_, _24833_);
  and (_24836_, _24832_, _24089_);
  and (_24837_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  or (_27198_, _24837_, _24836_);
  and (_24838_, _24832_, _24134_);
  and (_24839_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  or (_08724_, _24839_, _24838_);
  and (_24840_, _24805_, _24781_);
  nor (_24841_, _24840_, _24747_);
  not (_24842_, _24841_);
  and (_24843_, _24842_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_24844_, _24747_);
  nor (_24845_, _24769_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_24846_, _24845_, _24777_);
  not (_24847_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_24848_, _24773_, _24750_);
  or (_24849_, _24848_, _24847_);
  nand (_24850_, _24849_, _24846_);
  and (_24851_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_24852_, _24851_, _24778_);
  and (_24853_, _24852_, _24850_);
  or (_24854_, _24853_, _24762_);
  not (_24855_, _24760_);
  not (_24856_, _24762_);
  or (_24857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _24750_);
  or (_24858_, _24857_, _24856_);
  and (_24859_, _24858_, _24855_);
  and (_24860_, _24859_, _24854_);
  and (_24861_, _24851_, _24760_);
  or (_24862_, _24861_, _24757_);
  or (_24863_, _24862_, _24860_);
  nor (_24864_, _24857_, _24758_);
  nor (_24865_, _24864_, _24781_);
  and (_24866_, _24865_, _24863_);
  or (_24867_, _24857_, _24797_);
  and (_24868_, _24785_, _24750_);
  nor (_24869_, _24868_, _24790_);
  and (_24870_, _24787_, _24750_);
  or (_24871_, _24870_, _24847_);
  nand (_24872_, _24871_, _24869_);
  or (_24873_, _24851_, _24791_);
  and (_24874_, _24873_, _24872_);
  or (_24875_, _24874_, _24801_);
  not (_24876_, _24799_);
  not (_24877_, _24801_);
  or (_24878_, _24857_, _24877_);
  and (_24879_, _24878_, _24876_);
  and (_24880_, _24879_, _24875_);
  and (_24881_, _24851_, _24799_);
  or (_24882_, _24881_, _24795_);
  or (_24883_, _24882_, _24880_);
  and (_24884_, _24883_, _24807_);
  and (_24885_, _24884_, _24867_);
  or (_24886_, _24885_, _24866_);
  and (_24887_, _24886_, _24844_);
  or (_24888_, _24887_, _24843_);
  and (_08746_, _24888_, _22731_);
  and (_24889_, _24006_, _22974_);
  and (_24890_, _24889_, _24219_);
  not (_24891_, _24889_);
  and (_24892_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or (_08767_, _24892_, _24890_);
  nand (_24893_, _24840_, _24748_);
  and (_24894_, _24781_, _24844_);
  or (_24895_, _24894_, _24750_);
  and (_24896_, _24895_, _22731_);
  and (_08845_, _24896_, _24893_);
  and (_24897_, _24832_, _23996_);
  and (_24898_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  or (_08971_, _24898_, _24897_);
  and (_24899_, _24014_, _23940_);
  and (_24900_, _24899_, _24365_);
  and (_24902_, _24900_, _23548_);
  not (_24903_, _24900_);
  and (_24904_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_09008_, _24904_, _24902_);
  and (_24905_, _24900_, _23583_);
  and (_24906_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_09032_, _24906_, _24905_);
  and (_24907_, _24900_, _24051_);
  and (_24908_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_09093_, _24908_, _24907_);
  not (_24909_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor (_24910_, _24841_, _24909_);
  or (_24911_, _24778_, _24762_);
  and (_24912_, _24911_, _24855_);
  and (_24913_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _24750_);
  or (_24914_, _24913_, _24912_);
  and (_24915_, _24773_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_24916_, _24915_, _24909_);
  nor (_24917_, _24769_, _24750_);
  nor (_24918_, _24917_, _24777_);
  nand (_24919_, _24918_, _24763_);
  or (_24920_, _24919_, _24916_);
  and (_24921_, _24920_, _24914_);
  or (_24922_, _24921_, _24757_);
  or (_24923_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_24924_, _24856_, _24760_);
  and (_24925_, _24924_, _24758_);
  nor (_24926_, _24925_, _24923_);
  nor (_24927_, _24926_, _24781_);
  and (_24928_, _24927_, _24922_);
  and (_24929_, _24785_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_24930_, _24929_, _24790_);
  and (_24931_, _24787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_24932_, _24931_, _24909_);
  nand (_24933_, _24932_, _24930_);
  or (_24934_, _24913_, _24791_);
  and (_24935_, _24934_, _24933_);
  or (_24936_, _24935_, _24801_);
  or (_24937_, _24923_, _24877_);
  and (_24938_, _24937_, _24876_);
  and (_24939_, _24938_, _24936_);
  and (_24940_, _24913_, _24799_);
  or (_24941_, _24940_, _24795_);
  or (_24942_, _24941_, _24939_);
  and (_24943_, _24807_, _24797_);
  and (_24944_, _24923_, _24807_);
  or (_24945_, _24944_, _24943_);
  and (_24946_, _24945_, _24942_);
  or (_24947_, _24946_, _24928_);
  and (_24948_, _24947_, _24844_);
  or (_24949_, _24948_, _24910_);
  and (_09118_, _24949_, _22731_);
  and (_24950_, _24900_, _24134_);
  and (_24951_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_27200_, _24951_, _24950_);
  and (_24952_, _24365_, _23941_);
  and (_24953_, _24952_, _23548_);
  not (_24954_, _24952_);
  and (_24955_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_27201_, _24955_, _24953_);
  and (_24956_, _24952_, _23887_);
  and (_24957_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_09448_, _24957_, _24956_);
  and (_24959_, _24952_, _24089_);
  and (_24960_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_09479_, _24960_, _24959_);
  and (_24961_, _24952_, _24134_);
  and (_24962_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_09499_, _24962_, _24961_);
  and (_24963_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_24964_, _24963_, _24841_);
  and (_09539_, _24964_, _22731_);
  or (_24965_, _24801_, _24790_);
  nor (_24966_, _24799_, _24795_);
  nand (_24967_, _24966_, _24782_);
  or (_24968_, _24967_, _24965_);
  nor (_24969_, _24968_, _24788_);
  and (_24970_, _24969_, _24781_);
  and (_24971_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor (_24972_, _24777_, _24755_);
  not (_24973_, _24764_);
  nor (_24974_, _24775_, _24973_);
  and (_24975_, _24974_, _24972_);
  and (_24976_, _24975_, _24844_);
  or (_24977_, _24976_, _24971_);
  or (_24978_, _24977_, _24970_);
  and (_09560_, _24978_, _22731_);
  and (_24979_, _24788_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_24980_, _24979_, _24965_);
  and (_24981_, _24980_, _24966_);
  and (_24982_, _24981_, _24807_);
  nor (_24983_, _24760_, _24757_);
  or (_24984_, _24777_, _24762_);
  and (_24985_, _24775_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_24986_, _24985_, _24984_);
  nand (_24987_, _24986_, _24983_);
  nor (_24988_, _24987_, _24781_);
  or (_24989_, _24988_, _24747_);
  or (_24990_, _24989_, _24982_);
  or (_24991_, _24844_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_24992_, _24991_, _22731_);
  and (_09580_, _24992_, _24990_);
  and (_24993_, _24367_, _24219_);
  and (_24994_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  or (_09600_, _24994_, _24993_);
  nor (_24995_, _24787_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_24996_, _24995_, _24785_);
  or (_24997_, _24996_, _24790_);
  and (_24998_, _24997_, _24877_);
  or (_24999_, _24998_, _24799_);
  and (_25000_, _24999_, _24943_);
  or (_25001_, _24773_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_25002_, _25001_, _24769_);
  or (_25003_, _25002_, _24777_);
  and (_25004_, _25003_, _24856_);
  or (_25005_, _25004_, _24760_);
  nor (_25006_, _24781_, _24757_);
  and (_25007_, _25006_, _25005_);
  or (_25008_, _25007_, _24747_);
  or (_25009_, _25008_, _25000_);
  not (_25010_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nand (_25011_, _24747_, _25010_);
  and (_25012_, _25011_, _22731_);
  and (_09621_, _25012_, _25009_);
  and (_25013_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _22731_);
  and (_09650_, _25013_, _24747_);
  and (_25014_, _24367_, _23548_);
  and (_25015_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  or (_09745_, _25015_, _25014_);
  and (_25016_, _22906_, _22867_);
  and (_25017_, _25016_, _22844_);
  and (_25018_, _25017_, _24538_);
  and (_25019_, _25018_, _24533_);
  nand (_25020_, _25019_, _23504_);
  or (_25021_, _25019_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_25022_, _25021_, _24539_);
  and (_25023_, _25022_, _25020_);
  and (_25024_, _24577_, _22867_);
  and (_25025_, _25024_, _24548_);
  and (_25026_, _25025_, _23944_);
  not (_25027_, _25026_);
  or (_25028_, _25027_, _23577_);
  or (_25029_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_25030_, _25029_, _24179_);
  and (_25032_, _25030_, _25028_);
  not (_25033_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_25034_, _24178_, _25033_);
  or (_25035_, _25034_, rst);
  or (_25036_, _25035_, _25032_);
  or (_09786_, _25036_, _25023_);
  and (_25038_, _24367_, _23583_);
  and (_25039_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  or (_09809_, _25039_, _25038_);
  and (_25040_, _25018_, _24562_);
  nand (_25041_, _25040_, _23504_);
  or (_25042_, _25040_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_25043_, _25042_, _24539_);
  and (_25044_, _25043_, _25041_);
  or (_25045_, _25027_, _23880_);
  or (_25046_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_25047_, _25046_, _24179_);
  and (_25048_, _25047_, _25045_);
  not (_25049_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_25050_, _24178_, _25049_);
  or (_25051_, _25050_, rst);
  or (_25052_, _25051_, _25048_);
  or (_09868_, _25052_, _25044_);
  and (_25053_, _25018_, _24177_);
  nand (_25054_, _25053_, _23504_);
  or (_25055_, _25053_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_25056_, _25055_, _24539_);
  and (_25057_, _25056_, _25054_);
  nand (_25058_, _25026_, _23542_);
  or (_25059_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_25060_, _25059_, _24179_);
  and (_25061_, _25060_, _25058_);
  not (_25062_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_25063_, _24178_, _25062_);
  or (_25064_, _25063_, rst);
  or (_25065_, _25064_, _25061_);
  or (_09894_, _25065_, _25057_);
  and (_25066_, _25018_, _24577_);
  nand (_25067_, _25066_, _23504_);
  or (_25068_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_25069_, _25068_, _24539_);
  and (_25070_, _25069_, _25067_);
  nand (_25071_, _25026_, _24210_);
  and (_25072_, _25071_, _24179_);
  and (_25073_, _25072_, _25068_);
  not (_25074_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_25075_, _24178_, _25074_);
  or (_25077_, _25075_, rst);
  or (_25078_, _25077_, _25073_);
  or (_09922_, _25078_, _25070_);
  and (_25080_, _24367_, _24051_);
  and (_25081_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  or (_09986_, _25081_, _25080_);
  and (_25083_, _24485_, _24051_);
  and (_25084_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  or (_10012_, _25084_, _25083_);
  and (_25085_, _24485_, _24089_);
  and (_25086_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  or (_10107_, _25086_, _25085_);
  and (_25088_, _25018_, _24594_);
  nand (_25089_, _25088_, _23504_);
  or (_25090_, _25088_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_25091_, _25090_, _24539_);
  and (_25092_, _25091_, _25089_);
  nand (_25093_, _25026_, _24126_);
  or (_25094_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_25096_, _25094_, _24179_);
  and (_25097_, _25096_, _25093_);
  not (_25098_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_25099_, _24178_, _25098_);
  or (_25100_, _25099_, rst);
  or (_25101_, _25100_, _25097_);
  or (_10136_, _25101_, _25092_);
  and (_25102_, _24478_, _23583_);
  and (_25103_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_10250_, _25103_, _25102_);
  and (_25104_, _25018_, _24607_);
  nand (_25105_, _25104_, _23504_);
  or (_25106_, _25104_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_25107_, _25106_, _24539_);
  and (_25108_, _25107_, _25105_);
  nand (_25109_, _25026_, _24043_);
  or (_25110_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_25111_, _25110_, _24179_);
  and (_25112_, _25111_, _25109_);
  not (_25113_, _24178_);
  and (_25115_, _25113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_25116_, _25115_, rst);
  or (_25117_, _25116_, _25112_);
  or (_10293_, _25117_, _25108_);
  and (_25118_, _24485_, _23583_);
  and (_25119_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  or (_10347_, _25119_, _25118_);
  and (_25120_, _24478_, _23887_);
  and (_25121_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_10382_, _25121_, _25120_);
  and (_25122_, _22905_, _22867_);
  and (_25123_, _25122_, _22844_);
  and (_25124_, _25123_, _24538_);
  and (_25125_, _25124_, _24177_);
  nand (_25126_, _25125_, _23504_);
  or (_25127_, _25125_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_25128_, _25127_, _24539_);
  and (_25129_, _25128_, _25126_);
  and (_25130_, _25024_, _24626_);
  nand (_25131_, _25130_, _23542_);
  or (_25132_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_25133_, _25132_, _24179_);
  and (_25134_, _25133_, _25131_);
  not (_25135_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_25136_, _24178_, _25135_);
  or (_25137_, _25136_, rst);
  or (_25138_, _25137_, _25134_);
  or (_10460_, _25138_, _25129_);
  and (_25139_, _25124_, _24607_);
  nand (_25140_, _25139_, _23504_);
  or (_25141_, _25139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_25142_, _25141_, _24539_);
  and (_25143_, _25142_, _25140_);
  nand (_25144_, _25130_, _24043_);
  or (_25145_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_25146_, _25145_, _24179_);
  and (_25147_, _25146_, _25144_);
  and (_25148_, _25113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_25149_, _25148_, rst);
  or (_25150_, _25149_, _25147_);
  or (_10482_, _25150_, _25143_);
  and (_25151_, _25124_, _24636_);
  nand (_25152_, _25151_, _23504_);
  or (_25153_, _25151_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_25154_, _25153_, _24539_);
  and (_25155_, _25154_, _25152_);
  nand (_25156_, _25130_, _24082_);
  or (_25157_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_25158_, _25157_, _24179_);
  and (_25159_, _25158_, _25156_);
  not (_25160_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor (_25161_, _24178_, _25160_);
  or (_25162_, _25161_, rst);
  or (_25163_, _25162_, _25159_);
  or (_10516_, _25163_, _25155_);
  and (_25164_, _25124_, _24533_);
  nand (_25165_, _25164_, _23504_);
  or (_25166_, _25164_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_25167_, _25166_, _24539_);
  and (_25168_, _25167_, _25165_);
  not (_25169_, _25130_);
  or (_25171_, _25169_, _23577_);
  or (_25172_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_25173_, _25172_, _24179_);
  and (_25174_, _25173_, _25171_);
  not (_25175_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor (_25176_, _24178_, _25175_);
  or (_25177_, _25176_, rst);
  or (_25178_, _25177_, _25174_);
  or (_10541_, _25178_, _25168_);
  and (_25179_, _25124_, _24562_);
  nand (_25180_, _25179_, _23504_);
  or (_25181_, _25179_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_25182_, _25181_, _24539_);
  and (_25183_, _25182_, _25180_);
  or (_25184_, _25169_, _23880_);
  or (_25185_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_25186_, _25185_, _24179_);
  and (_25187_, _25186_, _25184_);
  not (_25188_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_25189_, _24178_, _25188_);
  or (_25190_, _25189_, rst);
  or (_25191_, _25190_, _25187_);
  or (_10565_, _25191_, _25183_);
  and (_25192_, _25124_, _24577_);
  nand (_25193_, _25192_, _23504_);
  or (_25194_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_25195_, _25194_, _24539_);
  and (_25196_, _25195_, _25193_);
  nand (_25197_, _25130_, _24210_);
  and (_25198_, _25197_, _24179_);
  and (_25199_, _25198_, _25194_);
  not (_25200_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_25201_, _24178_, _25200_);
  or (_25202_, _25201_, rst);
  or (_25203_, _25202_, _25199_);
  or (_10592_, _25203_, _25196_);
  and (_25204_, _24237_, _23996_);
  and (_25205_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_27065_, _25205_, _25204_);
  and (_25206_, _24372_, _23945_);
  and (_25207_, _25206_, _24089_);
  not (_25208_, _25206_);
  and (_25209_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_10727_, _25209_, _25207_);
  and (_25210_, _24476_, _24056_);
  and (_25211_, _25210_, _23583_);
  not (_25212_, _25210_);
  and (_25213_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  or (_10764_, _25213_, _25211_);
  and (_25214_, _25210_, _23887_);
  and (_25215_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  or (_10780_, _25215_, _25214_);
  and (_25216_, _25210_, _23548_);
  and (_25217_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  or (_10796_, _25217_, _25216_);
  and (_25218_, _25206_, _24051_);
  and (_25219_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_10814_, _25219_, _25218_);
  and (_25220_, _25017_, _24698_);
  and (_25221_, _25220_, _24533_);
  nand (_25222_, _25221_, _23504_);
  or (_25223_, _25221_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_25224_, _25223_, _24539_);
  and (_25225_, _25224_, _25222_);
  and (_25226_, _22936_, _22906_);
  and (_25227_, _25226_, _23944_);
  and (_25228_, _25227_, _25024_);
  not (_25229_, _25228_);
  or (_25230_, _25229_, _23577_);
  or (_25231_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_25232_, _25231_, _24179_);
  and (_25233_, _25232_, _25230_);
  not (_25234_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_25235_, _24178_, _25234_);
  or (_25236_, _25235_, rst);
  or (_25238_, _25236_, _25233_);
  or (_10934_, _25238_, _25225_);
  and (_25240_, _25220_, _24562_);
  nand (_25241_, _25240_, _23504_);
  or (_25242_, _25240_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_25243_, _25242_, _24539_);
  and (_25244_, _25243_, _25241_);
  or (_25246_, _25229_, _23880_);
  or (_25247_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_25248_, _25247_, _24179_);
  and (_25249_, _25248_, _25246_);
  not (_25250_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_25251_, _24178_, _25250_);
  or (_25252_, _25251_, rst);
  or (_25253_, _25252_, _25249_);
  or (_10960_, _25253_, _25244_);
  and (_25254_, _25220_, _24177_);
  nand (_25255_, _25254_, _23504_);
  or (_25256_, _25254_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_25257_, _25256_, _24539_);
  and (_25258_, _25257_, _25255_);
  nand (_25259_, _25228_, _23542_);
  or (_25260_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_25261_, _25260_, _24179_);
  and (_25262_, _25261_, _25259_);
  not (_25263_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_25264_, _24178_, _25263_);
  or (_25266_, _25264_, rst);
  or (_25267_, _25266_, _25262_);
  or (_10987_, _25267_, _25258_);
  and (_25268_, _25220_, _24577_);
  nand (_25269_, _25268_, _23504_);
  or (_25270_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_25271_, _25270_, _24539_);
  and (_25272_, _25271_, _25269_);
  nand (_25274_, _25228_, _24210_);
  and (_25275_, _25274_, _24179_);
  and (_25276_, _25275_, _25270_);
  not (_25277_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_25278_, _24178_, _25277_);
  or (_25279_, _25278_, rst);
  or (_25280_, _25279_, _25276_);
  or (_11035_, _25280_, _25272_);
  and (_25281_, _25210_, _24134_);
  and (_25283_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  or (_27155_, _25283_, _25281_);
  and (_25284_, _25210_, _24051_);
  and (_25285_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  or (_11161_, _25285_, _25284_);
  and (_25286_, _25220_, _24594_);
  nand (_25287_, _25286_, _23504_);
  or (_25288_, _25286_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_25289_, _25288_, _24539_);
  and (_25290_, _25289_, _25287_);
  nand (_25291_, _25228_, _24126_);
  or (_25292_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_25293_, _25292_, _24179_);
  and (_25294_, _25293_, _25291_);
  not (_25295_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_25296_, _24178_, _25295_);
  or (_25297_, _25296_, rst);
  or (_25298_, _25297_, _25294_);
  or (_11255_, _25298_, _25290_);
  and (_25299_, _25220_, _24607_);
  nand (_25300_, _25299_, _23504_);
  or (_25301_, _25299_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_25302_, _25301_, _24539_);
  and (_25303_, _25302_, _25300_);
  nand (_25305_, _25228_, _24043_);
  or (_25306_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_25307_, _25306_, _24179_);
  and (_25308_, _25307_, _25305_);
  and (_25309_, _25113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_25310_, _25309_, rst);
  or (_25311_, _25310_, _25308_);
  or (_11356_, _25311_, _25303_);
  and (_25312_, _25206_, _24134_);
  and (_25313_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_11416_, _25313_, _25312_);
  and (_25314_, _24476_, _24223_);
  and (_25315_, _25314_, _24051_);
  not (_25316_, _25314_);
  and (_25318_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_11589_, _25318_, _25315_);
  and (_25319_, _25123_, _24698_);
  and (_25320_, _25319_, _24562_);
  nand (_25321_, _25320_, _23504_);
  or (_25322_, _25320_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_25323_, _25322_, _24539_);
  and (_25325_, _25323_, _25321_);
  and (_25327_, _25319_, _24577_);
  not (_25328_, _25327_);
  or (_25329_, _25328_, _23880_);
  or (_25330_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_25331_, _25330_, _24179_);
  and (_25332_, _25331_, _25329_);
  not (_25333_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_25334_, _24178_, _25333_);
  or (_25335_, _25334_, rst);
  or (_25336_, _25335_, _25332_);
  or (_11618_, _25336_, _25325_);
  and (_25338_, _25319_, _24177_);
  nand (_25339_, _25338_, _23504_);
  or (_25340_, _25338_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_25341_, _25340_, _24539_);
  and (_25342_, _25341_, _25339_);
  nand (_25343_, _25327_, _23542_);
  or (_25344_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_25345_, _25344_, _24179_);
  and (_25346_, _25345_, _25343_);
  not (_25347_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_25349_, _24178_, _25347_);
  or (_25350_, _25349_, rst);
  or (_25351_, _25350_, _25346_);
  or (_11644_, _25351_, _25342_);
  nand (_25353_, _25327_, _23504_);
  or (_25354_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_25355_, _25354_, _24539_);
  and (_25356_, _25355_, _25353_);
  nand (_25357_, _25327_, _24210_);
  and (_25358_, _25357_, _24179_);
  and (_25359_, _25358_, _25354_);
  not (_25360_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_25361_, _24178_, _25360_);
  or (_25362_, _25361_, rst);
  or (_25363_, _25362_, _25359_);
  or (_11669_, _25363_, _25356_);
  and (_25364_, _25314_, _24089_);
  and (_25365_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_27122_, _25365_, _25364_);
  and (_25366_, _25319_, _24607_);
  nand (_25367_, _25366_, _23504_);
  or (_25368_, _25366_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_25369_, _25368_, _24539_);
  and (_25370_, _25369_, _25367_);
  nand (_25371_, _25327_, _24043_);
  or (_25372_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_25374_, _25372_, _24179_);
  and (_25375_, _25374_, _25371_);
  and (_25376_, _25113_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_25377_, _25376_, rst);
  or (_25378_, _25377_, _25375_);
  or (_11891_, _25378_, _25370_);
  and (_25380_, _25206_, _24219_);
  and (_25381_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_27036_, _25381_, _25380_);
  and (_25382_, _25319_, _24594_);
  nand (_25383_, _25382_, _23504_);
  or (_25384_, _25382_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_25385_, _25384_, _24539_);
  and (_25386_, _25385_, _25383_);
  nand (_25387_, _25327_, _24126_);
  or (_25388_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_25390_, _25388_, _24179_);
  and (_25391_, _25390_, _25387_);
  not (_25392_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_25393_, _24178_, _25392_);
  or (_25394_, _25393_, rst);
  or (_25395_, _25394_, _25391_);
  or (_11973_, _25395_, _25386_);
  not (_25396_, _25319_);
  or (_25397_, _25396_, _24643_);
  and (_25398_, _25397_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_25400_, _24638_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_25401_, _25400_, _24637_);
  and (_25402_, _25401_, _25319_);
  or (_25403_, _25402_, _25398_);
  and (_25404_, _25403_, _24539_);
  nand (_25405_, _25327_, _24082_);
  or (_25406_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_25407_, _25406_, _24179_);
  and (_25408_, _25407_, _25405_);
  not (_25409_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_25410_, _24178_, _25409_);
  or (_25411_, _25410_, rst);
  or (_25412_, _25411_, _25408_);
  or (_11994_, _25412_, _25404_);
  and (_25413_, _24004_, _23943_);
  and (_25414_, _25413_, _24146_);
  and (_25415_, _25414_, _23548_);
  not (_25416_, _25414_);
  and (_25417_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or (_12065_, _25417_, _25415_);
  and (_25418_, _25314_, _23996_);
  and (_25420_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_12243_, _25420_, _25418_);
  and (_25421_, _25314_, _24134_);
  and (_25422_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_12266_, _25422_, _25421_);
  and (_25423_, _25206_, _23887_);
  and (_25424_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_12515_, _25424_, _25423_);
  and (_25425_, _25206_, _23548_);
  and (_25426_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_12616_, _25426_, _25425_);
  and (_25428_, _25314_, _24219_);
  and (_25429_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_12637_, _25429_, _25428_);
  and (_25430_, _24302_, _24051_);
  and (_25431_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  or (_27231_, _25431_, _25430_);
  and (_25432_, _24476_, _24319_);
  and (_25433_, _25432_, _23996_);
  not (_25434_, _25432_);
  and (_25435_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_27100_, _25435_, _25433_);
  and (_25436_, _25432_, _24134_);
  and (_25438_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_12748_, _25438_, _25436_);
  and (_25440_, _24302_, _24089_);
  and (_25441_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  or (_14268_, _25441_, _25440_);
  and (_25442_, _24146_, _23945_);
  and (_25443_, _25442_, _24089_);
  not (_25444_, _25442_);
  and (_25445_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_15162_, _25445_, _25443_);
  and (_25446_, _25314_, _23887_);
  and (_25447_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_15213_, _25447_, _25446_);
  and (_25448_, _25442_, _23583_);
  and (_25449_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_15234_, _25449_, _25448_);
  and (_25450_, _25314_, _23548_);
  and (_25451_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_15619_, _25451_, _25450_);
  nor (_25453_, _22737_, _23011_);
  not (_25454_, _22737_);
  and (_25455_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_25456_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  not (_25457_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_25458_, _23601_, _25457_);
  nor (_25459_, _25458_, _25456_);
  and (_25460_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_25461_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_25462_, _25461_, _25460_);
  and (_25463_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_25465_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_25466_, _25465_, _25463_);
  and (_25467_, _25466_, _25462_);
  and (_25469_, _25467_, _25459_);
  nor (_25470_, _25469_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_25472_, _25470_, _25455_);
  nor (_25473_, _25472_, _25454_);
  nor (_25475_, _25473_, _25453_);
  nor (_26877_[7], _25475_, rst);
  nor (_26840_[3], _23615_, rst);
  or (_25477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor (_25478_, _22968_, _22937_);
  and (_25479_, _25478_, _24620_);
  or (_25480_, _25479_, _25477_);
  and (_25481_, _24532_, _24550_);
  and (_25482_, _25481_, _24531_);
  not (_25483_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_25484_, _25481_, _25483_);
  nand (_25485_, _25484_, _25479_);
  or (_25486_, _25485_, _25482_);
  and (_25487_, _25486_, _25480_);
  and (_25488_, _24173_, _24004_);
  and (_25489_, _25488_, _24628_);
  or (_25490_, _25489_, _25487_);
  nand (_25491_, _25489_, _23989_);
  and (_25492_, _25491_, _22731_);
  and (_17618_, _25492_, _25490_);
  and (_25493_, _25442_, _24134_);
  and (_25494_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_27034_, _25494_, _25493_);
  and (_25495_, _25432_, _24219_);
  and (_25496_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_27099_, _25496_, _25495_);
  and (_25497_, _24636_, _24181_);
  and (_25499_, _25497_, _25488_);
  and (_25500_, _24607_, _24181_);
  and (_25501_, _25500_, _25488_);
  nor (_25502_, _25501_, _25499_);
  or (_25503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_25504_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_25505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _25504_);
  and (_25506_, _25505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_25507_, _25506_, _25503_);
  and (_25508_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_25509_, _25508_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_25510_, _25509_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_25511_, _25510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_25512_, _25511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_25513_, _25512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_25514_, _25513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_25515_, _25514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_25516_, _25515_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_25517_, _25516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_25518_, _25517_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_25519_, _25518_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_25520_, _25519_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_25521_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_25522_, _25521_, _25520_);
  and (_25523_, _25522_, _25507_);
  nor (_25524_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  not (_25526_, _25524_);
  not (_25527_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_25528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_25529_, _25528_, _25524_);
  and (_25531_, _25529_, _25527_);
  nor (_25532_, _25531_, _25526_);
  nand (_25533_, _25532_, _25523_);
  nand (_25534_, _25533_, _25502_);
  or (_25535_, _25502_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_25536_, _25535_, _22731_);
  and (_17752_, _25536_, _25534_);
  and (_25538_, _25524_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not (_25539_, _25538_);
  or (_25540_, _25529_, _25523_);
  and (_25541_, _25540_, _25539_);
  and (_25542_, _25541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_25543_, _25520_, _25507_);
  and (_25544_, _25543_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_25545_, _25544_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor (_25546_, _25531_, _25523_);
  or (_25547_, _25546_, _25499_);
  and (_25548_, _25547_, _25545_);
  or (_25549_, _25548_, _25542_);
  not (_25550_, _25499_);
  nor (_25551_, _25550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor (_25552_, _25551_, _25501_);
  and (_25553_, _25552_, _25549_);
  not (_25554_, _23989_);
  and (_25556_, _24607_, _22868_);
  and (_25557_, _25556_, _24179_);
  and (_25558_, _25557_, _25488_);
  and (_25560_, _25558_, _25554_);
  or (_25561_, _25560_, _25553_);
  and (_17768_, _25561_, _22731_);
  nor (_25563_, _22737_, _23133_);
  and (_25564_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_25565_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_25566_, _25565_, _25564_);
  and (_25567_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_25568_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_25569_, _25568_, _25567_);
  and (_25571_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_25572_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_25573_, _25572_, _25571_);
  and (_25574_, _25573_, _25569_);
  and (_25575_, _25574_, _25566_);
  nor (_25576_, _25575_, _24471_);
  nor (_25577_, _25576_, _25563_);
  nor (_26867_[4], _25577_, rst);
  nor (_25578_, _25550_, _23989_);
  not (_25579_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor (_25580_, _25538_, _25579_);
  and (_25581_, _25580_, _25523_);
  and (_25582_, _25513_, _25507_);
  or (_25583_, _25582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_25584_, _25582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_25585_, _25584_, _25583_);
  or (_25586_, _25585_, _25531_);
  or (_25587_, _25586_, _25581_);
  nand (_25588_, _25531_, _25579_);
  and (_25589_, _25588_, _25502_);
  and (_25590_, _25589_, _25587_);
  and (_25591_, _25558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_25592_, _25591_, _25590_);
  or (_25593_, _25592_, _25578_);
  and (_17818_, _25593_, _22731_);
  and (_25594_, _25526_, _25507_);
  and (_25596_, _25594_, _25502_);
  or (_25597_, _25596_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_25598_, _25522_);
  nand (_25599_, _25596_, _25598_);
  and (_25600_, _25599_, _22731_);
  and (_17853_, _25600_, _25597_);
  and (_25601_, _24533_, _22868_);
  and (_25602_, _25601_, _24179_);
  and (_25603_, _25602_, _25488_);
  nand (_25604_, _25603_, _23989_);
  and (_25605_, _25538_, _25528_);
  not (_25606_, _25605_);
  and (_25607_, _24562_, _24181_);
  and (_25608_, _25607_, _25488_);
  nor (_25609_, _25608_, _25606_);
  not (_25610_, _25609_);
  and (_25611_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_25612_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_25613_, _25612_, _25611_);
  or (_25614_, _25603_, _25613_);
  and (_25615_, _25614_, _22731_);
  and (_17922_, _25615_, _25604_);
  nand (_25616_, _25608_, _23989_);
  not (_25617_, _25603_);
  nor (_25618_, _25605_, _25579_);
  and (_25619_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_25620_, _25619_, _25618_);
  or (_25621_, _25620_, _25608_);
  and (_25622_, _25621_, _25617_);
  and (_25623_, _25622_, _25616_);
  and (_25625_, _25603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_25626_, _25625_, _25623_);
  and (_17942_, _25626_, _22731_);
  and (_17956_, t2ex_i, _22731_);
  and (_25627_, _24476_, _22974_);
  and (_25628_, _25627_, _23996_);
  not (_25629_, _25627_);
  and (_25630_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  or (_17998_, _25630_, _25628_);
  and (_25631_, _24350_, _24089_);
  and (_25632_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_27060_, _25632_, _25631_);
  nand (_25633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _22731_);
  nor (_18105_, _25633_, t2ex_i);
  nor (_25634_, t2_i, rst);
  and (_18119_, _25634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  and (_18134_, t2_i, _22731_);
  and (_25635_, _24350_, _23996_);
  and (_25636_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_18155_, _25636_, _25635_);
  and (_25637_, _24301_, _24223_);
  and (_25639_, _25637_, _24219_);
  not (_25640_, _25637_);
  and (_25642_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_18176_, _25642_, _25639_);
  and (_25643_, _25432_, _23887_);
  and (_25644_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_18441_, _25644_, _25643_);
  and (_25645_, _25432_, _23583_);
  and (_25647_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_18950_, _25647_, _25645_);
  and (_25648_, _24140_, _23945_);
  and (_25649_, _25648_, _23996_);
  not (_25650_, _25648_);
  and (_25651_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  or (_19201_, _25651_, _25649_);
  and (_25652_, _25627_, _24219_);
  and (_25654_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  or (_19605_, _25654_, _25652_);
  and (_25656_, _25627_, _23887_);
  and (_25657_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  or (_19639_, _25657_, _25656_);
  and (_25658_, _24496_, _24056_);
  and (_25659_, _25658_, _24134_);
  not (_25660_, _25658_);
  and (_25661_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or (_19907_, _25661_, _25659_);
  and (_25662_, _25627_, _23548_);
  and (_25663_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  or (_27090_, _25663_, _25662_);
  and (_25664_, _25442_, _24219_);
  and (_25665_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_27033_, _25665_, _25664_);
  and (_25666_, _25627_, _24051_);
  and (_25668_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  or (_21388_, _25668_, _25666_);
  and (_25669_, _25627_, _24089_);
  and (_25670_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  or (_21519_, _25670_, _25669_);
  and (_25672_, _24365_, _24016_);
  and (_25673_, _25672_, _24051_);
  not (_25674_, _25672_);
  and (_25675_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_21620_, _25675_, _25673_);
  and (_25677_, _25627_, _23583_);
  and (_25679_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  or (_21642_, _25679_, _25677_);
  and (_26865_[0], _23685_, _22731_);
  and (_26865_[1], _23664_, _22731_);
  and (_26865_[2], _23643_, _22731_);
  and (_25681_, _25024_, _24179_);
  and (_25682_, _25226_, _24004_);
  and (_25683_, _25682_, _25681_);
  not (_25684_, _25683_);
  and (_25685_, _25684_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_25686_, _25683_, _23577_);
  or (_25687_, _25686_, _25685_);
  and (_26865_[3], _25687_, _22731_);
  and (_25689_, _25648_, _24089_);
  and (_25691_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  or (_27031_, _25691_, _25689_);
  nor (_25692_, _23592_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_25693_, _25692_, _25454_);
  nor (_25694_, _25693_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_25695_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  not (_25696_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nand (_25697_, _25694_, _25696_);
  and (_25698_, _25697_, _22731_);
  and (_26883_[0], _25698_, _25695_);
  or (_25699_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  not (_25700_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand (_25701_, _25694_, _25700_);
  and (_25703_, _25701_, _22731_);
  and (_26883_[1], _25703_, _25699_);
  or (_25704_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  not (_25705_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand (_25707_, _25694_, _25705_);
  and (_25709_, _25707_, _22731_);
  and (_26883_[2], _25709_, _25704_);
  or (_25710_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  not (_25711_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nand (_25712_, _25694_, _25711_);
  and (_25713_, _25712_, _22731_);
  and (_26883_[3], _25713_, _25710_);
  or (_25714_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  not (_25715_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand (_25716_, _25694_, _25715_);
  and (_25718_, _25716_, _22731_);
  and (_26883_[4], _25718_, _25714_);
  or (_25719_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  not (_25720_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand (_25721_, _25694_, _25720_);
  and (_25722_, _25721_, _22731_);
  and (_26883_[5], _25722_, _25719_);
  or (_25723_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  not (_25724_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand (_25726_, _25694_, _25724_);
  and (_25727_, _25726_, _22731_);
  and (_26883_[6], _25727_, _25723_);
  or (_25728_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  not (_25729_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nand (_25730_, _25694_, _25729_);
  and (_25732_, _25730_, _22731_);
  and (_26883_[7], _25732_, _25728_);
  or (_25734_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not (_25735_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_25736_, _25694_, _25735_);
  and (_25737_, _25736_, _22731_);
  and (_26883_[8], _25737_, _25734_);
  or (_25738_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  not (_25739_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_25740_, _25694_, _25739_);
  and (_25741_, _25740_, _22731_);
  and (_26883_[9], _25741_, _25738_);
  or (_25743_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  not (_25744_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand (_25745_, _25694_, _25744_);
  and (_25746_, _25745_, _22731_);
  and (_26883_[10], _25746_, _25743_);
  or (_25748_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  not (_25750_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_25751_, _25694_, _25750_);
  and (_25752_, _25751_, _22731_);
  and (_26883_[11], _25752_, _25748_);
  or (_25753_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  not (_25754_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nand (_25755_, _25694_, _25754_);
  and (_25756_, _25755_, _22731_);
  and (_26883_[12], _25756_, _25753_);
  or (_25757_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  not (_25758_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_25759_, _25694_, _25758_);
  and (_25760_, _25759_, _22731_);
  and (_26883_[13], _25760_, _25757_);
  or (_25761_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  not (_25763_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_25764_, _25694_, _25763_);
  and (_25765_, _25764_, _22731_);
  and (_26883_[14], _25765_, _25761_);
  or (_25766_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  not (_25767_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_25768_, _25694_, _25767_);
  and (_25769_, _25768_, _22731_);
  and (_26883_[15], _25769_, _25766_);
  or (_25770_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  not (_25771_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand (_25772_, _25694_, _25771_);
  and (_25773_, _25772_, _22731_);
  and (_26883_[16], _25773_, _25770_);
  or (_25775_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  not (_25776_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand (_25777_, _25694_, _25776_);
  and (_25778_, _25777_, _22731_);
  and (_26883_[17], _25778_, _25775_);
  or (_25779_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  not (_25780_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand (_25781_, _25694_, _25780_);
  and (_25782_, _25781_, _22731_);
  and (_26883_[18], _25782_, _25779_);
  or (_25783_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  not (_25784_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand (_25785_, _25694_, _25784_);
  and (_25786_, _25785_, _22731_);
  and (_26883_[19], _25786_, _25783_);
  or (_25787_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  not (_25788_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand (_25789_, _25694_, _25788_);
  and (_25790_, _25789_, _22731_);
  and (_26883_[20], _25790_, _25787_);
  or (_25791_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  not (_25792_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand (_25793_, _25694_, _25792_);
  and (_25794_, _25793_, _22731_);
  and (_26883_[21], _25794_, _25791_);
  or (_25795_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  not (_25796_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand (_25797_, _25694_, _25796_);
  and (_25798_, _25797_, _22731_);
  and (_26883_[22], _25798_, _25795_);
  or (_25799_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  not (_25800_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand (_25801_, _25694_, _25800_);
  and (_25802_, _25801_, _22731_);
  and (_26883_[23], _25802_, _25799_);
  or (_25803_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  not (_25804_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand (_25805_, _25694_, _25804_);
  and (_25806_, _25805_, _22731_);
  and (_26883_[24], _25806_, _25803_);
  or (_25807_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  not (_25808_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_25809_, _25694_, _25808_);
  and (_25810_, _25809_, _22731_);
  and (_26883_[25], _25810_, _25807_);
  or (_25811_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  not (_25812_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_25813_, _25694_, _25812_);
  and (_25814_, _25813_, _22731_);
  and (_26883_[26], _25814_, _25811_);
  or (_25815_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  not (_25816_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand (_25817_, _25694_, _25816_);
  and (_25818_, _25817_, _22731_);
  and (_26883_[27], _25818_, _25815_);
  or (_25819_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  not (_25820_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand (_25821_, _25694_, _25820_);
  and (_25822_, _25821_, _22731_);
  and (_26883_[28], _25822_, _25819_);
  or (_25823_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  not (_25825_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_25826_, _25694_, _25825_);
  and (_25827_, _25826_, _22731_);
  and (_26883_[29], _25827_, _25823_);
  or (_25828_, _25694_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  not (_25829_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand (_25830_, _25694_, _25829_);
  and (_25831_, _25830_, _22731_);
  and (_26883_[30], _25831_, _25828_);
  and (_25832_, _25684_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_25833_, _25684_, _24082_);
  nor (_25834_, _25833_, _25832_);
  nor (_25835_, _25834_, _22906_);
  and (_25836_, _25834_, _22906_);
  nor (_25837_, _25836_, _25835_);
  or (_25838_, _25687_, _22867_);
  nor (_25839_, _25686_, _25685_);
  or (_25840_, _25839_, _22868_);
  and (_25841_, _23685_, _22886_);
  nor (_25842_, _23685_, _22886_);
  nor (_25844_, _25842_, _25841_);
  and (_25845_, _24176_, _22978_);
  and (_25846_, _25845_, _24298_);
  and (_25848_, _25846_, _25844_);
  and (_25849_, _25848_, _22936_);
  and (_25850_, _25849_, _25840_);
  and (_25851_, _25850_, _25838_);
  and (_25852_, _25851_, _25837_);
  and (_25854_, _25852_, _24210_);
  not (_25855_, _25834_);
  and (_25856_, _25687_, _23685_);
  and (_25858_, _25856_, _25855_);
  nand (_25859_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_25860_, _25839_, _23791_);
  and (_25861_, _25860_, _25834_);
  nand (_25862_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_25863_, _25862_, _25859_);
  and (_25864_, _25687_, _23791_);
  and (_25865_, _25864_, _25855_);
  nand (_25866_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_25867_, _25856_, _25834_);
  nand (_25868_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_25869_, _25868_, _25866_);
  and (_25870_, _25869_, _25863_);
  not (_25872_, _25852_);
  and (_25873_, _25839_, _23685_);
  and (_25874_, _25873_, _25855_);
  nand (_25876_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_25877_, _25873_, _25834_);
  nand (_25878_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_25879_, _25878_, _25876_);
  and (_25880_, _25860_, _25855_);
  nand (_25881_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_25882_, _25864_, _25834_);
  nand (_25884_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_25885_, _25884_, _25881_);
  and (_25886_, _25885_, _25879_);
  and (_25888_, _25886_, _25872_);
  and (_25890_, _25888_, _25870_);
  nor (_25891_, _25890_, _25854_);
  and (_26866_[0], _25891_, _22731_);
  and (_25892_, _25852_, _23542_);
  and (_25893_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_25894_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_25895_, _25894_, _25893_);
  and (_25896_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_25897_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor (_25898_, _25897_, _25896_);
  and (_25899_, _25898_, _25895_);
  and (_25900_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_25901_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_25902_, _25901_, _25900_);
  and (_25903_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_25905_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_25907_, _25905_, _25903_);
  and (_25908_, _25907_, _25902_);
  and (_25909_, _25908_, _25872_);
  and (_25910_, _25909_, _25899_);
  nor (_25911_, _25910_, _25892_);
  and (_26866_[1], _25911_, _22731_);
  nor (_25912_, _25872_, _23880_);
  and (_25913_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_25914_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_25915_, _25914_, _25913_);
  and (_25916_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_25917_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_25918_, _25917_, _25916_);
  and (_25919_, _25918_, _25915_);
  and (_25920_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_25921_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_25922_, _25921_, _25920_);
  and (_25923_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_25924_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_25925_, _25924_, _25923_);
  and (_25926_, _25925_, _25922_);
  and (_25928_, _25926_, _25872_);
  and (_25929_, _25928_, _25919_);
  nor (_25930_, _25929_, _25912_);
  and (_26866_[2], _25930_, _22731_);
  and (_25931_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_25932_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_25933_, _25932_, _25931_);
  and (_25934_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_25935_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_25936_, _25935_, _25934_);
  and (_25937_, _25936_, _25933_);
  nand (_25938_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nand (_25940_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_25941_, _25940_, _25938_);
  nand (_25942_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nand (_25944_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_25945_, _25944_, _25942_);
  and (_25947_, _25945_, _25941_);
  and (_25948_, _25947_, _25872_);
  and (_25950_, _25948_, _25937_);
  not (_25951_, _23577_);
  and (_25952_, _25852_, _25951_);
  nor (_25954_, _25952_, _25950_);
  and (_26866_[3], _25954_, _22731_);
  and (_25955_, _25852_, _24082_);
  and (_25956_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  and (_25958_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_25959_, _25958_, _25956_);
  and (_25961_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_25962_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_25963_, _25962_, _25961_);
  and (_25964_, _25963_, _25959_);
  and (_25965_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_25967_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor (_25968_, _25967_, _25965_);
  and (_25969_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_25970_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_25971_, _25970_, _25969_);
  and (_25973_, _25971_, _25968_);
  and (_25974_, _25973_, _25872_);
  and (_25975_, _25974_, _25964_);
  nor (_25976_, _25975_, _25955_);
  and (_26866_[4], _25976_, _22731_);
  and (_25977_, _25852_, _24043_);
  and (_25978_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_25979_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_25980_, _25979_, _25978_);
  and (_25981_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_25982_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_25983_, _25982_, _25981_);
  and (_25984_, _25983_, _25980_);
  and (_25985_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_25986_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_25987_, _25986_, _25985_);
  and (_25988_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_25989_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_25990_, _25989_, _25988_);
  and (_25991_, _25990_, _25987_);
  and (_25992_, _25991_, _25872_);
  and (_25994_, _25992_, _25984_);
  nor (_25995_, _25994_, _25977_);
  and (_26866_[5], _25995_, _22731_);
  and (_25997_, _25852_, _24126_);
  and (_25998_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_25999_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_26000_, _25999_, _25998_);
  and (_26001_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_26002_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor (_26003_, _26002_, _26001_);
  and (_26005_, _26003_, _26000_);
  and (_26006_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_26007_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_26008_, _26007_, _26006_);
  and (_26010_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_26011_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_26013_, _26011_, _26010_);
  and (_26014_, _26013_, _26008_);
  and (_26016_, _26014_, _25872_);
  and (_26017_, _26016_, _26005_);
  nor (_26018_, _26017_, _25997_);
  and (_26866_[6], _26018_, _22731_);
  and (_26020_, _24476_, _24095_);
  and (_26021_, _26020_, _23583_);
  not (_26022_, _26020_);
  and (_26023_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  or (_22612_, _26023_, _26021_);
  and (_26024_, _26020_, _23887_);
  and (_26025_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  or (_22613_, _26025_, _26024_);
  and (_26027_, _25648_, _23583_);
  and (_26028_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  or (_27030_, _26028_, _26027_);
  and (_26031_, _24051_, _22983_);
  and (_26032_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  or (_22614_, _26032_, _26031_);
  and (_26034_, _26020_, _23548_);
  and (_26035_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  or (_22615_, _26035_, _26034_);
  nor (_26036_, _22737_, _23097_);
  and (_26037_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_26038_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_26039_, _26038_, _26037_);
  and (_26040_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_26041_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_26042_, _26041_, _26040_);
  and (_26043_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_26044_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_26045_, _26044_, _26043_);
  and (_26047_, _26045_, _26042_);
  and (_26048_, _26047_, _26039_);
  nor (_26049_, _26048_, _24471_);
  nor (_26050_, _26049_, _26036_);
  nor (_26867_[5], _26050_, rst);
  nor (_26051_, _22737_, _23248_);
  and (_26053_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_26054_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_26055_, _26054_, _26053_);
  and (_26057_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_26058_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_26059_, _26058_, _26057_);
  and (_26060_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_26061_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_26063_, _26061_, _26060_);
  and (_26064_, _26063_, _26059_);
  and (_26066_, _26064_, _26055_);
  nor (_26067_, _26066_, _24471_);
  nor (_26068_, _26067_, _26051_);
  nor (_26867_[1], _26068_, rst);
  and (_26840_[4], _23703_, _22731_);
  nor (_26070_, _22737_, _23095_);
  and (_26071_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_26072_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_26073_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_26074_, _26073_, _26072_);
  and (_26076_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_26077_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_26079_, _26077_, _26076_);
  and (_26080_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_26081_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_26082_, _26081_, _26080_);
  and (_26083_, _26082_, _26079_);
  and (_26084_, _26083_, _26074_);
  nor (_26085_, _26084_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_26087_, _26085_, _26071_);
  nor (_26088_, _26087_, _25454_);
  nor (_26089_, _26088_, _26070_);
  nor (_26877_[5], _26089_, rst);
  nor (_26090_, _22737_, _23060_);
  and (_26091_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_26092_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_26093_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_26094_, _26093_, _26092_);
  and (_26095_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_26097_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_26098_, _26097_, _26095_);
  and (_26099_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_26100_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_26101_, _26100_, _26099_);
  and (_26102_, _26101_, _26098_);
  and (_26103_, _26102_, _26094_);
  nor (_26104_, _26103_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_26106_, _26104_, _26091_);
  nor (_26107_, _26106_, _25454_);
  nor (_26108_, _26107_, _26090_);
  nor (_26877_[6], _26108_, rst);
  and (_26110_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_26111_, _22740_, _22806_);
  or (_26112_, _26111_, _26110_);
  and (_26862_[14], _26112_, _22731_);
  and (_26113_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_26114_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_26115_, _22740_, _26114_);
  or (_26116_, _26115_, _26113_);
  and (_26862_[13], _26116_, _22731_);
  and (_26118_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_26119_, _22740_, _22797_);
  or (_26120_, _26119_, _26118_);
  and (_26862_[12], _26120_, _22731_);
  and (_26121_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_26122_, _22740_, _22793_);
  or (_26123_, _26122_, _26121_);
  and (_26862_[11], _26123_, _22731_);
  and (_26124_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_26125_, _22740_, _22789_);
  or (_26126_, _26125_, _26124_);
  and (_26862_[10], _26126_, _22731_);
  and (_26127_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not (_26128_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_26129_, _22740_, _26128_);
  or (_26130_, _26129_, _26127_);
  and (_26862_[9], _26130_, _22731_);
  and (_26131_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_26132_, _22740_, _22780_);
  or (_26133_, _26132_, _26131_);
  and (_26862_[8], _26133_, _22731_);
  and (_26135_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_26136_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_26137_, _22740_, _26136_);
  or (_26138_, _26137_, _26135_);
  and (_26862_[7], _26138_, _22731_);
  and (_26139_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_26140_, _22740_, _22772_);
  or (_26141_, _26140_, _26139_);
  and (_26862_[6], _26141_, _22731_);
  and (_26142_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_26143_, _22740_, _22767_);
  or (_26144_, _26143_, _26142_);
  and (_26862_[5], _26144_, _22731_);
  and (_26145_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_26146_, _22740_, _22762_);
  or (_26147_, _26146_, _26145_);
  and (_26862_[4], _26147_, _22731_);
  and (_26148_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_26149_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_26150_, _22740_, _26149_);
  or (_26151_, _26150_, _26148_);
  and (_26862_[3], _26151_, _22731_);
  and (_26152_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_26153_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_26154_, _22740_, _26153_);
  or (_26155_, _26154_, _26152_);
  and (_26862_[2], _26155_, _22731_);
  nor (_26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_26157_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and (_26158_, _26156_, _23296_);
  nor (_26159_, _26158_, _26157_);
  not (_26160_, _26159_);
  and (_26161_, _23301_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_26162_, _26161_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26163_, _23086_, _23049_);
  nor (_26164_, _26163_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_26165_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_26166_, _23237_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_26167_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26168_, _23156_, _26167_);
  nand (_26169_, _26168_, _26166_);
  or (_26170_, _23156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26171_, _23084_, _26167_);
  nand (_26172_, _26171_, _26170_);
  and (_26173_, _26172_, _26169_);
  or (_26174_, _23371_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26175_, _23122_, _26167_);
  nand (_26176_, _26175_, _26174_);
  or (_26177_, _23122_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_26178_, _23049_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_26180_, _26178_, _26177_);
  and (_26181_, _26180_, _26176_);
  nand (_26182_, _26181_, _26173_);
  and (_26183_, _26182_, _26165_);
  nor (_26184_, _26183_, _26164_);
  or (_26185_, _23269_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26186_, _23371_, _26167_);
  nand (_26187_, _26186_, _26185_);
  and (_26188_, _26187_, _26165_);
  and (_26189_, _26180_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_26190_, _26189_, _26188_);
  not (_26191_, _26190_);
  nand (_26192_, _26156_, _23039_);
  nor (_26193_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_26194_, _26193_);
  and (_26195_, _26194_, _26192_);
  not (_26196_, _26195_);
  or (_26197_, _23301_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26198_, _23237_, _26167_);
  and (_26199_, _26198_, _26197_);
  or (_26200_, _26199_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26201_, _26172_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26202_, _26201_, _26200_);
  or (_26203_, _26202_, _26196_);
  and (_26204_, _23269_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_26205_, _26204_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26206_, _26176_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_26207_, _26206_, _26205_);
  nand (_26208_, _26156_, _23079_);
  nor (_26209_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_26210_, _26209_);
  and (_26211_, _26210_, _26208_);
  not (_26212_, _26211_);
  or (_26213_, _26212_, _26207_);
  nand (_26214_, _26201_, _26200_);
  or (_26215_, _26214_, _26195_);
  and (_26216_, _26215_, _26203_);
  not (_26217_, _26216_);
  or (_26218_, _26217_, _26213_);
  and (_26219_, _26218_, _26203_);
  nand (_26220_, _26206_, _26205_);
  or (_26221_, _26211_, _26220_);
  and (_26222_, _26221_, _26213_);
  and (_26223_, _26222_, _26216_);
  not (_26224_, _26156_);
  or (_26225_, _26224_, _23115_);
  nor (_26226_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_26227_, _26226_);
  and (_26228_, _26227_, _26225_);
  or (_26229_, _26161_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26230_, _26169_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_26231_, _26230_, _26229_);
  nand (_26232_, _26231_, _26228_);
  or (_26233_, _26231_, _26228_);
  nand (_26234_, _26233_, _26232_);
  nor (_26235_, _26187_, _26165_);
  nand (_26236_, _26156_, _23150_);
  nor (_26237_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_26238_, _26237_);
  and (_26239_, _26238_, _26236_);
  not (_26240_, _26239_);
  or (_26241_, _26240_, _26235_);
  or (_26242_, _26241_, _26234_);
  nand (_26243_, _26242_, _26232_);
  nand (_26244_, _26243_, _26223_);
  and (_26245_, _26244_, _26219_);
  and (_26246_, _26199_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_26247_, _26246_);
  nor (_26248_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_26249_, _26248_);
  nand (_26250_, _26156_, _23199_);
  and (_26251_, _26250_, _26249_);
  nand (_26252_, _26251_, _26247_);
  or (_26253_, _26251_, _26247_);
  nand (_26254_, _26253_, _26252_);
  nand (_26255_, _26204_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_26256_, _26224_, _23232_);
  nor (_26257_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_26258_, _26257_);
  and (_26259_, _26258_, _26256_);
  nand (_26260_, _26259_, _26255_);
  or (_26261_, _26224_, _23264_);
  nor (_26262_, _26156_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_26263_, _26262_);
  nand (_26264_, _26263_, _26261_);
  and (_26265_, _26264_, _26162_);
  or (_26266_, _26259_, _26255_);
  nand (_26267_, _26266_, _26260_);
  or (_26268_, _26267_, _26265_);
  and (_26269_, _26268_, _26260_);
  or (_26271_, _26269_, _26254_);
  nand (_26272_, _26271_, _26252_);
  and (_26273_, _26233_, _26232_);
  not (_26274_, _26235_);
  or (_26275_, _26239_, _26274_);
  and (_26276_, _26275_, _26241_);
  and (_26277_, _26276_, _26273_);
  and (_26278_, _26277_, _26223_);
  nand (_26279_, _26278_, _26272_);
  nand (_26280_, _26279_, _26245_);
  and (_26281_, _26191_, _26184_);
  nand (_26282_, _26281_, _26280_);
  and (_26283_, _26282_, _26195_);
  not (_26284_, _26283_);
  and (_26285_, _26281_, _26280_);
  and (_26286_, _26276_, _26272_);
  not (_26287_, _26286_);
  and (_26288_, _26287_, _26241_);
  or (_26289_, _26288_, _26234_);
  and (_26290_, _26289_, _26232_);
  not (_26291_, _26290_);
  nand (_26292_, _26291_, _26222_);
  and (_26293_, _26292_, _26213_);
  nand (_26294_, _26293_, _26216_);
  or (_26295_, _26293_, _26216_);
  nand (_26296_, _26295_, _26294_);
  nand (_26297_, _26296_, _26285_);
  nand (_26298_, _26297_, _26284_);
  or (_26299_, _26298_, _26191_);
  nand (_26300_, _26298_, _26191_);
  or (_26301_, _26291_, _26222_);
  nand (_26302_, _26301_, _26292_);
  nand (_26303_, _26302_, _26285_);
  and (_26304_, _26282_, _26212_);
  not (_26305_, _26304_);
  and (_26306_, _26305_, _26303_);
  and (_26307_, _26306_, _26214_);
  not (_26308_, _26307_);
  nand (_26309_, _26308_, _26300_);
  nand (_26310_, _26309_, _26299_);
  and (_26311_, _26300_, _26299_);
  nor (_26312_, _26306_, _26214_);
  nor (_26313_, _26312_, _26307_);
  and (_26314_, _26313_, _26311_);
  nand (_26315_, _26288_, _26234_);
  nand (_26316_, _26315_, _26289_);
  nand (_26317_, _26316_, _26285_);
  nor (_26318_, _26285_, _26228_);
  not (_26319_, _26318_);
  and (_26320_, _26319_, _26317_);
  and (_26321_, _26320_, _26220_);
  nor (_26322_, _26276_, _26272_);
  nor (_26323_, _26322_, _26286_);
  nor (_26324_, _26323_, _26282_);
  and (_26325_, _26282_, _26240_);
  nor (_26326_, _26325_, _26324_);
  and (_26327_, _26326_, _26231_);
  not (_26328_, _26327_);
  nor (_26329_, _26320_, _26220_);
  or (_26330_, _26321_, _26329_);
  nor (_26331_, _26330_, _26328_);
  or (_26332_, _26331_, _26321_);
  and (_26333_, _26269_, _26254_);
  not (_26334_, _26333_);
  and (_26335_, _26334_, _26271_);
  or (_26336_, _26335_, _26282_);
  or (_26337_, _26285_, _26251_);
  and (_26338_, _26337_, _26336_);
  nor (_26339_, _26338_, _26274_);
  not (_26340_, _26339_);
  not (_26341_, _26162_);
  or (_26342_, _26282_, _26341_);
  nand (_26343_, _26342_, _26264_);
  or (_26344_, _26342_, _26264_);
  and (_26345_, _26344_, _26343_);
  nand (_26346_, _26345_, _26255_);
  or (_26347_, _26345_, _26255_);
  and (_26348_, _26347_, _26346_);
  nor (_26349_, _26341_, _26159_);
  not (_26350_, _26349_);
  nand (_26351_, _26350_, _26348_);
  and (_26352_, _26351_, _26346_);
  and (_26353_, _26267_, _26265_);
  not (_26354_, _26353_);
  and (_26355_, _26354_, _26268_);
  or (_26356_, _26355_, _26282_);
  or (_26357_, _26285_, _26259_);
  and (_26358_, _26357_, _26356_);
  nand (_26359_, _26358_, _26247_);
  or (_26360_, _26358_, _26247_);
  and (_26361_, _26360_, _26359_);
  not (_26362_, _26361_);
  or (_26363_, _26362_, _26352_);
  and (_26364_, _26338_, _26274_);
  not (_26365_, _26364_);
  and (_26366_, _26365_, _26359_);
  nand (_26367_, _26366_, _26363_);
  and (_26368_, _26367_, _26340_);
  nor (_26369_, _26326_, _26231_);
  nor (_26370_, _26369_, _26327_);
  not (_26371_, _26330_);
  and (_26372_, _26371_, _26370_);
  and (_26373_, _26372_, _26368_);
  or (_26374_, _26373_, _26332_);
  nand (_26375_, _26374_, _26314_);
  nand (_26376_, _26375_, _26310_);
  and (_26377_, _26376_, _26184_);
  and (_26378_, _26377_, _26162_);
  nor (_26379_, _26378_, _26160_);
  and (_26380_, _26378_, _26160_);
  or (_26381_, _26380_, _26379_);
  nand (_26382_, _26381_, _23528_);
  and (_26383_, _23364_, _23403_);
  nor (_26384_, _26383_, _23404_);
  nand (_26385_, _23390_, _26384_);
  and (_26386_, _23477_, _23487_);
  nor (_26387_, _23484_, _23461_);
  nor (_26388_, _26387_, _23296_);
  nor (_26389_, _26388_, _26386_);
  and (_26390_, _26389_, _24197_);
  and (_26391_, _26390_, _24201_);
  and (_26392_, _26391_, _26385_);
  nor (_26393_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_26394_, _26393_);
  and (_26395_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  nand (_26396_, _26393_, _23049_);
  not (_26397_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_26398_, _26397_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_26399_, _26398_);
  or (_26400_, _26399_, _23120_);
  not (_26401_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_26402_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _26401_);
  not (_26403_, _26402_);
  or (_26404_, _26403_, _23205_);
  and (_26405_, _26404_, _26400_);
  nor (_26406_, _26402_, _26398_);
  or (_26407_, _23269_, _26401_);
  nand (_26408_, _26407_, _26406_);
  nand (_26409_, _26408_, _26405_);
  and (_26410_, _26409_, _26396_);
  and (_26411_, _26410_, _23264_);
  or (_26412_, _26394_, _23084_);
  or (_26413_, _26399_, _23169_);
  or (_26414_, _26403_, _23310_);
  and (_26415_, _26414_, _26413_);
  or (_26416_, _23301_, _26401_);
  nand (_26417_, _26416_, _26406_);
  nand (_26418_, _26417_, _26415_);
  and (_26419_, _26418_, _26412_);
  and (_26420_, _26419_, _23232_);
  nand (_26421_, _26420_, _26411_);
  and (_26422_, _26419_, _23563_);
  nand (_26423_, _26418_, _26412_);
  or (_26424_, _26423_, _23509_);
  and (_26425_, _26410_, _23232_);
  and (_26426_, _26425_, _26424_);
  nand (_26427_, _26426_, _26422_);
  nand (_26428_, _26427_, _26421_);
  nand (_26429_, _26409_, _26396_);
  or (_26430_, _26429_, _23199_);
  or (_26431_, _26423_, _23150_);
  or (_26432_, _26431_, _26430_);
  nand (_26433_, _26431_, _26430_);
  and (_26434_, _26433_, _26432_);
  and (_26435_, _26434_, _26428_);
  and (_26436_, _26410_, _23460_);
  and (_26437_, _26436_, _26422_);
  or (_26438_, _26429_, _23457_);
  or (_26439_, _26438_, _26431_);
  and (_26440_, _26419_, _23115_);
  or (_26441_, _26440_, _26436_);
  and (_26442_, _26441_, _26439_);
  nand (_26443_, _26442_, _26437_);
  or (_26444_, _26442_, _26437_);
  and (_26445_, _26444_, _26443_);
  nand (_26446_, _26445_, _26435_);
  not (_26447_, _26438_);
  or (_26448_, _26439_, _23079_);
  and (_26449_, _26419_, _23959_);
  not (_26450_, _26449_);
  nand (_26451_, _26450_, _26439_);
  and (_26452_, _26451_, _26448_);
  nand (_26453_, _26452_, _26447_);
  or (_26454_, _26449_, _26447_);
  nand (_26455_, _26454_, _26453_);
  or (_26456_, _26455_, _26446_);
  and (_26457_, _26419_, _23491_);
  and (_26458_, _26457_, _26411_);
  or (_26459_, _26420_, _26411_);
  and (_26460_, _26459_, _26421_);
  and (_26461_, _26460_, _26458_);
  or (_26462_, _26426_, _26422_);
  and (_26463_, _26462_, _26427_);
  nand (_26464_, _26463_, _26461_);
  not (_26465_, _26464_);
  nand (_26466_, _26434_, _26428_);
  or (_26467_, _26434_, _26428_);
  and (_26468_, _26467_, _26466_);
  nand (_26469_, _26468_, _26465_);
  or (_26470_, _26445_, _26435_);
  nand (_26471_, _26470_, _26446_);
  or (_26472_, _26471_, _26469_);
  and (_26473_, _26446_, _26443_);
  nand (_26474_, _26473_, _26455_);
  or (_26475_, _26473_, _26455_);
  nand (_26476_, _26475_, _26474_);
  or (_26477_, _26476_, _26472_);
  and (_26478_, _26477_, _26456_);
  nor (_26479_, _26455_, _26443_);
  not (_26480_, _26448_);
  and (_26481_, _26452_, _26447_);
  or (_26482_, _26423_, _23039_);
  or (_26483_, _26429_, _23079_);
  or (_26484_, _26483_, _26482_);
  nand (_26485_, _26483_, _26482_);
  and (_26486_, _26485_, _26484_);
  nand (_26487_, _26486_, _26481_);
  or (_26488_, _26486_, _26481_);
  and (_26489_, _26488_, _26487_);
  nand (_26490_, _26489_, _26480_);
  or (_26491_, _26489_, _26480_);
  and (_26492_, _26491_, _26490_);
  nand (_26493_, _26492_, _26479_);
  or (_26494_, _26492_, _26479_);
  nand (_26495_, _26494_, _26493_);
  or (_26496_, _26495_, _26478_);
  nand (_26497_, _26495_, _26478_);
  and (_26498_, _26497_, _26496_);
  nand (_26499_, _26498_, _26395_);
  or (_26500_, _26498_, _26395_);
  and (_26501_, _26500_, _26499_);
  and (_26502_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nand (_26503_, _26476_, _26472_);
  and (_26504_, _26503_, _26477_);
  nand (_26505_, _26504_, _26502_);
  or (_26506_, _26504_, _26502_);
  nand (_26507_, _26506_, _26505_);
  and (_26508_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nand (_26509_, _26471_, _26469_);
  and (_26510_, _26509_, _26472_);
  nand (_26511_, _26510_, _26508_);
  or (_26512_, _26510_, _26508_);
  nand (_26513_, _26512_, _26511_);
  and (_26514_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or (_26515_, _26468_, _26465_);
  and (_26516_, _26515_, _26469_);
  nand (_26517_, _26516_, _26514_);
  and (_26518_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or (_26519_, _26463_, _26461_);
  and (_26520_, _26519_, _26464_);
  nand (_26521_, _26520_, _26518_);
  and (_26522_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand (_26523_, _26460_, _26458_);
  or (_26524_, _26460_, _26458_);
  and (_26525_, _26524_, _26523_);
  and (_26526_, _26525_, _26522_);
  not (_26527_, _26526_);
  or (_26528_, _26520_, _26518_);
  nand (_26529_, _26528_, _26521_);
  or (_26530_, _26529_, _26527_);
  and (_26531_, _26530_, _26521_);
  or (_26532_, _26516_, _26514_);
  nand (_26533_, _26532_, _26517_);
  or (_26534_, _26533_, _26531_);
  and (_26535_, _26534_, _26517_);
  or (_26536_, _26535_, _26513_);
  and (_26537_, _26536_, _26511_);
  or (_26538_, _26537_, _26507_);
  nand (_26539_, _26538_, _26505_);
  nand (_26540_, _26539_, _26501_);
  nand (_26541_, _26540_, _26499_);
  and (_26542_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  nand (_26543_, _26496_, _26493_);
  and (_26544_, _26410_, _23487_);
  and (_26545_, _26544_, _26450_);
  and (_26546_, _26490_, _26487_);
  not (_26547_, _26546_);
  nand (_26548_, _26547_, _26545_);
  or (_26549_, _26547_, _26545_);
  and (_26550_, _26549_, _26548_);
  nand (_26551_, _26550_, _26543_);
  or (_26552_, _26550_, _26543_);
  and (_26553_, _26552_, _26551_);
  nand (_26554_, _26553_, _26542_);
  or (_26555_, _26553_, _26542_);
  nand (_26556_, _26555_, _26554_);
  not (_26557_, _26556_);
  and (_26558_, _26557_, _26541_);
  nor (_26559_, _26557_, _26541_);
  nor (_26560_, _26559_, _26558_);
  and (_26561_, _26560_, _23531_);
  and (_26562_, _26384_, _22995_);
  and (_26563_, _23488_, _23456_);
  nand (_26564_, _23534_, _23264_);
  nand (_26565_, _24206_, _26564_);
  or (_26566_, _26565_, _26563_);
  or (_26567_, _26566_, _26562_);
  nor (_26568_, _26567_, _26561_);
  and (_26569_, _26568_, _26392_);
  nand (_26570_, _26569_, _26382_);
  not (_26571_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_26572_, \oc8051_top_1.oc8051_decoder1.state [1], _22735_);
  and (_26573_, _26572_, _26571_);
  and (_26574_, _24251_, _26573_);
  not (_26575_, _26573_);
  and (_26576_, _23816_, _23772_);
  nor (_26577_, _26576_, _24251_);
  and (_26578_, _23825_, _23805_);
  or (_26579_, _23898_, _23807_);
  nor (_26580_, _26579_, _26578_);
  and (_26581_, _23818_, _23816_);
  and (_26582_, _23903_, _23816_);
  nor (_26583_, _26582_, _26581_);
  and (_26584_, _23816_, _23810_);
  nor (_26585_, _26584_, _23897_);
  and (_26586_, _26585_, _26583_);
  and (_26587_, _26586_, _26580_);
  and (_26588_, _26587_, _26577_);
  nor (_26589_, _26588_, _26575_);
  and (_26590_, _23816_, _24278_);
  and (_26591_, _26590_, _23903_);
  nor (_26592_, _26591_, _26589_);
  and (_26593_, _23802_, _23778_);
  and (_26594_, _23800_, _23792_);
  nor (_26595_, _26594_, _26593_);
  nor (_26596_, _26595_, _24279_);
  nor (_26597_, _26574_, _26596_);
  or (_26598_, _26579_, _23897_);
  nand (_26599_, _26598_, _26573_);
  or (_26600_, _26583_, _26575_);
  and (_26601_, \oc8051_top_1.oc8051_decoder1.state [0], _22735_);
  and (_26602_, _26601_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_26603_, _23903_, _23792_);
  and (_26605_, _26603_, _26602_);
  and (_26606_, _26594_, _24278_);
  nor (_26607_, _26606_, _26605_);
  not (_26608_, _26591_);
  and (_26609_, _26608_, _26607_);
  and (_26610_, _26609_, _26600_);
  and (_26611_, _26610_, _26599_);
  and (_26612_, _26611_, _26597_);
  and (_26613_, _26612_, _26592_);
  or (_26614_, _26613_, _26574_);
  and (_26615_, _26614_, _26570_);
  nor (_26616_, _22737_, _23280_);
  and (_26617_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_26618_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_26619_, _26618_, _26617_);
  and (_26620_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_26622_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_26623_, _26622_, _26620_);
  and (_26624_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_26625_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_26626_, _26625_, _26624_);
  and (_26627_, _26626_, _26623_);
  and (_26628_, _26627_, _26619_);
  nor (_26629_, _26628_, _24471_);
  nor (_26630_, _26629_, _26616_);
  not (_26631_, _26630_);
  nand (_26632_, _26582_, _24278_);
  and (_26633_, _26632_, _26600_);
  and (_26634_, _26607_, _26599_);
  nand (_26635_, _26634_, _26633_);
  or (_26636_, _26635_, _26631_);
  and (_26637_, _26634_, _26633_);
  nor (_26638_, _22737_, _23278_);
  or (_26639_, _23623_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_26640_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_26641_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_26642_, _26641_, _26640_);
  and (_26643_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_26644_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_26645_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_26646_, _26645_, _26644_);
  or (_26647_, _26646_, _26643_);
  or (_26648_, _26647_, _26642_);
  and (_26649_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_26650_, _26649_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_26651_, _26650_, _26648_);
  and (_26652_, _26651_, _22737_);
  and (_26653_, _26652_, _26639_);
  nor (_26654_, _26653_, _26638_);
  not (_26655_, _26654_);
  or (_26656_, _26655_, _26637_);
  and (_26657_, _26656_, _26636_);
  and (_26658_, _26657_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_26659_, _26657_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_26660_, _26635_, _26597_);
  nor (_26662_, _26660_, _26592_);
  nand (_26663_, _26662_, _26659_);
  nor (_26664_, _26663_, _26658_);
  and (_26665_, _26660_, _26592_);
  and (_26666_, _26665_, _26631_);
  and (_26667_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_26668_, _26667_, _26666_);
  or (_26669_, _26668_, _26664_);
  or (_26670_, _26669_, _26615_);
  nor (_26671_, _26583_, _26601_);
  and (_26672_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_26673_, _23911_, _23780_);
  nor (_26674_, _24255_, _26673_);
  nor (_26675_, _24244_, _23773_);
  and (_26676_, _26675_, _26674_);
  nor (_26677_, _26676_, _24279_);
  and (_26678_, _26584_, _26573_);
  not (_26679_, _22736_);
  nor (_26680_, _26675_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_26681_, _26680_, _26679_);
  nor (_26682_, _26681_, _26678_);
  not (_26683_, _26682_);
  nor (_26684_, _26683_, _26677_);
  nor (_26686_, _26684_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_26687_, _26686_, _26672_);
  and (_26688_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_26689_, _26688_);
  and (_26690_, _23816_, _23806_);
  and (_26691_, _23814_, _23772_);
  nor (_26692_, _26691_, _26690_);
  and (_26693_, _23788_, _23708_);
  and (_26694_, _26693_, _23814_);
  nor (_26695_, _26694_, _26603_);
  and (_26696_, _26695_, _26692_);
  nor (_26697_, _23910_, _23841_);
  and (_26698_, _23810_, _23708_);
  nand (_26699_, _26698_, _23814_);
  and (_26700_, _26699_, _26697_);
  and (_26701_, _23814_, _23784_);
  nor (_26702_, _26701_, _23840_);
  not (_26703_, _26702_);
  nor (_26704_, _26703_, _24269_);
  and (_26705_, _26704_, _26700_);
  and (_26706_, _26705_, _26696_);
  nand (_26707_, _26706_, _26674_);
  nand (_26708_, _26707_, _24278_);
  and (_26709_, _26678_, _23769_);
  nor (_26710_, _26709_, _26671_);
  and (_26711_, _26710_, _26678_);
  nor (_26712_, _26711_, _26605_);
  nand (_26713_, _26712_, _26708_);
  nand (_26714_, _26713_, _22735_);
  and (_26715_, _26714_, _26689_);
  not (_26716_, _26715_);
  and (_26717_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_26718_, _26717_);
  nor (_26719_, _24274_, _23930_);
  and (_26720_, _26719_, _24260_);
  and (_26721_, _23838_, _23783_);
  not (_26722_, _26721_);
  and (_26723_, _23801_, _23803_);
  and (_26724_, _23803_, _23772_);
  nor (_26726_, _26724_, _26723_);
  and (_26727_, _26726_, _26722_);
  and (_26729_, _26727_, _26720_);
  and (_26730_, _23926_, _23708_);
  and (_26731_, _26730_, _23797_);
  and (_26732_, _26731_, _23685_);
  nor (_26733_, _26732_, _23845_);
  and (_26734_, _23911_, _23792_);
  and (_26735_, _23923_, _23791_);
  nor (_26736_, _26735_, _26734_);
  and (_26737_, _26736_, _26733_);
  and (_26738_, _26737_, _26729_);
  or (_26739_, _23819_, _23807_);
  nand (_26740_, _26739_, _23685_);
  not (_26741_, _23817_);
  and (_26742_, _23844_, _23792_);
  nor (_26743_, _26742_, _23793_);
  and (_26744_, _26743_, _26741_);
  and (_26745_, _26744_, _26740_);
  not (_26747_, _23803_);
  nor (_26748_, _23903_, _23812_);
  nor (_26749_, _26748_, _26747_);
  or (_26750_, _23911_, _23784_);
  nand (_26751_, _26750_, _23803_);
  nand (_26752_, _26751_, _26583_);
  nor (_26753_, _26752_, _26749_);
  and (_26754_, _26693_, _23803_);
  nor (_26755_, _26754_, _26603_);
  and (_26756_, _23892_, _23814_);
  and (_26757_, _26730_, _23779_);
  nor (_26758_, _26757_, _26756_);
  and (_26759_, _26758_, _26755_);
  and (_26760_, _23816_, _23805_);
  nor (_26761_, _26760_, _23893_);
  and (_26762_, _26761_, _24265_);
  and (_26763_, _26762_, _26759_);
  and (_26764_, _26763_, _26753_);
  and (_26765_, _26764_, _26745_);
  nand (_26766_, _26765_, _26738_);
  nand (_26767_, _26766_, _24278_);
  nor (_26768_, _26605_, _26678_);
  nand (_26769_, _26768_, _26767_);
  nand (_26770_, _26769_, _22735_);
  and (_26772_, _26770_, _26718_);
  and (_26773_, _26772_, _26716_);
  and (_26775_, _26773_, _26687_);
  nand (_26776_, _26775_, _25954_);
  nor (_26777_, _26772_, _26715_);
  and (_26778_, _26777_, _26687_);
  and (_26779_, _24177_, _22867_);
  and (_26780_, _26779_, _24188_);
  and (_26781_, _26780_, _23577_);
  and (_26782_, _26780_, _23880_);
  not (_26783_, _26780_);
  and (_26784_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_26786_, _26784_, _26782_);
  and (_26787_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_26788_, _26783_, _23542_);
  nor (_26789_, _26788_, _26787_);
  nand (_26790_, _26780_, _24671_);
  or (_26791_, _26780_, _22874_);
  and (_26792_, _26791_, _26790_);
  and (_26793_, _26792_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_26794_, _26793_, _26789_);
  and (_26795_, _26794_, _26786_);
  and (_26796_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_26797_, _26796_, _26781_);
  and (_26798_, _26797_, _26795_);
  nor (_26799_, _26797_, _26795_);
  nor (_26800_, _26799_, _26798_);
  nor (_26801_, _26800_, _22815_);
  nor (_26802_, _26801_, _22857_);
  nor (_26803_, _26802_, _26780_);
  nor (_26804_, _26803_, _26781_);
  not (_26805_, _26804_);
  nand (_26806_, _26805_, _26778_);
  and (_26807_, _26715_, _26687_);
  and (_26808_, _26807_, _26772_);
  nand (_26809_, _26808_, _25687_);
  not (_26810_, _24473_);
  not (_26811_, _26772_);
  and (_26812_, _26807_, _26811_);
  nand (_26813_, _26812_, _26810_);
  and (_26814_, _26813_, _26809_);
  and (_26815_, _26814_, _26806_);
  and (_26816_, _26815_, _26776_);
  nor (_26818_, _26816_, _22867_);
  and (_26819_, _26816_, _22867_);
  nor (_26820_, _26819_, _26818_);
  not (_26821_, _26820_);
  and (_00001_, _26775_, _25976_);
  not (_00002_, _00001_);
  not (_00003_, _26778_);
  nor (_00004_, _26783_, _24082_);
  and (_00005_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_00006_, _00005_, _00004_);
  and (_00008_, _00006_, _26798_);
  nor (_00009_, _00006_, _26798_);
  nor (_00010_, _00009_, _00008_);
  nor (_00011_, _00010_, _22815_);
  nor (_00012_, _00011_, _22896_);
  nor (_00013_, _00012_, _26780_);
  nor (_00014_, _00013_, _00004_);
  nor (_00015_, _00014_, _00003_);
  and (_00016_, _26808_, _25855_);
  not (_00017_, _00016_);
  or (_00018_, _26772_, _26716_);
  nor (_00020_, _00018_, _25577_);
  not (_00021_, _26687_);
  and (_00023_, _26715_, _00021_);
  nor (_00024_, _00023_, _00020_);
  nand (_00025_, _00024_, _00017_);
  nor (_00026_, _00025_, _00015_);
  and (_00027_, _00026_, _00002_);
  nor (_00028_, _00027_, _22905_);
  and (_00029_, _00027_, _22905_);
  nor (_00030_, _00029_, _00028_);
  and (_00031_, _26775_, _25995_);
  not (_00033_, _26050_);
  and (_00034_, _26812_, _00033_);
  nor (_00035_, _00034_, _00031_);
  nor (_00036_, _26783_, _24043_);
  and (_00037_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_00038_, _00037_, _00036_);
  and (_00039_, _00038_, _00008_);
  nor (_00040_, _00038_, _00008_);
  nor (_00041_, _00040_, _00039_);
  nor (_00042_, _00041_, _22815_);
  nor (_00043_, _00042_, _22927_);
  nor (_00045_, _00043_, _26780_);
  nor (_00046_, _00045_, _00036_);
  nor (_00047_, _00046_, _00003_);
  nor (_00048_, _26773_, _26687_);
  and (_00049_, _00048_, _00018_);
  nor (_00050_, _00049_, _00047_);
  and (_00051_, _00050_, _00035_);
  nor (_00052_, _00051_, _22936_);
  and (_00053_, _00051_, _22936_);
  nor (_00054_, _00053_, _00052_);
  nor (_00055_, _00054_, _00030_);
  nor (_00056_, _22737_, _23062_);
  and (_00057_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00058_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_00059_, _00058_, _00057_);
  and (_00060_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00061_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_00062_, _00061_, _00060_);
  and (_00063_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_00064_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_00065_, _00064_, _00063_);
  and (_00066_, _00065_, _00062_);
  and (_00067_, _00066_, _00059_);
  nor (_00068_, _00067_, _24471_);
  nor (_00069_, _00068_, _00056_);
  not (_00070_, _00069_);
  and (_00071_, _00070_, _26812_);
  nor (_00072_, _26783_, _24126_);
  and (_00073_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_00075_, _00073_, _00072_);
  and (_00076_, _00075_, _00039_);
  nor (_00077_, _00075_, _00039_);
  nor (_00078_, _00077_, _00076_);
  nor (_00080_, _00078_, _22815_);
  nor (_00081_, _00080_, _22960_);
  nor (_00083_, _00081_, _26780_);
  nor (_00084_, _00083_, _00072_);
  nor (_00085_, _00084_, _00003_);
  and (_00086_, _26775_, _26018_);
  or (_00088_, _00048_, _00086_);
  or (_00089_, _00088_, _00085_);
  nor (_00090_, _00089_, _00071_);
  nor (_00091_, _00090_, _22968_);
  and (_00092_, _00090_, _22968_);
  nor (_00093_, _00092_, _00091_);
  and (_00094_, _26783_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nand (_00095_, _00094_, _00076_);
  or (_00096_, _00094_, _00076_);
  and (_00097_, _00096_, _22854_);
  nand (_00098_, _00097_, _00095_);
  nor (_00099_, _26780_, _22826_);
  nand (_00100_, _00099_, _00098_);
  and (_00101_, _26780_, _23989_);
  not (_00102_, _00101_);
  nand (_00104_, _00102_, _00100_);
  not (_00105_, _00104_);
  nand (_00106_, _00105_, _26777_);
  nand (_00107_, _25852_, _23989_);
  nand (_00108_, _25865_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand (_00109_, _25877_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_00110_, _00109_, _00108_);
  nand (_00111_, _25858_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nand (_00112_, _25882_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_00113_, _00112_, _00111_);
  and (_00114_, _00113_, _00110_);
  nand (_00115_, _25867_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand (_00116_, _25861_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_00117_, _00116_, _00115_);
  nand (_00118_, _25874_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nand (_00119_, _25880_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_00120_, _00119_, _00118_);
  and (_00121_, _00120_, _00117_);
  and (_00122_, _00121_, _25872_);
  nand (_00123_, _00122_, _00114_);
  and (_00124_, _00123_, _00107_);
  nand (_00125_, _00124_, _26773_);
  nor (_00126_, _22737_, _23008_);
  and (_00127_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00128_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_00129_, _00128_, _00127_);
  and (_00130_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00131_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_00132_, _00131_, _00130_);
  and (_00133_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_00134_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_00135_, _00134_, _00133_);
  and (_00136_, _00135_, _00132_);
  and (_00137_, _00136_, _00129_);
  nor (_00138_, _00137_, _24471_);
  nor (_00139_, _00138_, _00126_);
  or (_00140_, _00139_, _00018_);
  and (_00141_, _00140_, _26687_);
  and (_00142_, _00141_, _00125_);
  nand (_00143_, _00142_, _00106_);
  and (_00144_, _00143_, _22844_);
  nor (_00145_, _00143_, _22844_);
  nor (_00146_, _00145_, _00144_);
  nor (_00147_, _00146_, _00093_);
  and (_00148_, _00147_, _00055_);
  and (_00149_, _00148_, _26821_);
  nor (_00150_, _25481_, _24180_);
  and (_00151_, _00150_, _00149_);
  and (_00152_, _00151_, _26671_);
  not (_00153_, _00152_);
  and (_00154_, _26775_, _25911_);
  not (_00155_, _00154_);
  and (_00156_, _26808_, _23664_);
  not (_00157_, _26068_);
  and (_00158_, _26812_, _00157_);
  nor (_00159_, _00158_, _00156_);
  and (_00160_, _26773_, _00021_);
  nor (_00161_, _26793_, _26789_);
  nor (_00162_, _00161_, _26794_);
  nor (_00163_, _00162_, _22815_);
  nor (_00164_, _00163_, _22911_);
  nor (_00165_, _00164_, _26780_);
  nor (_00166_, _00165_, _26788_);
  not (_00167_, _00166_);
  and (_00168_, _00167_, _26778_);
  nor (_00169_, _00168_, _00160_);
  and (_00170_, _00169_, _00159_);
  and (_00171_, _00170_, _00155_);
  nor (_00173_, _00171_, _22919_);
  and (_00174_, _00171_, _22919_);
  nor (_00175_, _00174_, _00173_);
  or (_00176_, _26820_, _25113_);
  and (_00177_, _26775_, _25891_);
  and (_00178_, _26631_, _26812_);
  nor (_00179_, _00178_, _00177_);
  nor (_00180_, _26792_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_00181_, _00180_, _26793_);
  nor (_00182_, _00181_, _22815_);
  nor (_00183_, _00182_, _22875_);
  nor (_00185_, _00183_, _26780_);
  not (_00186_, _00185_);
  and (_00187_, _00186_, _26790_);
  nor (_00188_, _00187_, _00003_);
  and (_00189_, _26808_, _23685_);
  nor (_00190_, _00189_, _00188_);
  and (_00191_, _00190_, _00179_);
  and (_00192_, _00191_, _24175_);
  nor (_00193_, _00191_, _24175_);
  or (_00194_, _00193_, _00192_);
  and (_00195_, _26775_, _25930_);
  not (_00196_, _00195_);
  and (_00197_, _26808_, _23643_);
  nor (_00198_, _26794_, _26786_);
  nor (_00199_, _00198_, _26795_);
  nor (_00200_, _00199_, _22815_);
  nor (_00201_, _00200_, _22942_);
  nor (_00202_, _00201_, _26780_);
  nor (_00204_, _00202_, _26782_);
  not (_00205_, _00204_);
  and (_00206_, _00205_, _26778_);
  nor (_00207_, _22737_, _23226_);
  and (_00208_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00210_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_00211_, _00210_, _00208_);
  and (_00213_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00214_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_00216_, _00214_, _00213_);
  and (_00217_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_00218_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_00219_, _00218_, _00217_);
  and (_00220_, _00219_, _00216_);
  and (_00221_, _00220_, _00211_);
  nor (_00222_, _00221_, _24471_);
  nor (_00223_, _00222_, _00207_);
  not (_00224_, _00223_);
  and (_00225_, _00224_, _26812_);
  or (_00226_, _00225_, _00206_);
  nor (_00227_, _00226_, _00197_);
  and (_00228_, _00227_, _00196_);
  nor (_00229_, _00228_, _22951_);
  and (_00230_, _00228_, _22951_);
  nor (_00231_, _00230_, _00229_);
  or (_00232_, _00231_, _00194_);
  or (_00233_, _00232_, _00176_);
  nor (_00234_, _00233_, _00175_);
  and (_00235_, _00234_, _00148_);
  and (_00236_, _22844_, _22869_);
  and (_00237_, _00236_, _00235_);
  and (_00238_, _26698_, _23816_);
  and (_00239_, _26582_, _23708_);
  or (_00240_, _00239_, _26581_);
  and (_00241_, _23380_, _23393_);
  nor (_00242_, _23380_, _23393_);
  nor (_00243_, _00242_, _00241_);
  not (_00244_, _00243_);
  nor (_00245_, _23376_, _23173_);
  and (_00246_, _23376_, _23173_);
  nor (_00247_, _00246_, _00245_);
  and (_00248_, _23369_, _23316_);
  nor (_00249_, _00248_, _23370_);
  nor (_00250_, _23367_, _23319_);
  nor (_00251_, _00250_, _23368_);
  nor (_00252_, _26678_, _23321_);
  and (_00253_, _00252_, _00251_);
  nand (_00254_, _00253_, _00249_);
  nor (_00255_, _00254_, _00247_);
  not (_00256_, _26384_);
  nor (_00257_, _23377_, _23168_);
  nor (_00258_, _00257_, _23378_);
  and (_00259_, _00258_, _00256_);
  and (_00260_, _00259_, _00255_);
  nor (_00261_, _23378_, _23164_);
  nor (_00263_, _00261_, _23379_);
  and (_00264_, _00263_, _26710_);
  and (_00265_, _00264_, _00260_);
  and (_00266_, _00265_, _00244_);
  not (_00267_, _00266_);
  and (_00268_, _26709_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  not (_00269_, _00268_);
  and (_00271_, _26671_, _23478_);
  nor (_00272_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_00273_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00274_, _00273_, _00272_);
  nor (_00275_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_00277_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_00278_, _00277_, _00275_);
  and (_00279_, _00278_, _00274_);
  and (_00281_, _00279_, _26711_);
  nor (_00282_, _00281_, _00271_);
  and (_00283_, _00282_, _00269_);
  and (_00284_, _00283_, _00267_);
  or (_00285_, _00284_, _00240_);
  nor (_00286_, _00285_, _00238_);
  and (_00287_, _26582_, _23707_);
  not (_00288_, _00287_);
  and (_00290_, _26584_, _23707_);
  nor (_00292_, _00290_, _23897_);
  and (_00293_, _00292_, _00288_);
  and (_00294_, _00293_, _26580_);
  and (_00295_, _00294_, _00284_);
  nor (_00296_, _00295_, _00286_);
  not (_00297_, _26603_);
  and (_00298_, _26577_, _00297_);
  not (_00300_, _00298_);
  nor (_00301_, _00300_, _00296_);
  nor (_00303_, _26605_, _26573_);
  nor (_00304_, _00303_, _00301_);
  nor (_00306_, _00304_, _26596_);
  and (_00307_, _25478_, _24539_);
  and (_00308_, _00307_, _25017_);
  not (_00309_, _00308_);
  nor (_00311_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not (_00312_, _00311_);
  nor (_00313_, _00312_, _25683_);
  and (_00314_, _00313_, _00309_);
  not (_00315_, _00314_);
  and (_00316_, _00315_, _26709_);
  not (_00317_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_00318_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _22735_);
  and (_00319_, _00318_, _00317_);
  not (_00320_, _00319_);
  nor (_00321_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00322_, _00321_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_00323_, _24625_, _24004_);
  and (_00324_, _00323_, _25681_);
  nor (_00325_, _00324_, _00322_);
  and (_00326_, _00325_, _00320_);
  nor (_00327_, _22968_, _22936_);
  and (_00328_, _00327_, _24539_);
  and (_00329_, _00328_, _25123_);
  not (_00330_, _00329_);
  and (_00331_, _00330_, _00326_);
  not (_00332_, _00331_);
  and (_00333_, _00332_, _26711_);
  nor (_00334_, _00333_, _00316_);
  not (_00335_, _00334_);
  nor (_00336_, _00335_, _00306_);
  not (_00337_, _00336_);
  nor (_00338_, _00337_, _00237_);
  and (_00339_, _00338_, _00153_);
  nand (_00340_, _26655_, _26606_);
  nand (_00341_, _00340_, _00339_);
  or (_00342_, _00341_, _26670_);
  or (_00343_, _00339_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_00344_, _00343_, _22731_);
  and (_26870_[0], _00344_, _00342_);
  or (_00345_, _00339_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_00346_, _00345_, _22731_);
  nand (_00347_, _26376_, _26184_);
  or (_00348_, _26350_, _26348_);
  and (_00349_, _00348_, _26351_);
  or (_00350_, _00349_, _00347_);
  or (_00351_, _26377_, _26345_);
  and (_00352_, _00351_, _00350_);
  nand (_00353_, _00352_, _23528_);
  and (_00354_, _26553_, _26542_);
  nor (_00355_, _26558_, _00354_);
  and (_00356_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  and (_00357_, _26548_, _26484_);
  nand (_00358_, _00357_, _26551_);
  nand (_00359_, _00358_, _00356_);
  or (_00360_, _00358_, _00356_);
  nand (_00361_, _00360_, _00359_);
  nand (_00362_, _00361_, _00355_);
  or (_00363_, _00361_, _00355_);
  and (_00364_, _00363_, _00362_);
  nand (_00365_, _00364_, _23531_);
  nor (_00366_, _23463_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_00367_, _00366_, _23264_);
  nor (_00368_, _00366_, _23264_);
  nor (_00369_, _00368_, _00367_);
  nor (_00370_, _00369_, _23470_);
  not (_00371_, _00370_);
  nand (_00372_, _23534_, _23232_);
  and (_00373_, _23484_, _23264_);
  not (_00374_, _23535_);
  nor (_00375_, _00374_, _23296_);
  nor (_00376_, _00375_, _00373_);
  and (_00377_, _00376_, _00372_);
  and (_00378_, _00377_, _23527_);
  and (_00379_, _00378_, _00371_);
  and (_00380_, _00379_, _23518_);
  nor (_00381_, _23324_, _23272_);
  or (_00382_, _00381_, _23396_);
  and (_00383_, _00382_, _23404_);
  nor (_00384_, _00382_, _23404_);
  or (_00385_, _00384_, _00383_);
  and (_00386_, _00385_, _23390_);
  nor (_00387_, _23366_, _23322_);
  nor (_00388_, _00387_, _23367_);
  nor (_00389_, _00388_, _22996_);
  nor (_00390_, _00389_, _00386_);
  and (_00391_, _00390_, _00380_);
  and (_00392_, _00391_, _00365_);
  nand (_00393_, _00392_, _00353_);
  and (_00394_, _00393_, _26614_);
  and (_00395_, _26665_, _00157_);
  and (_00396_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_00397_, _00396_, _00395_);
  or (_00398_, _26635_, _00157_);
  nor (_00399_, _22737_, _23246_);
  and (_00400_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_00401_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00402_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00403_, _00402_, _00401_);
  and (_00404_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00405_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_00406_, _00405_, _00404_);
  or (_00407_, _00406_, _00403_);
  and (_00408_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00409_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00410_, _00409_, _00408_);
  or (_00411_, _00410_, _00407_);
  and (_00412_, _00411_, _23623_);
  or (_00413_, _00412_, _00400_);
  and (_00414_, _00413_, _22737_);
  nor (_00415_, _00414_, _00399_);
  not (_00416_, _00415_);
  or (_00417_, _00416_, _26637_);
  and (_00418_, _00417_, _00398_);
  nand (_00419_, _00418_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_00420_, _00418_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_00421_, _00420_, _00419_);
  or (_00422_, _00421_, _26658_);
  and (_00423_, _00421_, _26658_);
  not (_00424_, _00423_);
  and (_00425_, _00424_, _26662_);
  and (_00426_, _00425_, _00422_);
  or (_00427_, _00426_, _00397_);
  or (_00428_, _00427_, _00394_);
  nand (_00429_, _00416_, _26606_);
  nand (_00430_, _00429_, _00339_);
  or (_00431_, _00430_, _00428_);
  and (_26870_[1], _00431_, _00346_);
  not (_00432_, _26363_);
  and (_00433_, _26362_, _26352_);
  nor (_00434_, _00433_, _00432_);
  or (_00435_, _00434_, _00347_);
  or (_00436_, _26377_, _26358_);
  and (_00437_, _00436_, _00435_);
  nand (_00438_, _00437_, _23528_);
  and (_00439_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  not (_00440_, _26541_);
  or (_00441_, _00361_, _26556_);
  or (_00442_, _00441_, _00440_);
  nand (_00443_, _00360_, _00354_);
  and (_00444_, _00443_, _00359_);
  and (_00445_, _00444_, _00442_);
  not (_00446_, _00445_);
  nand (_00447_, _00446_, _00439_);
  or (_00448_, _00446_, _00439_);
  and (_00449_, _00448_, _00447_);
  nand (_00450_, _00449_, _23531_);
  nor (_00451_, _00251_, _22996_);
  and (_00452_, _23484_, _23232_);
  not (_00453_, _00452_);
  nand (_00454_, _23535_, _23264_);
  not (_00455_, _23534_);
  or (_00456_, _00455_, _23199_);
  and (_00457_, _00456_, _00454_);
  and (_00458_, _00457_, _00453_);
  and (_00459_, _00458_, _23876_);
  not (_00460_, _00459_);
  nor (_00461_, _00460_, _00451_);
  nor (_00462_, _23407_, _23405_);
  nor (_00463_, _00462_, _23391_);
  and (_00464_, _00463_, _23409_);
  and (_00465_, _23462_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_00466_, _00368_, _23872_);
  nor (_00467_, _00466_, _00465_);
  nor (_00468_, _00467_, _23470_);
  nor (_00469_, _00468_, _00464_);
  and (_00470_, _00469_, _00461_);
  and (_00471_, _00470_, _23868_);
  and (_00472_, _00471_, _00450_);
  nand (_00473_, _00472_, _00438_);
  and (_00474_, _00473_, _26614_);
  and (_00475_, _26665_, _00224_);
  and (_00476_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_00477_, _00476_, _00475_);
  nand (_00478_, _00424_, _00419_);
  or (_00479_, _26635_, _00224_);
  nor (_00480_, _22737_, _23228_);
  and (_00481_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_00482_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00483_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_00484_, _00483_, _00482_);
  and (_00485_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00486_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_00487_, _00486_, _00485_);
  and (_00488_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00489_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_00490_, _00489_, _00488_);
  and (_00491_, _00490_, _00487_);
  and (_00492_, _00491_, _00484_);
  nor (_00493_, _00492_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_00494_, _00493_, _00481_);
  nor (_00495_, _00494_, _25454_);
  nor (_00496_, _00495_, _00480_);
  not (_00497_, _00496_);
  or (_00498_, _00497_, _26637_);
  nand (_00499_, _00498_, _00479_);
  or (_00500_, _00499_, _23213_);
  nand (_00501_, _00499_, _23213_);
  and (_00502_, _00501_, _00500_);
  or (_00503_, _00502_, _00478_);
  and (_00504_, _00502_, _00478_);
  not (_00505_, _00504_);
  and (_00506_, _00505_, _26662_);
  and (_00507_, _00506_, _00503_);
  or (_00508_, _00507_, _00477_);
  or (_00509_, _00508_, _00474_);
  nand (_00510_, _00497_, _26606_);
  nand (_00511_, _00510_, _00339_);
  or (_00512_, _00511_, _00509_);
  not (_00513_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00514_, _25694_, _00513_);
  and (_00516_, _25694_, _00513_);
  nor (_00517_, _00516_, _00514_);
  or (_00518_, _00517_, _00339_);
  and (_00519_, _00518_, _22731_);
  and (_26870_[2], _00519_, _00512_);
  and (_00520_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_00521_, _00520_, _00439_);
  not (_00522_, _00521_);
  nor (_00523_, _00522_, _00444_);
  nor (_00524_, _00522_, _00441_);
  and (_00525_, _00524_, _26541_);
  nor (_00526_, _00525_, _00523_);
  not (_00528_, _00520_);
  nand (_00529_, _00528_, _00447_);
  and (_00530_, _00529_, _00526_);
  nand (_00531_, _00530_, _23531_);
  not (_00532_, _26338_);
  or (_00533_, _26377_, _00532_);
  or (_00534_, _26364_, _26339_);
  and (_00535_, _26363_, _26359_);
  nand (_00536_, _00535_, _00534_);
  or (_00537_, _00535_, _00534_);
  and (_00538_, _00537_, _00536_);
  nand (_00539_, _00538_, _26377_);
  nand (_00540_, _00539_, _00533_);
  nand (_00542_, _00540_, _23528_);
  nor (_00543_, _00249_, _22996_);
  not (_00544_, _00543_);
  not (_00545_, _23463_);
  not (_00546_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_00547_, _23462_, _00546_);
  nor (_00548_, _00547_, _23563_);
  nor (_00549_, _00548_, _23470_);
  and (_00550_, _00549_, _00545_);
  not (_00551_, _00550_);
  and (_00552_, _23409_, _23402_);
  or (_00553_, _00552_, _23391_);
  nor (_00554_, _00553_, _23410_);
  not (_00555_, _00554_);
  or (_00556_, _00455_, _23150_);
  and (_00557_, _23484_, _23563_);
  nand (_00558_, _23535_, _23232_);
  not (_00559_, _00558_);
  nor (_00560_, _00559_, _00557_);
  and (_00561_, _00560_, _00556_);
  and (_00562_, _00561_, _23561_);
  not (_00563_, _00562_);
  nor (_00564_, _00563_, _23575_);
  and (_00565_, _00564_, _00555_);
  and (_00566_, _00565_, _00551_);
  and (_00567_, _00566_, _00544_);
  and (_00568_, _00567_, _00542_);
  nand (_00569_, _00568_, _00531_);
  and (_00570_, _00569_, _26614_);
  and (_00571_, _26665_, _26810_);
  and (_00572_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_00573_, _00572_, _00571_);
  nand (_00574_, _00505_, _00500_);
  and (_00575_, _26637_, _24473_);
  nor (_00576_, _22737_, _23181_);
  and (_00577_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_00578_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00579_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_00580_, _00579_, _00578_);
  and (_00581_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00582_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or (_00583_, _00582_, _00581_);
  or (_00584_, _00583_, _00580_);
  and (_00585_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00586_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_00587_, _00586_, _00585_);
  or (_00588_, _00587_, _00584_);
  and (_00589_, _00588_, _23623_);
  or (_00590_, _00589_, _00577_);
  and (_00591_, _00590_, _22737_);
  nor (_00592_, _00591_, _00576_);
  and (_00593_, _00592_, _26635_);
  nor (_00594_, _00593_, _00575_);
  and (_00595_, _00594_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_00597_, _00594_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_00598_, _00597_, _00595_);
  nand (_00599_, _00598_, _00574_);
  or (_00600_, _00598_, _00574_);
  and (_00601_, _00600_, _26662_);
  and (_00602_, _00601_, _00599_);
  or (_00603_, _00602_, _00573_);
  or (_00604_, _00603_, _00570_);
  not (_00605_, _00592_);
  nand (_00606_, _00605_, _26606_);
  nand (_00607_, _00606_, _00339_);
  or (_00608_, _00607_, _00604_);
  and (_00609_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  not (_00610_, _00609_);
  nor (_00611_, _00610_, _25694_);
  nor (_00612_, _00514_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00613_, _00612_, _00611_);
  or (_00614_, _00613_, _00339_);
  and (_00615_, _00614_, _22731_);
  and (_26870_[3], _00615_, _00608_);
  nand (_00616_, _26370_, _26368_);
  or (_00617_, _26370_, _26368_);
  nand (_00618_, _00617_, _00616_);
  nand (_00619_, _00618_, _26377_);
  or (_00620_, _26377_, _26326_);
  and (_00621_, _00620_, _00619_);
  nand (_00622_, _00621_, _23528_);
  or (_00623_, _00525_, _00523_);
  and (_00624_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  nand (_00625_, _00624_, _00623_);
  or (_00626_, _00624_, _00623_);
  and (_00627_, _00626_, _00625_);
  nand (_00628_, _00627_, _23531_);
  and (_00629_, _00247_, _22995_);
  not (_00630_, _00629_);
  nor (_00631_, _23413_, _23173_);
  not (_00632_, _00631_);
  nor (_00633_, _23414_, _23391_);
  and (_00634_, _00633_, _00632_);
  not (_00635_, _00634_);
  and (_00636_, _23484_, _23460_);
  not (_00637_, _00636_);
  or (_00638_, _00374_, _23199_);
  nand (_00639_, _23534_, _23115_);
  and (_00640_, _00639_, _00638_);
  and (_00641_, _00640_, _00637_);
  nand (_00642_, _00641_, _24075_);
  nor (_00643_, _23464_, _23460_);
  not (_00644_, _00643_);
  nor (_00645_, _23465_, _23470_);
  and (_00646_, _00645_, _00644_);
  not (_00647_, _00646_);
  nand (_00648_, _00647_, _24072_);
  or (_00649_, _00648_, _00642_);
  nor (_00650_, _00649_, _24079_);
  and (_00651_, _00650_, _00635_);
  and (_00652_, _00651_, _00630_);
  and (_00653_, _00652_, _00628_);
  nand (_00654_, _00653_, _00622_);
  and (_00655_, _00654_, _26614_);
  not (_00656_, _25577_);
  and (_00658_, _26665_, _00656_);
  nor (_00659_, _22737_, _23131_);
  and (_00660_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_00661_, _23593_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00662_, _23602_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00663_, _00662_, _00661_);
  and (_00664_, _23607_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00665_, _23597_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_00666_, _00665_, _00664_);
  or (_00667_, _00666_, _00663_);
  and (_00668_, _23605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00669_, _23590_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00670_, _00669_, _00668_);
  or (_00671_, _00670_, _00667_);
  and (_00672_, _00671_, _23623_);
  or (_00673_, _00672_, _00660_);
  and (_00675_, _00673_, _22737_);
  nor (_00676_, _00675_, _00659_);
  not (_00677_, _00676_);
  and (_00678_, _00677_, _26606_);
  and (_00679_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00680_, _00679_, _00678_);
  or (_00681_, _00680_, _00658_);
  and (_00682_, _26637_, _25577_);
  and (_00683_, _00676_, _26635_);
  nor (_00684_, _00683_, _00682_);
  nand (_00685_, _00684_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_00686_, _00684_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00687_, _00686_, _00685_);
  nor (_00688_, _00595_, _00574_);
  nor (_00689_, _00688_, _00597_);
  or (_00690_, _00689_, _00687_);
  nand (_00691_, _00689_, _00687_);
  and (_00692_, _00691_, _26662_);
  and (_00693_, _00692_, _00690_);
  nor (_00694_, _00693_, _00681_);
  nand (_00695_, _00694_, _00339_);
  or (_00696_, _00695_, _00655_);
  and (_00697_, _00611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00698_, _00611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_00699_, _00698_, _00697_);
  or (_00700_, _00699_, _00339_);
  and (_00701_, _00700_, _22731_);
  and (_26870_[4], _00701_, _00696_);
  nand (_00702_, _00347_, _26320_);
  and (_00703_, _00616_, _26328_);
  nand (_00704_, _00703_, _26371_);
  or (_00705_, _00703_, _26371_);
  nand (_00706_, _00705_, _00704_);
  nand (_00707_, _00706_, _26377_);
  nand (_00708_, _00707_, _00702_);
  nand (_00709_, _00708_, _23528_);
  and (_00710_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_00711_, _00710_, _00624_);
  nand (_00712_, _00711_, _00623_);
  not (_00713_, _00710_);
  nand (_00714_, _00713_, _00625_);
  and (_00715_, _00714_, _00712_);
  nand (_00716_, _00715_, _23531_);
  nor (_00717_, _23417_, _23414_);
  nor (_00718_, _00717_, _23418_);
  and (_00719_, _00718_, _23390_);
  not (_00720_, _00719_);
  nor (_00721_, _00258_, _22996_);
  nor (_00722_, _23458_, _23039_);
  nor (_00723_, _00722_, _23464_);
  and (_00724_, _00723_, _23364_);
  and (_00725_, _00724_, _23457_);
  not (_00726_, _00724_);
  nor (_00727_, _23465_, _23115_);
  and (_00728_, _23465_, _23115_);
  nor (_00729_, _00728_, _00727_);
  and (_00730_, _00729_, _00726_);
  or (_00731_, _00730_, _23470_);
  nor (_00732_, _00731_, _00725_);
  and (_00733_, _23484_, _23115_);
  not (_00734_, _00733_);
  or (_00735_, _00374_, _23150_);
  or (_00736_, _00455_, _23079_);
  and (_00737_, _00736_, _00735_);
  and (_00738_, _00737_, _00734_);
  and (_00739_, _00738_, _24039_);
  not (_00740_, _00739_);
  nor (_00741_, _00740_, _00732_);
  and (_00742_, _00741_, _24032_);
  not (_00743_, _00742_);
  nor (_00744_, _00743_, _00721_);
  and (_00745_, _00744_, _00720_);
  and (_00746_, _00745_, _00716_);
  nand (_00747_, _00746_, _00709_);
  and (_00748_, _00747_, _26614_);
  and (_00749_, _26665_, _00033_);
  not (_00750_, _26089_);
  and (_00751_, _26606_, _00750_);
  and (_00752_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_00753_, _00752_, _00751_);
  or (_00754_, _00753_, _00749_);
  nand (_00755_, _00691_, _00685_);
  and (_00756_, _26637_, _26050_);
  and (_00757_, _26635_, _26089_);
  nor (_00758_, _00757_, _00756_);
  and (_00759_, _00758_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_00760_, _00758_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_00761_, _00760_, _00759_);
  or (_00762_, _00761_, _00755_);
  and (_00763_, _00761_, _00755_);
  not (_00764_, _00763_);
  and (_00765_, _00764_, _26662_);
  and (_00766_, _00765_, _00762_);
  nor (_00767_, _00766_, _00754_);
  nand (_00768_, _00767_, _00339_);
  or (_00769_, _00768_, _00748_);
  and (_00770_, _00697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00771_, _00697_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00772_, _00771_, _00770_);
  or (_00773_, _00772_, _00339_);
  and (_00774_, _00773_, _22731_);
  and (_26870_[5], _00774_, _00769_);
  and (_00775_, _26374_, _26313_);
  nor (_00776_, _26374_, _26313_);
  or (_00777_, _00776_, _00775_);
  and (_00778_, _00777_, _26377_);
  nor (_00779_, _26377_, _26306_);
  or (_00780_, _00779_, _00778_);
  or (_00781_, _00780_, _23529_);
  not (_00782_, _23531_);
  and (_00783_, _26394_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  not (_00784_, _00783_);
  nor (_00785_, _00784_, _00712_);
  and (_00786_, _00784_, _00712_);
  or (_00787_, _00786_, _00785_);
  or (_00788_, _00787_, _00782_);
  nor (_00789_, _00263_, _22996_);
  not (_00790_, _00789_);
  nor (_00791_, _23423_, _23418_);
  nor (_00792_, _00791_, _23391_);
  and (_00793_, _00792_, _23425_);
  and (_00794_, _00726_, _23466_);
  and (_00795_, _00726_, _00727_);
  nor (_00796_, _00795_, _23079_);
  nor (_00797_, _00796_, _00794_);
  nor (_00798_, _00797_, _23470_);
  and (_00799_, _23484_, _23959_);
  not (_00800_, _00799_);
  or (_00801_, _00455_, _23039_);
  nand (_00802_, _23535_, _23115_);
  and (_00803_, _00802_, _00801_);
  and (_00804_, _00803_, _00800_);
  and (_00805_, _00804_, _24122_);
  not (_00806_, _00805_);
  nor (_00807_, _00806_, _00798_);
  and (_00808_, _00807_, _24115_);
  not (_00809_, _00808_);
  nor (_00810_, _00809_, _00793_);
  and (_00811_, _00810_, _00790_);
  and (_00812_, _00811_, _00788_);
  and (_00813_, _00812_, _00781_);
  not (_00814_, _00813_);
  and (_00815_, _00814_, _26614_);
  not (_00816_, _26108_);
  and (_00817_, _26606_, _00816_);
  and (_00818_, _26665_, _00070_);
  and (_00819_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00820_, _00819_, _00818_);
  or (_00821_, _00820_, _00817_);
  or (_00822_, _00763_, _00759_);
  and (_00823_, _26637_, _00069_);
  and (_00824_, _26635_, _26108_);
  nor (_00825_, _00824_, _00823_);
  nand (_00826_, _00825_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_00827_, _00825_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00828_, _00827_, _00826_);
  or (_00829_, _00828_, _00822_);
  nand (_00830_, _00828_, _00822_);
  and (_00831_, _00830_, _26662_);
  and (_00832_, _00831_, _00829_);
  or (_00833_, _00832_, _00821_);
  or (_00834_, _00833_, _00815_);
  and (_00835_, _00834_, _00339_);
  and (_00836_, _00770_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00837_, _00770_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_00838_, _00837_, _00836_);
  nor (_00839_, _00838_, _00339_);
  or (_00840_, _00839_, _00835_);
  and (_26870_[6], _00840_, _22731_);
  nor (_00841_, _00836_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_00842_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_00843_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_00844_, _00843_, _00842_);
  and (_00845_, _00844_, _00609_);
  not (_00846_, _00845_);
  nor (_00847_, _00846_, _25694_);
  nor (_00848_, _00847_, _00841_);
  or (_00849_, _00848_, _00339_);
  and (_00850_, _00849_, _22731_);
  or (_00851_, _26377_, _26298_);
  nor (_00852_, _00775_, _26307_);
  nor (_00853_, _00852_, _26311_);
  or (_00854_, _00853_, _00347_);
  and (_00855_, _00854_, _00851_);
  and (_00856_, _00855_, _23528_);
  not (_00857_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  and (_00858_, _00785_, _00857_);
  or (_00859_, _26393_, _00857_);
  nor (_00860_, _00859_, _00785_);
  or (_00861_, _00860_, _00858_);
  and (_00862_, _00861_, _23531_);
  and (_00863_, _00243_, _22995_);
  nand (_00864_, _23427_, _23393_);
  and (_00865_, _00864_, _23429_);
  and (_00866_, _00865_, _23390_);
  nor (_00867_, _00724_, _23466_);
  nor (_00868_, _00867_, _23487_);
  or (_00869_, _23467_, _23470_);
  or (_00870_, _00869_, _00868_);
  and (_00871_, _23492_, _23456_);
  nor (_00872_, _00374_, _23079_);
  and (_00873_, _23484_, _23487_);
  and (_00874_, _23441_, _23491_);
  or (_00875_, _00874_, _00873_);
  or (_00876_, _00875_, _00872_);
  nor (_00877_, _00876_, _00871_);
  and (_00878_, _00877_, _00870_);
  nand (_00879_, _00878_, _23988_);
  or (_00880_, _00879_, _00866_);
  or (_00881_, _00880_, _00863_);
  or (_00882_, _00881_, _00862_);
  or (_00883_, _00882_, _00856_);
  and (_00884_, _00883_, _26614_);
  not (_00885_, _00139_);
  and (_00886_, _26665_, _00885_);
  and (_00887_, _26605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_00888_, _00887_, _00886_);
  nand (_00889_, _00830_, _00826_);
  and (_00890_, _26637_, _00139_);
  and (_00891_, _26635_, _25475_);
  nor (_00892_, _00891_, _00890_);
  and (_00893_, _00892_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_00894_, _00892_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_00895_, _00894_, _00893_);
  nand (_00896_, _00895_, _00889_);
  or (_00897_, _00895_, _00889_);
  and (_00898_, _00897_, _26662_);
  and (_00899_, _00898_, _00896_);
  or (_00900_, _00899_, _00888_);
  or (_00901_, _00900_, _00884_);
  not (_00902_, _25475_);
  nand (_00903_, _26606_, _00902_);
  nand (_00904_, _00903_, _00339_);
  or (_00905_, _00904_, _00901_);
  and (_26870_[7], _00905_, _00850_);
  and (_00906_, _00847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00907_, _00847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_00908_, _00907_, _00906_);
  or (_00909_, _00908_, _00339_);
  and (_00910_, _00909_, _22731_);
  and (_00911_, _26570_, _26605_);
  and (_00912_, _26606_, _26631_);
  nor (_00913_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00914_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23275_);
  nor (_00915_, _00914_, _00913_);
  not (_00916_, _00915_);
  or (_00917_, _00916_, _23430_);
  and (_00918_, _00916_, _23430_);
  nor (_00919_, _00918_, _23391_);
  and (_00920_, _00919_, _00917_);
  nand (_00921_, _26377_, _23528_);
  nor (_00922_, _23975_, _23472_);
  not (_00923_, _00922_);
  nor (_00924_, _00923_, _23966_);
  nor (_00925_, _00924_, _23301_);
  and (_00926_, _00924_, _23301_);
  or (_00927_, _00926_, _23953_);
  nor (_00928_, _00927_, _00925_);
  and (_00929_, _23484_, _23301_);
  and (_00930_, _26457_, _23531_);
  and (_00931_, _23488_, _23460_);
  nor (_00932_, _23974_, _23296_);
  or (_00933_, _00932_, _00931_);
  or (_00934_, _00933_, _00930_);
  nor (_00935_, _00934_, _00929_);
  not (_00936_, _00935_);
  nor (_00937_, _00936_, _00928_);
  nand (_00938_, _00937_, _00921_);
  or (_00939_, _00938_, _00920_);
  and (_00940_, _00939_, _26574_);
  and (_00941_, _26665_, _23765_);
  and (_00942_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_00943_, _00942_, _00941_);
  or (_00944_, _00943_, _00940_);
  or (_00945_, _00944_, _00912_);
  or (_00946_, _00945_, _00911_);
  not (_00947_, _00339_);
  not (_00948_, _00894_);
  and (_00949_, _00948_, _00889_);
  or (_00950_, _00949_, _00893_);
  and (_00951_, _00950_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not (_00952_, _00951_);
  or (_00953_, _00950_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00954_, _00953_, _00952_);
  or (_00955_, _00954_, _00892_);
  nand (_00956_, _00954_, _00892_);
  and (_00957_, _00956_, _00955_);
  and (_00958_, _00957_, _26662_);
  or (_00959_, _00958_, _00947_);
  or (_00960_, _00959_, _00946_);
  and (_26870_[8], _00960_, _00910_);
  not (_00961_, _00892_);
  nor (_00962_, _00953_, _00961_);
  and (_00963_, _00951_, _00961_);
  nor (_00964_, _00963_, _00962_);
  nand (_00965_, _00964_, _23243_);
  or (_00966_, _00964_, _23243_);
  and (_00967_, _00966_, _00965_);
  and (_00968_, _00967_, _26662_);
  and (_00969_, _00393_, _26605_);
  not (_00970_, _26574_);
  nor (_00971_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_00973_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23243_);
  nor (_00974_, _00973_, _00971_);
  not (_00975_, _00974_);
  or (_00976_, _00975_, _00917_);
  and (_00977_, _00975_, _00917_);
  nor (_00978_, _00977_, _23391_);
  and (_00979_, _00978_, _00976_);
  not (_00980_, _00979_);
  and (_00981_, _26285_, _23528_);
  not (_00982_, _00981_);
  and (_00983_, _23484_, _23269_);
  nor (_00984_, _23323_, _23039_);
  and (_00986_, _00984_, _23964_);
  and (_00987_, _00986_, _23364_);
  and (_00988_, _23323_, _23039_);
  and (_00989_, _00988_, _23957_);
  and (_00990_, _00989_, _23456_);
  nor (_00991_, _00990_, _00987_);
  nor (_00992_, _00991_, _23305_);
  and (_00993_, _00991_, _23305_);
  or (_00995_, _00993_, _23953_);
  nor (_00996_, _00995_, _00992_);
  and (_00997_, _26410_, _23491_);
  not (_00998_, _00997_);
  and (_00999_, _00998_, _26424_);
  nor (_01000_, _00999_, _26458_);
  and (_01001_, _01000_, _23531_);
  and (_01002_, _23488_, _23115_);
  and (_01003_, _23506_, _23264_);
  or (_01004_, _01003_, _01002_);
  or (_01005_, _01004_, _01001_);
  or (_01006_, _01005_, _00996_);
  nor (_01007_, _01006_, _00983_);
  and (_01008_, _01007_, _00982_);
  and (_01009_, _01008_, _00980_);
  nor (_01010_, _01009_, _00970_);
  and (_01011_, _26665_, _23745_);
  and (_01012_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01013_, _26606_, _00157_);
  or (_01014_, _01013_, _01012_);
  or (_01015_, _01014_, _01011_);
  or (_01016_, _01015_, _01010_);
  or (_01017_, _01016_, _00969_);
  or (_01018_, _01017_, _00968_);
  and (_01019_, _01018_, _00339_);
  nor (_01020_, _00906_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01021_, _00906_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_01022_, _01021_, _01020_);
  nor (_01023_, _01022_, _00339_);
  or (_01024_, _01023_, _01019_);
  and (_26870_[9], _01024_, _22731_);
  nor (_01025_, _01021_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01026_, _01021_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01027_, _01026_, _01025_);
  or (_01028_, _01027_, _00339_);
  and (_01029_, _01028_, _22731_);
  and (_01030_, _00473_, _26605_);
  nor (_01031_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01032_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23215_);
  nor (_01033_, _01032_, _01031_);
  not (_01034_, _01033_);
  and (_01035_, _01034_, _00976_);
  not (_01036_, _01035_);
  or (_01037_, _01034_, _00976_);
  and (_01038_, _01037_, _23390_);
  and (_01039_, _01038_, _01036_);
  not (_01040_, _01039_);
  nor (_01041_, _26525_, _26522_);
  nor (_01042_, _01041_, _26526_);
  and (_01043_, _01042_, _23531_);
  and (_01044_, _23488_, _23959_);
  and (_01045_, _23484_, _23237_);
  or (_01046_, _01045_, _01044_);
  nor (_01047_, _01046_, _01043_);
  and (_01048_, _00990_, _23305_);
  and (_01049_, _00986_, _23269_);
  and (_01050_, _01049_, _23364_);
  nor (_01051_, _01050_, _01048_);
  nor (_01052_, _01051_, _23310_);
  and (_01053_, _01051_, _23310_);
  or (_01054_, _01053_, _23953_);
  nor (_01055_, _01054_, _01052_);
  and (_01056_, _23506_, _23232_);
  and (_01057_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  or (_01058_, _01057_, _01056_);
  nor (_01059_, _01058_, _01055_);
  and (_01060_, _01059_, _01047_);
  and (_01061_, _01060_, _01040_);
  nor (_01062_, _01061_, _00970_);
  and (_01063_, _26665_, _23724_);
  and (_01064_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_01065_, _01064_, _01063_);
  or (_01066_, _01065_, _01062_);
  or (_01067_, _01066_, _01030_);
  and (_01068_, _00962_, _23243_);
  and (_01069_, _00963_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_01071_, _01069_, _01068_);
  nand (_01072_, _01071_, _23215_);
  or (_01073_, _01071_, _23215_);
  and (_01074_, _01073_, _01072_);
  and (_01075_, _01074_, _26662_);
  or (_01076_, _01075_, _01067_);
  nand (_01077_, _26606_, _00224_);
  nand (_01078_, _01077_, _00339_);
  or (_01079_, _01078_, _01076_);
  and (_26870_[10], _01079_, _01029_);
  nor (_01080_, _01026_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01081_, _01026_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_01082_, _01081_, _01080_);
  or (_01083_, _01082_, _00339_);
  and (_01084_, _01083_, _22731_);
  and (_01085_, _00569_, _26605_);
  nor (_01086_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01087_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23177_);
  nor (_01088_, _01087_, _01086_);
  not (_01089_, _01088_);
  and (_01090_, _01089_, _01037_);
  not (_01091_, _01090_);
  or (_01092_, _01089_, _01037_);
  and (_01094_, _01092_, _23390_);
  and (_01095_, _01094_, _01091_);
  not (_01096_, _01095_);
  and (_01097_, _26529_, _26527_);
  not (_01098_, _01097_);
  and (_01099_, _01098_, _26530_);
  and (_01100_, _01099_, _23531_);
  not (_01101_, _01100_);
  and (_01102_, _01049_, _23237_);
  nor (_01103_, _01102_, _23456_);
  nor (_01104_, _23269_, _23237_);
  and (_01105_, _01104_, _00989_);
  nor (_01106_, _01105_, _23364_);
  or (_01107_, _01106_, _01103_);
  and (_01108_, _01107_, _23205_);
  nor (_01109_, _01107_, _23205_);
  nor (_01110_, _01109_, _01108_);
  and (_01111_, _01110_, _23514_);
  and (_01112_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor (_01113_, _23974_, _23199_);
  and (_01114_, _23484_, _23371_);
  or (_01115_, _01114_, _01113_);
  or (_01116_, _01115_, _23489_);
  nor (_01117_, _01116_, _01112_);
  not (_01118_, _01117_);
  nor (_01119_, _01118_, _01111_);
  and (_01120_, _01119_, _01101_);
  and (_01121_, _01120_, _01096_);
  nor (_01122_, _01121_, _00970_);
  and (_01123_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01124_, _26606_, _26810_);
  or (_01125_, _01124_, _01123_);
  or (_01126_, _01125_, _01122_);
  or (_01127_, _01126_, _01085_);
  and (_01128_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01129_, _01128_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01130_, _01129_, _00949_);
  nor (_01131_, _01130_, _00892_);
  or (_01132_, \oc8051_top_1.oc8051_memory_interface1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_01133_, _01132_, _00953_);
  and (_01134_, _01133_, _00892_);
  nor (_01135_, _01134_, _01131_);
  or (_01136_, _01135_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand (_01137_, _01135_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01138_, _01137_, _01136_);
  and (_01139_, _01138_, _26662_);
  or (_01140_, _01139_, _01127_);
  and (_01141_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01142_, \oc8051_top_1.oc8051_memory_interface1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_01143_, _01142_, _01141_);
  and (_01144_, \oc8051_top_1.oc8051_memory_interface1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01145_, _01144_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01146_, _01145_, _01143_);
  and (_01147_, _01146_, _01129_);
  and (_01148_, _01147_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_01149_, _01147_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_01150_, _01149_, _01148_);
  nand (_01151_, _01150_, _26665_);
  nand (_01152_, _01151_, _00339_);
  or (_01153_, _01152_, _01140_);
  and (_26870_[11], _01153_, _01084_);
  and (_01154_, _00654_, _26605_);
  nor (_01155_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01156_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23128_);
  nor (_01157_, _01156_, _01155_);
  not (_01158_, _01157_);
  and (_01159_, _01158_, _01092_);
  not (_01160_, _01159_);
  or (_01161_, _01158_, _01092_);
  and (_01162_, _01161_, _23390_);
  and (_01163_, _01162_, _01160_);
  not (_01164_, _01163_);
  and (_01165_, _26533_, _26531_);
  not (_01166_, _01165_);
  and (_01167_, _01166_, _26534_);
  and (_01168_, _01167_, _23531_);
  not (_01169_, _01168_);
  and (_01170_, _01105_, _23205_);
  and (_01171_, _01170_, _23456_);
  and (_01172_, _01102_, _23371_);
  and (_01173_, _01172_, _23364_);
  nor (_01174_, _01173_, _01171_);
  and (_01175_, _01174_, _23169_);
  nor (_01176_, _01174_, _23169_);
  nor (_01177_, _01176_, _01175_);
  and (_01178_, _01177_, _23514_);
  and (_01179_, _23506_, _23364_);
  nor (_01180_, _01179_, _23484_);
  or (_01181_, _01180_, _23169_);
  or (_01182_, _23974_, _23150_);
  or (_01183_, _01182_, _23364_);
  and (_01184_, _23488_, _23491_);
  and (_01185_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_01186_, _01185_, _01184_);
  and (_01187_, _01186_, _01183_);
  and (_01188_, _01187_, _01181_);
  not (_01189_, _01188_);
  nor (_01190_, _01189_, _01178_);
  and (_01191_, _01190_, _01169_);
  and (_01192_, _01191_, _01164_);
  nor (_01193_, _01192_, _00970_);
  and (_01194_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_01195_, _26606_, _00656_);
  or (_01197_, _01195_, _01194_);
  or (_01198_, _01197_, _01193_);
  or (_01199_, _01198_, _01154_);
  and (_01200_, _01129_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand (_01201_, _01200_, _00950_);
  nor (_01202_, _01201_, _00892_);
  nor (_01203_, _01133_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01204_, _01203_, _00892_);
  nor (_01205_, _01204_, _01202_);
  nand (_01206_, _01205_, _23128_);
  or (_01207_, _01205_, _23128_);
  and (_01208_, _01207_, _01206_);
  and (_01209_, _01208_, _26662_);
  or (_01210_, _01209_, _01199_);
  or (_01211_, _01148_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01212_, _01148_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_01213_, _01212_);
  and (_01214_, _01213_, _26665_);
  nand (_01215_, _01214_, _01211_);
  nand (_01216_, _01215_, _00339_);
  or (_01217_, _01216_, _01210_);
  not (_01218_, _25694_);
  and (_01219_, _00845_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_01220_, _01219_, _01218_);
  not (_01221_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand (_01222_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_01223_, _01222_, _01221_);
  nand (_01225_, _01223_, _01220_);
  nor (_01226_, _01225_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_01227_, _01225_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_01228_, _01227_, _01226_);
  or (_01229_, _01228_, _00339_);
  and (_01230_, _01229_, _22731_);
  and (_26870_[12], _01230_, _01217_);
  not (_01231_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_01232_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_01233_, _01225_, _01232_);
  nand (_01234_, _01233_, _01231_);
  or (_01236_, _01233_, _01231_);
  and (_01237_, _01236_, _01234_);
  or (_01238_, _01237_, _00339_);
  and (_01239_, _01238_, _22731_);
  and (_01240_, _00747_, _26605_);
  nor (_01241_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_01242_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23092_);
  nor (_01243_, _01242_, _01241_);
  not (_01244_, _01243_);
  and (_01245_, _01244_, _01161_);
  not (_01246_, _01245_);
  or (_01247_, _01244_, _01161_);
  and (_01248_, _01247_, _23390_);
  and (_01249_, _01248_, _01246_);
  not (_01250_, _01249_);
  and (_01251_, _26535_, _26513_);
  not (_01252_, _01251_);
  and (_01253_, _01252_, _26536_);
  and (_01255_, _01253_, _23531_);
  and (_01256_, _01172_, _23156_);
  nor (_01257_, _01256_, _23456_);
  and (_01258_, _23205_, _23169_);
  and (_01259_, _01258_, _01105_);
  nor (_01260_, _01259_, _23364_);
  or (_01261_, _01260_, _01257_);
  nor (_01262_, _01261_, _23122_);
  and (_01263_, _01261_, _23122_);
  nor (_01264_, _01263_, _01262_);
  nor (_01265_, _01264_, _23953_);
  and (_01266_, _23364_, _23122_);
  nor (_01267_, _23364_, _23457_);
  nor (_01268_, _01267_, _01266_);
  nor (_01269_, _01268_, _23974_);
  and (_01270_, _23484_, _23122_);
  and (_01271_, _23488_, _23264_);
  and (_01272_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or (_01273_, _01272_, _01271_);
  nor (_01274_, _01273_, _01270_);
  not (_01275_, _01274_);
  nor (_01276_, _01275_, _01269_);
  not (_01277_, _01276_);
  nor (_01278_, _01277_, _01265_);
  not (_01279_, _01278_);
  nor (_01280_, _01279_, _01255_);
  and (_01281_, _01280_, _01250_);
  nor (_01282_, _01281_, _00970_);
  and (_01283_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_01284_, _26606_, _00033_);
  or (_01285_, _01284_, _01283_);
  or (_01286_, _01285_, _01282_);
  or (_01287_, _01286_, _01240_);
  nor (_01288_, _00892_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_01289_, _01202_);
  nand (_01290_, _01203_, _23128_);
  and (_01291_, _01290_, _01289_);
  or (_01292_, _01291_, _01288_);
  nand (_01293_, _01292_, _23092_);
  or (_01294_, _01292_, _23092_);
  and (_01295_, _01294_, _01293_);
  and (_01296_, _01295_, _26662_);
  or (_01297_, _01296_, _01287_);
  and (_01298_, _01212_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_01299_, _01212_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_01300_, _01299_, _26665_);
  nor (_01302_, _01300_, _01298_);
  or (_01303_, _01302_, _00947_);
  or (_01304_, _01303_, _01297_);
  and (_26870_[13], _01304_, _01239_);
  or (_01305_, _01298_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01306_, _01298_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_01308_, _01306_);
  and (_01309_, _01308_, _26665_);
  and (_01310_, _01309_, _01305_);
  not (_01311_, _26605_);
  nor (_01312_, _00813_, _01311_);
  nor (_01313_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_01314_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _23057_);
  nor (_01315_, _01314_, _01313_);
  not (_01316_, _01315_);
  and (_01317_, _01316_, _01247_);
  not (_01318_, _01317_);
  or (_01319_, _01316_, _01247_);
  and (_01320_, _01319_, _23390_);
  and (_01321_, _01320_, _01318_);
  not (_01322_, _01321_);
  and (_01323_, _26537_, _26507_);
  not (_01324_, _01323_);
  and (_01325_, _01324_, _26538_);
  and (_01326_, _01325_, _23531_);
  and (_01327_, _01259_, _24022_);
  and (_01328_, _01256_, _23122_);
  and (_01329_, _01328_, _23364_);
  nor (_01330_, _01329_, _01327_);
  nor (_01331_, _01330_, _23086_);
  and (_01333_, _01330_, _23086_);
  nor (_01335_, _01333_, _01331_);
  and (_01337_, _01335_, _23514_);
  and (_01338_, _23484_, _23084_);
  nor (_01339_, _23364_, _23959_);
  not (_01340_, _01339_);
  and (_01341_, _23364_, _23086_);
  nor (_01342_, _01341_, _23974_);
  and (_01343_, _01342_, _01340_);
  and (_01344_, _23488_, _23232_);
  and (_01345_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or (_01346_, _01345_, _01344_);
  or (_01347_, _01346_, _01343_);
  nor (_01348_, _01347_, _01338_);
  not (_01349_, _01348_);
  nor (_01350_, _01349_, _01337_);
  not (_01351_, _01350_);
  nor (_01352_, _01351_, _01326_);
  and (_01353_, _01352_, _01322_);
  nor (_01354_, _01353_, _00970_);
  and (_01356_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_01357_, _26606_, _00070_);
  or (_01358_, _01357_, _01356_);
  or (_01359_, _01358_, _01354_);
  or (_01360_, _01359_, _01312_);
  or (_01361_, _01290_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_01362_, _01361_, _00961_);
  nand (_01363_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_01364_, _01363_, _01201_);
  or (_01365_, _01364_, _00892_);
  and (_01366_, _01365_, _01362_);
  nand (_01367_, _01366_, _23057_);
  or (_01369_, _01366_, _23057_);
  and (_01370_, _01369_, _01367_);
  and (_01371_, _01370_, _26662_);
  or (_01372_, _01371_, _01360_);
  or (_01373_, _01372_, _01310_);
  or (_01374_, _01373_, _00947_);
  not (_01375_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_01376_, _01236_, _01375_);
  or (_01377_, _01236_, _01375_);
  and (_01378_, _01377_, _01376_);
  or (_01380_, _01378_, _00339_);
  and (_01381_, _01380_, _22731_);
  and (_26870_[14], _01381_, _01374_);
  and (_01382_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _22731_);
  and (_01383_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  not (_01384_, _23615_);
  nor (_01385_, _23639_, _01384_);
  nor (_01386_, _23681_, _23660_);
  and (_01387_, _01386_, _01385_);
  nor (_01389_, _23765_, _23703_);
  not (_01390_, _23724_);
  nor (_01391_, _23745_, _01390_);
  and (_01393_, _01391_, _01389_);
  and (_01394_, _01393_, _01387_);
  not (_01395_, _23660_);
  and (_01396_, _01395_, _23615_);
  not (_01397_, _23681_);
  nor (_01398_, _01397_, _23639_);
  and (_01399_, _01398_, _01396_);
  nor (_01400_, _01399_, _01394_);
  and (_01401_, _23745_, _01390_);
  not (_01402_, _23765_);
  and (_01403_, _01402_, _23703_);
  and (_01405_, _01403_, _01401_);
  and (_01406_, _01405_, _01387_);
  and (_01408_, _23765_, _23703_);
  nor (_01410_, _23745_, _23724_);
  and (_01411_, _01410_, _01408_);
  and (_01412_, _01411_, _01387_);
  nor (_01413_, _01412_, _01406_);
  and (_01414_, _01413_, _01400_);
  and (_01415_, _01396_, _23639_);
  and (_01416_, _01415_, _23681_);
  and (_01417_, _23745_, _23724_);
  and (_01418_, _01417_, _01389_);
  and (_01419_, _01418_, _01416_);
  and (_01420_, _01415_, _01397_);
  not (_01422_, _01420_);
  and (_01424_, _01408_, _01401_);
  and (_01425_, _01410_, _23765_);
  nor (_01427_, _01425_, _01424_);
  nor (_01428_, _01427_, _01422_);
  nor (_01429_, _01428_, _01419_);
  and (_01430_, _01429_, _01414_);
  and (_01431_, _01385_, _23660_);
  and (_01432_, _01431_, _01397_);
  not (_01433_, _01432_);
  and (_01434_, _01417_, _01403_);
  nor (_01435_, _01434_, _01424_);
  nor (_01436_, _01435_, _01433_);
  not (_01437_, _01436_);
  and (_01438_, _01408_, _01391_);
  and (_01439_, _01438_, _01387_);
  nor (_01440_, _01402_, _23703_);
  and (_01441_, _01440_, _01401_);
  and (_01442_, _01441_, _01431_);
  nor (_01443_, _01442_, _01439_);
  and (_01444_, _01401_, _01389_);
  and (_01445_, _01444_, _01387_);
  and (_01446_, _01401_, _23765_);
  and (_01447_, _01446_, _01387_);
  nor (_01448_, _01447_, _01445_);
  and (_01449_, _01448_, _01443_);
  and (_01450_, _01449_, _01437_);
  and (_01451_, _01450_, _01430_);
  and (_01452_, _01391_, _23765_);
  not (_01453_, _01452_);
  and (_01454_, _01453_, _01435_);
  nor (_01455_, _01454_, _23615_);
  not (_01456_, _01455_);
  not (_01457_, _01415_);
  and (_01458_, _01403_, _01391_);
  nor (_01459_, _01458_, _01441_);
  nor (_01460_, _01459_, _01457_);
  and (_01461_, _01416_, _01410_);
  nor (_01462_, _01461_, _01460_);
  and (_01463_, _01440_, _01391_);
  nor (_01464_, _01458_, _01463_);
  nor (_01465_, _01464_, _01433_);
  not (_01466_, _01387_);
  and (_01467_, _01402_, _23745_);
  and (_01468_, _01467_, _23724_);
  nor (_01469_, _01463_, _01468_);
  nor (_01470_, _01469_, _01466_);
  nor (_01471_, _01470_, _01465_);
  and (_01472_, _01471_, _01462_);
  and (_01473_, _01472_, _01456_);
  and (_01474_, _01473_, _01451_);
  and (_01475_, _01431_, _23681_);
  and (_01476_, _01475_, _01444_);
  and (_01477_, _01458_, _01387_);
  nor (_01478_, _01477_, _01476_);
  nor (_01479_, _01438_, _01418_);
  nor (_01480_, _01479_, _01433_);
  not (_01481_, _01405_);
  nor (_01482_, _01432_, _01415_);
  nor (_01483_, _01482_, _01481_);
  nor (_01484_, _01483_, _01480_);
  and (_01485_, _01484_, _01478_);
  not (_01486_, _23703_);
  and (_01487_, _23765_, _23724_);
  and (_01488_, _01487_, _23745_);
  and (_01489_, _01488_, _01486_);
  and (_01490_, _01489_, _01416_);
  not (_01491_, _01490_);
  and (_01492_, _01438_, _01416_);
  and (_01493_, _01475_, _01405_);
  nor (_01494_, _01493_, _01492_);
  and (_01496_, _01494_, _01491_);
  not (_01497_, _01393_);
  nor (_01498_, _01432_, _01384_);
  nor (_01499_, _01498_, _01497_);
  not (_01501_, _01424_);
  and (_01502_, _01391_, _01486_);
  nor (_01503_, _01502_, _01438_);
  and (_01505_, _01503_, _01501_);
  and (_01506_, _23660_, _23639_);
  and (_01507_, _01506_, _23615_);
  not (_01508_, _01507_);
  nor (_01509_, _01508_, _01505_);
  nor (_01510_, _01509_, _01499_);
  and (_01511_, _01510_, _01496_);
  and (_01512_, _01511_, _01485_);
  and (_01513_, _01488_, _23703_);
  and (_01514_, _01513_, _01416_);
  nor (_01515_, _01514_, _01444_);
  nor (_01516_, _01515_, _01482_);
  not (_01517_, _01516_);
  and (_01518_, _01434_, _01416_);
  and (_01519_, _01438_, _01420_);
  nor (_01520_, _01519_, _01518_);
  and (_01521_, _01410_, _01402_);
  and (_01522_, _01521_, _01432_);
  not (_01523_, _01522_);
  and (_01524_, _01410_, _01403_);
  and (_01525_, _01524_, _01387_);
  and (_01526_, _01440_, _01410_);
  and (_01527_, _01526_, _01387_);
  or (_01528_, _01527_, _01525_);
  or (_01529_, _01424_, _01393_);
  and (_01530_, _01529_, _01416_);
  nor (_01531_, _01530_, _01528_);
  and (_01532_, _01531_, _01523_);
  and (_01533_, _01532_, _01520_);
  and (_01534_, _01533_, _01517_);
  and (_01535_, _01534_, _01512_);
  and (_01536_, _01535_, _01474_);
  and (_01537_, _01475_, _01441_);
  or (_01538_, _01506_, _01384_);
  and (_01539_, _01538_, _01438_);
  or (_01540_, _01539_, _01412_);
  nor (_01541_, _01540_, _01537_);
  and (_01542_, _01541_, _01494_);
  and (_01543_, _01542_, _01478_);
  nand (_01544_, _01543_, _01533_);
  or (_01545_, _01544_, _01536_);
  and (_01546_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_01547_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_01548_, _01547_, _01546_);
  and (_01549_, _01548_, _01545_);
  nor (_01550_, _01548_, _01545_);
  nor (_01551_, _01550_, _01549_);
  or (_01552_, _01551_, _24471_);
  or (_01553_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_01554_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_01555_, _01554_, _01553_);
  and (_01556_, _01555_, _01552_);
  or (_26871_[0], _01556_, _01383_);
  not (_01557_, _01536_);
  and (_01558_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_01559_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_01560_, _01559_, _01558_);
  and (_01561_, _01560_, _01546_);
  nor (_01562_, _01560_, _01546_);
  nor (_01563_, _01562_, _01561_);
  nand (_01564_, _01563_, _01557_);
  or (_01565_, _01563_, _01557_);
  and (_01566_, _01565_, _01564_);
  nand (_01567_, _01566_, _01549_);
  or (_01568_, _01566_, _01549_);
  and (_01569_, _01568_, _01567_);
  or (_01570_, _01569_, _24471_);
  or (_01571_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01572_, _01571_, _01554_);
  and (_01573_, _01572_, _01570_);
  and (_01574_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_26871_[1], _01574_, _01573_);
  and (_01575_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nand (_01576_, _01567_, _01564_);
  nor (_01577_, _01561_, _01558_);
  not (_01578_, _01577_);
  and (_01579_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_01580_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_01581_, _01580_, _01579_);
  and (_01582_, _01581_, _01578_);
  nor (_01583_, _01581_, _01578_);
  nor (_01584_, _01583_, _01582_);
  and (_01585_, _01584_, _01576_);
  nor (_01586_, _01584_, _01576_);
  nor (_01587_, _01586_, _01585_);
  or (_01588_, _01587_, _24471_);
  or (_01589_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_01590_, _01589_, _01554_);
  and (_01591_, _01590_, _01588_);
  or (_26871_[2], _01591_, _01575_);
  nor (_01592_, _01582_, _01579_);
  nor (_01593_, _01592_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_01594_, _01592_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_01595_, _01594_, _01593_);
  and (_01596_, _01595_, _01585_);
  nor (_01597_, _01595_, _01585_);
  nor (_01598_, _01597_, _01596_);
  or (_01599_, _01598_, _24471_);
  or (_01601_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01602_, _01601_, _01554_);
  and (_01603_, _01602_, _01599_);
  and (_01605_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_26871_[3], _01605_, _01603_);
  and (_01607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_01608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_01609_, _01608_, _01607_);
  nand (_01610_, _01609_, _01593_);
  or (_01611_, _01609_, _01593_);
  and (_01612_, _01611_, _01610_);
  and (_01613_, _01612_, _01596_);
  nor (_01614_, _01612_, _01596_);
  nor (_01615_, _01614_, _01613_);
  or (_01616_, _01615_, _24471_);
  or (_01617_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01618_, _01617_, _01554_);
  and (_01619_, _01618_, _01616_);
  and (_01620_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_26871_[4], _01620_, _01619_);
  not (_01621_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _01621_);
  and (_01623_, _01622_, _22731_);
  nand (_01624_, _01608_, _01592_);
  and (_01625_, _01624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not (_01626_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_01627_, _01608_, _01626_);
  and (_01628_, _01627_, _01592_);
  or (_01629_, _01628_, _01625_);
  or (_01630_, _01629_, _01613_);
  and (_01631_, _01629_, _01612_);
  and (_01632_, _01631_, _01596_);
  nor (_01633_, _01632_, _24471_);
  and (_01634_, _01633_, _01630_);
  nor (_01635_, _24470_, _23090_);
  or (_01636_, _01635_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01637_, _01636_, _01634_);
  and (_26871_[5], _01637_, _01623_);
  not (_01638_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_01639_, _01628_, _01638_);
  and (_01640_, _01627_, _01638_);
  and (_01641_, _01640_, _01592_);
  nor (_01642_, _01641_, _01639_);
  not (_01643_, _01642_);
  and (_01644_, _01643_, _01632_);
  nor (_01645_, _01643_, _01632_);
  nor (_01646_, _01645_, _01644_);
  or (_01647_, _01646_, _24471_);
  or (_01648_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01649_, _01648_, _01554_);
  and (_01650_, _01649_, _01647_);
  and (_01651_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_26871_[6], _01651_, _01650_);
  and (_01652_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_01653_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_01654_, _01640_, _01653_);
  and (_01655_, _01654_, _01592_);
  nor (_01656_, _01641_, _01653_);
  nor (_01657_, _01656_, _01655_);
  not (_01658_, _01657_);
  and (_01659_, _01658_, _01644_);
  nor (_01660_, _01658_, _01644_);
  nor (_01661_, _01660_, _01659_);
  or (_01663_, _01661_, _24471_);
  or (_01664_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01665_, _01664_, _01554_);
  and (_01666_, _01665_, _01663_);
  or (_26871_[7], _01666_, _01652_);
  not (_01667_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_01668_, _01655_, _01667_);
  and (_01669_, _01654_, _01667_);
  and (_01670_, _01669_, _01592_);
  or (_01671_, _01670_, _01668_);
  and (_01672_, _01671_, _01659_);
  nor (_01673_, _01671_, _01659_);
  nor (_01674_, _01673_, _01672_);
  or (_01675_, _01674_, _24471_);
  or (_01676_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01677_, _01676_, _01554_);
  and (_01678_, _01677_, _01675_);
  and (_01679_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_26871_[8], _01679_, _01678_);
  not (_01680_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_01681_, _01669_, _01680_);
  and (_01682_, _01681_, _01592_);
  nor (_01683_, _01670_, _01680_);
  nor (_01684_, _01683_, _01682_);
  not (_01685_, _01684_);
  and (_01686_, _01685_, _01672_);
  or (_01687_, _01685_, _01672_);
  nand (_01689_, _01687_, _24470_);
  nor (_01690_, _01689_, _01686_);
  nor (_01691_, _24470_, _23243_);
  or (_01692_, _01691_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01693_, _01692_, _01690_);
  or (_01694_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _01621_);
  and (_01695_, _01694_, _22731_);
  and (_26871_[9], _01695_, _01693_);
  not (_01696_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01697_, _01682_, _01696_);
  and (_01699_, _01681_, _01696_);
  and (_01700_, _01699_, _01592_);
  nor (_01701_, _01700_, _01697_);
  not (_01702_, _01701_);
  and (_01703_, _01702_, _01686_);
  nor (_01704_, _01702_, _01686_);
  nor (_01705_, _01704_, _01703_);
  or (_01706_, _01705_, _24471_);
  or (_01707_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01708_, _01707_, _01554_);
  and (_01709_, _01708_, _01706_);
  and (_01710_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_26871_[10], _01710_, _01709_);
  and (_01711_, _01699_, _01221_);
  and (_01712_, _01711_, _01592_);
  nor (_01713_, _01700_, _01221_);
  nor (_01714_, _01713_, _01712_);
  not (_01715_, _01714_);
  and (_01716_, _01715_, _01703_);
  or (_01717_, _01715_, _01703_);
  nand (_01718_, _01717_, _24470_);
  nor (_01719_, _01718_, _01716_);
  nor (_01720_, _24470_, _23177_);
  or (_01721_, _01720_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01722_, _01721_, _01719_);
  or (_01723_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _01621_);
  and (_01724_, _01723_, _22731_);
  and (_26871_[11], _01724_, _01722_);
  nor (_01725_, _01712_, _01232_);
  and (_01726_, _01711_, _01232_);
  and (_01727_, _01726_, _01592_);
  or (_01728_, _01727_, _01725_);
  and (_01730_, _01728_, _01716_);
  nor (_01731_, _01728_, _01716_);
  nor (_01732_, _01731_, _01730_);
  or (_01733_, _01732_, _24471_);
  or (_01734_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01735_, _01734_, _01554_);
  and (_01736_, _01735_, _01733_);
  and (_01737_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_26871_[12], _01737_, _01736_);
  and (_01738_, _01727_, _01231_);
  nor (_01739_, _01727_, _01231_);
  nor (_01740_, _01739_, _01738_);
  not (_01741_, _01740_);
  and (_01742_, _01741_, _01730_);
  nor (_01743_, _01741_, _01730_);
  nor (_01744_, _01743_, _01742_);
  or (_01745_, _01744_, _24471_);
  or (_01746_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01747_, _01746_, _01554_);
  and (_01748_, _01747_, _01745_);
  and (_01749_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_26871_[13], _01749_, _01748_);
  nor (_01750_, _01738_, _01375_);
  and (_01751_, _01738_, _01375_);
  nor (_01752_, _01751_, _01750_);
  not (_01753_, _01752_);
  and (_01754_, _01753_, _01742_);
  nor (_01755_, _01753_, _01742_);
  nor (_01756_, _01755_, _01754_);
  or (_01757_, _01756_, _24471_);
  or (_01758_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01759_, _01758_, _01554_);
  and (_01760_, _01759_, _01757_);
  and (_01761_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_26871_[14], _01761_, _01760_);
  and (_01762_, _25648_, _24051_);
  and (_01763_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  or (_22617_, _01763_, _01762_);
  and (_01764_, _26020_, _24134_);
  and (_01765_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  or (_22618_, _01765_, _01764_);
  nor (_01766_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor (_01767_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_01768_, _01767_, _01766_);
  not (_01769_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor (_01770_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_01771_, _01770_, _01769_);
  and (_01772_, _01771_, _01768_);
  and (_01773_, _01772_, _25010_);
  and (_01774_, _01773_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_01775_, _01774_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_26875_[0], _01775_, _22731_);
  and (_01776_, _01773_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_01777_, _01776_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_26875_[1], _01777_, _22731_);
  and (_01778_, _01773_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or (_01779_, _01778_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_26875_[2], _01779_, _22731_);
  and (_01780_, _01772_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_01781_, _01780_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_26875_[3], _01781_, _22731_);
  and (_01782_, _01773_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_01783_, _01782_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_26875_[4], _01783_, _22731_);
  and (_01784_, _01773_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_01785_, _01784_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_26875_[5], _01785_, _22731_);
  and (_01786_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22731_);
  and (_01787_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _22731_);
  and (_01788_, _01787_, _01773_);
  or (_26875_[6], _01788_, _01786_);
  and (_01789_, _01545_, _22737_);
  nand (_01790_, _01789_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_01791_, _01789_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_01792_, _01791_, _01554_);
  and (_26876_[0], _01792_, _01790_);
  and (_01793_, _01545_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_01794_, _01536_, _23599_);
  nand (_01795_, _01536_, _23599_);
  and (_01796_, _01795_, _01794_);
  nand (_01797_, _01796_, _01793_);
  or (_01798_, _01796_, _01793_);
  and (_01800_, _01798_, _01797_);
  or (_01801_, _01800_, _25454_);
  or (_01802_, _22737_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01803_, _01802_, _01554_);
  and (_26876_[1], _01803_, _01801_);
  and (_01804_, _26020_, _24051_);
  and (_01805_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  or (_22619_, _01805_, _01804_);
  and (_01806_, _26020_, _24089_);
  and (_01807_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  or (_22621_, _01807_, _01806_);
  and (_01808_, _24320_, _23583_);
  and (_01809_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_22622_, _01809_, _01808_);
  and (_01810_, _24301_, _24095_);
  and (_01811_, _01810_, _24219_);
  not (_01812_, _01810_);
  and (_01813_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  or (_22623_, _01813_, _01811_);
  and (_01814_, _25497_, _24174_);
  nor (_01815_, _01814_, rst);
  and (_01816_, _25607_, _24174_);
  not (_01817_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  and (_01818_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor (_01819_, _01818_, _01817_);
  and (_01820_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_01821_, _01820_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_01822_, _01821_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_01823_, _01822_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_01824_, _01823_, _01818_);
  and (_01825_, _01824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_01826_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_01827_, _01826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01828_, _01827_, _01819_);
  and (_01829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_01830_, _01829_, _01828_);
  nor (_01831_, _01830_, _01816_);
  and (_22624_, _01831_, _01815_);
  and (_01832_, _24476_, _24372_);
  and (_01833_, _01832_, _24051_);
  not (_01834_, _01832_);
  and (_01835_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_22625_, _01835_, _01833_);
  not (_01836_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  and (_01837_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_01838_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_01839_, _01838_, _01837_);
  and (_26879_[0], _01839_, _22731_);
  and (_01840_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_01841_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01842_, _01841_, _01840_);
  and (_26879_[1], _01842_, _22731_);
  and (_01843_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_01844_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01845_, _01844_, _01843_);
  and (_26879_[2], _01845_, _22731_);
  and (_01846_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_01847_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01848_, _01847_, _01846_);
  and (_26879_[3], _01848_, _22731_);
  and (_01849_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_01850_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01851_, _01850_, _01849_);
  and (_26879_[4], _01851_, _22731_);
  and (_01852_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_01853_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01854_, _01853_, _01852_);
  and (_26879_[5], _01854_, _22731_);
  and (_01855_, _01836_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_01856_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_01857_, _01856_, _01855_);
  and (_26879_[6], _01857_, _22731_);
  not (_01858_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_01859_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor (_01860_, _01859_, _01858_);
  and (_01861_, _01859_, _01858_);
  nor (_01862_, _01861_, _01860_);
  and (_26882_[0], _01862_, _22731_);
  nor (_01863_, _01860_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_01864_, _01860_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_01865_, _01864_, _01863_);
  nor (_26882_[1], _01865_, rst);
  and (_01866_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_01867_, _01866_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01868_, _01866_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_01869_, _01868_, _01867_);
  or (_01870_, _01869_, _01859_);
  and (_26882_[2], _01870_, _22731_);
  and (_01871_, _01832_, _24089_);
  and (_01872_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_27066_, _01872_, _01871_);
  and (_01873_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_01874_, _25694_, _25696_);
  or (_01875_, _01874_, _01873_);
  and (_26884_[0], _01875_, _22731_);
  and (_01876_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_01877_, _25694_, _25700_);
  or (_01878_, _01877_, _01876_);
  and (_26884_[1], _01878_, _22731_);
  and (_01879_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_01880_, _25694_, _25705_);
  or (_01881_, _01880_, _01879_);
  and (_26884_[2], _01881_, _22731_);
  and (_01882_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_01883_, _25694_, _25711_);
  or (_01884_, _01883_, _01882_);
  and (_26884_[3], _01884_, _22731_);
  and (_01885_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_01886_, _25694_, _25715_);
  or (_01887_, _01886_, _01885_);
  and (_26884_[4], _01887_, _22731_);
  and (_01888_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_01889_, _25694_, _25720_);
  or (_01890_, _01889_, _01888_);
  and (_26884_[5], _01890_, _22731_);
  and (_01891_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_01892_, _25694_, _25724_);
  or (_01893_, _01892_, _01891_);
  and (_26884_[6], _01893_, _22731_);
  and (_01894_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_01895_, _25694_, _25729_);
  or (_01896_, _01895_, _01894_);
  and (_26884_[7], _01896_, _22731_);
  and (_01897_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_01898_, _25694_, _25735_);
  or (_01899_, _01898_, _01897_);
  and (_26884_[8], _01899_, _22731_);
  and (_01900_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_01901_, _25694_, _25739_);
  or (_01902_, _01901_, _01900_);
  and (_26884_[9], _01902_, _22731_);
  and (_01903_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_01904_, _25694_, _25744_);
  or (_01905_, _01904_, _01903_);
  and (_26884_[10], _01905_, _22731_);
  and (_01906_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_01907_, _25694_, _25750_);
  or (_01908_, _01907_, _01906_);
  and (_26884_[11], _01908_, _22731_);
  and (_01909_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_01910_, _25694_, _25754_);
  or (_01911_, _01910_, _01909_);
  and (_26884_[12], _01911_, _22731_);
  and (_01912_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_01913_, _25694_, _25758_);
  or (_01914_, _01913_, _01912_);
  and (_26884_[13], _01914_, _22731_);
  and (_01915_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_01916_, _25694_, _25763_);
  or (_01917_, _01916_, _01915_);
  and (_26884_[14], _01917_, _22731_);
  and (_01918_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_01919_, _25694_, _25767_);
  or (_01920_, _01919_, _01918_);
  and (_26884_[15], _01920_, _22731_);
  and (_01921_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_01922_, _25694_, _25771_);
  or (_01923_, _01922_, _01921_);
  and (_26884_[16], _01923_, _22731_);
  and (_01924_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_01926_, _25694_, _25776_);
  or (_01927_, _01926_, _01924_);
  and (_26884_[17], _01927_, _22731_);
  and (_01928_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_01929_, _25694_, _25780_);
  or (_01930_, _01929_, _01928_);
  and (_26884_[18], _01930_, _22731_);
  and (_01931_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_01932_, _25694_, _25784_);
  or (_01933_, _01932_, _01931_);
  and (_26884_[19], _01933_, _22731_);
  and (_01934_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_01935_, _25694_, _25788_);
  or (_01936_, _01935_, _01934_);
  and (_26884_[20], _01936_, _22731_);
  and (_01937_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_01938_, _25694_, _25792_);
  or (_01939_, _01938_, _01937_);
  and (_26884_[21], _01939_, _22731_);
  and (_01940_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_01941_, _25694_, _25796_);
  or (_01942_, _01941_, _01940_);
  and (_26884_[22], _01942_, _22731_);
  and (_01943_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_01944_, _25694_, _25800_);
  or (_01945_, _01944_, _01943_);
  and (_26884_[23], _01945_, _22731_);
  and (_01946_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_01947_, _25694_, _25804_);
  or (_01948_, _01947_, _01946_);
  and (_26884_[24], _01948_, _22731_);
  and (_01949_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_01950_, _25694_, _25808_);
  or (_01951_, _01950_, _01949_);
  and (_26884_[25], _01951_, _22731_);
  and (_01952_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_01953_, _25694_, _25812_);
  or (_01954_, _01953_, _01952_);
  and (_26884_[26], _01954_, _22731_);
  and (_01955_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_01956_, _25694_, _25816_);
  or (_01957_, _01956_, _01955_);
  and (_26884_[27], _01957_, _22731_);
  and (_01958_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_01959_, _25694_, _25820_);
  or (_01960_, _01959_, _01958_);
  and (_26884_[28], _01960_, _22731_);
  and (_01961_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_01962_, _25694_, _25825_);
  or (_01963_, _01962_, _01961_);
  and (_26884_[29], _01963_, _22731_);
  and (_01964_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_01965_, _25694_, _25829_);
  or (_01966_, _01965_, _01964_);
  and (_26884_[30], _01966_, _22731_);
  and (_01967_, _24257_, _23780_);
  and (_01968_, _23926_, _23780_);
  or (_01969_, _26673_, _24244_);
  or (_01970_, _01969_, _01968_);
  or (_01971_, _01970_, _01967_);
  or (_01972_, _01971_, _26749_);
  and (_01973_, _23844_, _23687_);
  or (_01974_, _23912_, _23790_);
  or (_01975_, _01974_, _01973_);
  or (_01976_, _23836_, _23773_);
  or (_01977_, _01976_, _24267_);
  and (_01978_, _23827_, _23687_);
  and (_01979_, _26693_, _23687_);
  or (_01980_, _01979_, _23898_);
  or (_01981_, _01980_, _01978_);
  or (_01982_, _01981_, _01977_);
  or (_01983_, _01982_, _01975_);
  or (_01984_, _24269_, _23916_);
  and (_01985_, _23911_, _23816_);
  and (_01986_, _23814_, _23789_);
  and (_01987_, _23825_, _23788_);
  or (_01988_, _01987_, _01986_);
  or (_01989_, _01988_, _01985_);
  and (_01990_, _23781_, _23786_);
  and (_01991_, _01990_, _23707_);
  and (_01992_, _01991_, _23803_);
  and (_01993_, _23911_, _23814_);
  or (_01994_, _01993_, _23830_);
  or (_01995_, _01994_, _01992_);
  or (_01996_, _01995_, _01989_);
  or (_01997_, _01996_, _01984_);
  or (_01998_, _01997_, _01983_);
  or (_01999_, _01998_, _01972_);
  and (_02000_, _01999_, _22737_);
  and (_02001_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_02002_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_02003_, _26601_, _02002_);
  nor (_02004_, _24246_, _23708_);
  and (_02005_, _23816_, _23788_);
  nor (_02006_, _02005_, _24246_);
  nand (_02007_, _23788_, _23779_);
  and (_02008_, _02007_, _02006_);
  nor (_02009_, _02008_, _02004_);
  and (_02010_, _02009_, _02003_);
  or (_02011_, _02010_, _26681_);
  or (_02012_, _02011_, _02001_);
  or (_02013_, _02012_, _02000_);
  and (_26849_[1], _02013_, _22731_);
  and (_02014_, _23830_, _23791_);
  and (_02015_, _26594_, _23707_);
  or (_02016_, _02015_, _24251_);
  or (_02017_, _02016_, _02014_);
  and (_02018_, _23803_, _23789_);
  and (_02019_, _01991_, _23814_);
  and (_02020_, _01991_, _23824_);
  and (_02021_, _26593_, _23707_);
  or (_02022_, _02021_, _02020_);
  or (_02023_, _02022_, _02019_);
  or (_02024_, _02023_, _02018_);
  and (_02025_, _23926_, _23687_);
  or (_02026_, _02025_, _23910_);
  or (_02027_, _24273_, _24258_);
  or (_02028_, _02027_, _02026_);
  or (_02029_, _02028_, _02024_);
  or (_02031_, _01984_, _24250_);
  or (_02032_, _02031_, _02029_);
  or (_02033_, _02032_, _02017_);
  or (_02034_, _02033_, _01983_);
  and (_02035_, _02034_, _22737_);
  and (_02036_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02037_, _02036_, _02011_);
  or (_02038_, _02037_, _02035_);
  and (_26849_[0], _02038_, _22731_);
  and (_02039_, _24097_, _23944_);
  and (_02040_, _02039_, _24159_);
  not (_02041_, _02040_);
  and (_02043_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_02044_, _02040_, _23996_);
  or (_22626_, _02044_, _02043_);
  nand (_26842_[0], _02009_, _23855_);
  and (_02045_, _24301_, _24159_);
  and (_02046_, _02045_, _23583_);
  not (_02047_, _02045_);
  and (_02048_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_27232_, _02048_, _02046_);
  nor (_02049_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_02050_, _02049_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  not (_02051_, _02050_);
  or (_02053_, _02051_, _26570_);
  or (_02054_, _02050_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_02055_, _02054_, _22731_);
  and (_26888_[0], _02055_, _02053_);
  or (_02056_, _02051_, _00393_);
  or (_02057_, _02050_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_02058_, _02057_, _22731_);
  and (_26888_[1], _02058_, _02056_);
  or (_02059_, _02051_, _00473_);
  or (_02060_, _02050_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_02061_, _02060_, _22731_);
  and (_26888_[2], _02061_, _02059_);
  or (_02062_, _02051_, _00569_);
  or (_02063_, _02050_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_02064_, _02063_, _22731_);
  and (_26888_[3], _02064_, _02062_);
  and (_02065_, _24236_, _24006_);
  and (_02066_, _02065_, _24219_);
  not (_02067_, _02065_);
  and (_02068_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  or (_22627_, _02068_, _02066_);
  and (_02069_, _02045_, _24089_);
  and (_02070_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_22628_, _02070_, _02069_);
  and (_02071_, _24553_, _24174_);
  or (_02072_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_02073_, _02072_, _22731_);
  not (_02074_, _02071_);
  or (_02075_, _02074_, _23880_);
  and (_22629_, _02075_, _02073_);
  and (_02076_, _01832_, _24134_);
  and (_02077_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_22630_, _02077_, _02076_);
  nor (_02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_02079_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _22731_);
  and (_02082_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_22631_, _02082_, _02079_);
  and (_02083_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_02084_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_22632_, _02084_, _02083_);
  and (_02085_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_02086_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_22633_, _02086_, _02085_);
  and (_02087_, _01832_, _23996_);
  and (_02088_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_22634_, _02088_, _02087_);
  and (_02089_, _02045_, _24051_);
  and (_02090_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_22635_, _02090_, _02089_);
  and (_02091_, _25648_, _23548_);
  and (_02092_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  or (_22636_, _02092_, _02091_);
  and (_02093_, _24476_, _24146_);
  and (_02094_, _02093_, _23583_);
  not (_02095_, _02093_);
  and (_02096_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_27037_, _02096_, _02094_);
  and (_02097_, _02093_, _24051_);
  and (_02098_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_22637_, _02098_, _02097_);
  and (_02100_, _02093_, _24089_);
  and (_02101_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_22638_, _02101_, _02100_);
  and (_22639_, _01786_, _24747_);
  and (_02102_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_02103_, _02102_, _24841_);
  and (_22640_, _02103_, _22731_);
  or (_02104_, _24844_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_02105_, _02104_, _22731_);
  not (_02106_, _24763_);
  or (_02107_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_02108_, _02107_, _02106_);
  nor (_02109_, _24915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or (_02110_, _02109_, _24919_);
  and (_02111_, _02110_, _02108_);
  or (_02112_, _02111_, _24757_);
  and (_02113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _24750_);
  nand (_02114_, _24777_, _24763_);
  nand (_02115_, _02114_, _24758_);
  nand (_02116_, _02115_, _02113_);
  nand (_02117_, _02116_, _02112_);
  and (_02118_, _02117_, _24809_);
  and (_02119_, _24805_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  not (_02120_, _24802_);
  and (_02121_, _02107_, _02120_);
  or (_02122_, _24931_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_02123_, _24930_, _24802_);
  and (_02124_, _02123_, _02122_);
  or (_02125_, _02124_, _02121_);
  and (_02126_, _02125_, _24797_);
  and (_02127_, _24802_, _24790_);
  or (_02129_, _02127_, _24795_);
  and (_02130_, _02129_, _02113_);
  or (_02131_, _02130_, _02126_);
  and (_02132_, _02131_, _24806_);
  or (_02133_, _02132_, _02119_);
  and (_02134_, _02133_, _24781_);
  or (_02135_, _02134_, _02118_);
  or (_02136_, _02135_, _24747_);
  and (_22641_, _02136_, _02105_);
  and (_02137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_02138_, _02137_, _24777_);
  or (_02139_, _24848_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_02140_, _02139_, _24846_);
  or (_02141_, _02140_, _02138_);
  and (_02142_, _02141_, _24763_);
  or (_02143_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _24750_);
  and (_02144_, _02143_, _02106_);
  or (_02145_, _02144_, _02142_);
  and (_02146_, _02145_, _25006_);
  and (_02147_, _02143_, _02120_);
  or (_02148_, _24870_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_02149_, _24869_, _24802_);
  and (_02150_, _02149_, _02148_);
  or (_02152_, _02150_, _02147_);
  and (_02153_, _02152_, _24943_);
  or (_02154_, _02153_, _02146_);
  and (_02155_, _02154_, _24844_);
  and (_02156_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_02157_, _02156_, _24805_);
  and (_02158_, _02157_, _24781_);
  nand (_02159_, _24757_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_02160_, _02159_, _24781_);
  or (_02161_, _02160_, _24747_);
  or (_02162_, _02161_, _02158_);
  and (_02163_, _02162_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or (_02164_, _02163_, _02155_);
  and (_22642_, _02164_, _22731_);
  and (_02166_, _24621_, _24607_);
  nand (_02167_, _02166_, _23504_);
  or (_02168_, _02166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_02169_, _02168_, _24630_);
  and (_02170_, _02169_, _02167_);
  nor (_02171_, _24630_, _24043_);
  or (_02172_, _02171_, _02170_);
  and (_22643_, _02172_, _22731_);
  and (_02173_, _24636_, _24544_);
  and (_02174_, _02173_, _23504_);
  nor (_02175_, _02173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_02176_, _02175_, _02174_);
  nand (_02177_, _02176_, _24557_);
  nand (_02178_, _24554_, _24082_);
  and (_02179_, _02178_, _22731_);
  and (_22644_, _02179_, _02177_);
  and (_02180_, _24451_, _23996_);
  and (_02181_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_22645_, _02181_, _02180_);
  and (_02182_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_02183_, _02040_, _23887_);
  or (_27028_, _02183_, _02182_);
  and (_02184_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_02185_, _02040_, _23583_);
  or (_27029_, _02185_, _02184_);
  and (_02186_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_02187_, _02040_, _23548_);
  or (_22646_, _02187_, _02186_);
  and (_02188_, _01832_, _24219_);
  and (_02189_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_22647_, _02189_, _02188_);
  and (_02190_, _02093_, _23996_);
  and (_02191_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_22648_, _02191_, _02190_);
  nand (_02192_, _01816_, _23989_);
  not (_02193_, _01814_);
  or (_02194_, _02193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_02195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_02196_, _02195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_02197_, _02195_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_02198_, _02197_, _02196_);
  not (_02199_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_02200_, _02199_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_02201_, t0_i);
  and (_02202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _02201_);
  and (_02203_, _02202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff );
  or (_02204_, _02203_, _02200_);
  and (_02205_, _02204_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_02206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_02207_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_02208_, _02207_, _02206_);
  and (_02209_, _02208_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_02210_, _02209_, _02205_);
  and (_02211_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_02212_, _02211_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_02213_, _02212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_02214_, _02213_, _02198_);
  nand (_02215_, _02196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_02216_, _02212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nand (_02217_, _02216_, _02215_);
  and (_02218_, _02217_, _02214_);
  nor (_02219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_02220_, _02219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_02221_, _02216_);
  and (_02222_, _02221_, _01829_);
  or (_02223_, _02222_, _02220_);
  and (_02224_, _02223_, _02213_);
  or (_02225_, _02224_, _02218_);
  or (_02226_, _02225_, _01814_);
  and (_02227_, _02226_, _02194_);
  or (_02228_, _02227_, _01816_);
  and (_02229_, _02228_, _22731_);
  and (_22649_, _02229_, _02192_);
  and (_02230_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_02231_, _02040_, _24051_);
  or (_22650_, _02231_, _02230_);
  and (_02232_, _24476_, _24140_);
  and (_02233_, _02232_, _24051_);
  not (_02234_, _02232_);
  and (_02235_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  or (_22651_, _02235_, _02233_);
  not (_02236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_02237_, _02236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  not (_02238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_02239_, t1_i);
  and (_02240_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _02239_);
  nor (_02241_, _02240_, _02238_);
  not (_02242_, _02241_);
  not (_02243_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_02244_, _02243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  nor (_02245_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_02246_, _02245_);
  and (_02247_, _02246_, _02244_);
  and (_02248_, _02247_, _02242_);
  not (_02249_, _02248_);
  and (_02250_, _02249_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and (_02251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_02252_, _02251_, _02248_);
  and (_02253_, _02252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_02254_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not (_02255_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_02256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_02257_, _02256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand (_02258_, _02257_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_02259_, _02258_, _02255_);
  and (_02260_, _02259_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_02262_, _02260_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_02263_, _02262_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_02264_, _02263_, _02254_);
  and (_02265_, _02264_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_02266_, _02265_, _02253_);
  and (_02267_, _02266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_02268_, _02267_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_02269_, _02268_, _02250_);
  and (_02270_, _02269_, _02237_);
  nor (_02271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_02272_, _02259_, _02254_);
  and (_02273_, _02272_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_02274_, _02273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_02275_, _02274_, _02251_);
  and (_02276_, _02275_, _02248_);
  and (_02277_, _02276_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_02278_, _02277_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_02279_, _02278_, _02250_);
  and (_02280_, _02279_, _02271_);
  and (_02281_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_02282_, _02281_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_02283_, _02236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_02284_, _02262_, _02248_);
  and (_02285_, _02284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or (_02286_, _02285_, _02250_);
  and (_02287_, _02286_, _02283_);
  or (_02288_, _02287_, _02282_);
  or (_02289_, _02288_, _02280_);
  nor (_02290_, _02289_, _02270_);
  and (_02291_, _25556_, _24174_);
  and (_02292_, _02291_, _24179_);
  nor (_02293_, _02292_, _02290_);
  and (_02294_, _25602_, _24174_);
  nor (_02295_, _02294_, rst);
  and (_22652_, _02295_, _02293_);
  and (_02296_, _02232_, _23996_);
  and (_02297_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  or (_27021_, _02297_, _02296_);
  and (_02298_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_02299_, _01814_, _23989_);
  not (_02300_, _01816_);
  not (_02301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_02302_, _01823_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_02303_, _02302_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_02304_, _02209_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_02305_, _02304_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_02306_, _02305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_02307_, _02306_, _02303_);
  nand (_02308_, _02307_, _02205_);
  nor (_02309_, _02308_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_02310_, _02309_, _02301_);
  and (_02311_, _02309_, _02301_);
  or (_02312_, _02311_, _02310_);
  and (_02313_, _02312_, _02198_);
  or (_02314_, _01826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not (_02315_, _01827_);
  and (_02316_, _01829_, _02315_);
  and (_02317_, _02316_, _02314_);
  and (_02318_, _02210_, _02303_);
  or (_02319_, _02318_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not (_02320_, _02219_);
  and (_02321_, _02303_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_02322_, _02210_, _02321_);
  nor (_02323_, _02322_, _02320_);
  and (_02324_, _02323_, _02319_);
  or (_02325_, _02324_, _02317_);
  or (_02326_, _02325_, _02313_);
  or (_02328_, _02326_, _01814_);
  and (_02329_, _02328_, _02300_);
  and (_02330_, _02329_, _02299_);
  or (_02331_, _02330_, _02298_);
  and (_22653_, _02331_, _22731_);
  and (_02332_, _02232_, _24134_);
  and (_02333_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  or (_27020_, _02333_, _02332_);
  and (_02334_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_02335_, _02040_, _24089_);
  or (_22654_, _02335_, _02334_);
  and (_02336_, _02093_, _23548_);
  and (_02337_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_22655_, _02337_, _02336_);
  and (_02338_, _02039_, _24297_);
  not (_02339_, _02338_);
  and (_02340_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  and (_02341_, _02338_, _24134_);
  or (_22656_, _02341_, _02340_);
  and (_02343_, _02093_, _24219_);
  and (_02344_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_22657_, _02344_, _02343_);
  and (_02345_, _02232_, _24219_);
  and (_02346_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  or (_22658_, _02346_, _02345_);
  and (_02347_, _24017_, _23583_);
  and (_02348_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  or (_22659_, _02348_, _02347_);
  or (_02349_, _02019_, _26756_);
  or (_02350_, _02349_, _23840_);
  or (_02351_, _02021_, _02015_);
  and (_02352_, _26760_, _23708_);
  or (_02353_, _02352_, _23841_);
  or (_02354_, _02353_, _02351_);
  or (_02355_, _02354_, _02350_);
  and (_02356_, _02355_, _22737_);
  and (_02357_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_02358_, _26675_);
  and (_02359_, _02358_, _02003_);
  and (_02360_, _02351_, _26573_);
  or (_02361_, _02360_, _02359_);
  or (_02362_, _02361_, _02357_);
  or (_02363_, _02362_, _02356_);
  and (_26848_[1], _02363_, _22731_);
  and (_02364_, _24365_, _24297_);
  and (_02365_, _02364_, _23583_);
  not (_02366_, _02364_);
  and (_02367_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_27208_, _02367_, _02365_);
  and (_02368_, _24408_, _24159_);
  and (_02369_, _02368_, _24051_);
  not (_02370_, _02368_);
  and (_02371_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  or (_27152_, _02371_, _02369_);
  and (_02372_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  and (_02373_, _02338_, _23996_);
  or (_22660_, _02373_, _02372_);
  and (_02374_, _26743_, _26736_);
  and (_02375_, _26698_, _23779_);
  or (_02376_, _01992_, _26760_);
  or (_02377_, _02376_, _02375_);
  or (_02378_, _23805_, _23800_);
  and (_02379_, _02378_, _23803_);
  or (_02380_, _02379_, _26724_);
  or (_02381_, _02380_, _02377_);
  nor (_02382_, _02381_, _02015_);
  nand (_02383_, _02382_, _02374_);
  or (_02384_, _02022_, _26721_);
  or (_02385_, _23841_, _23839_);
  and (_02386_, _23772_, _23824_);
  or (_02387_, _02386_, _02385_);
  or (_02388_, _02387_, _02384_);
  or (_02389_, _26691_, _23830_);
  or (_02390_, _02389_, _23828_);
  or (_02391_, _02390_, _02388_);
  or (_02392_, _02391_, _02350_);
  or (_02393_, _02392_, _02383_);
  and (_02394_, _02393_, _22737_);
  and (_02395_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_02396_, _26595_, _23708_);
  and (_02397_, _02396_, _26573_);
  and (_02398_, _26581_, _26573_);
  or (_02399_, _02398_, _02359_);
  or (_02400_, _02399_, _02397_);
  or (_02401_, _02400_, _02395_);
  or (_02402_, _02401_, _02394_);
  and (_26853_, _02402_, _22731_);
  and (_02403_, _02368_, _23583_);
  and (_02404_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  or (_22661_, _02404_, _02403_);
  and (_02405_, _02368_, _23548_);
  and (_02406_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  or (_22662_, _02406_, _02405_);
  and (_02407_, _02045_, _23887_);
  and (_02408_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_22663_, _02408_, _02407_);
  and (_02409_, _02368_, _24219_);
  and (_02410_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  or (_22664_, _02410_, _02409_);
  and (_02411_, _02065_, _23548_);
  and (_02412_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  or (_22665_, _02412_, _02411_);
  and (_02413_, _24408_, _24297_);
  and (_02414_, _02413_, _24134_);
  not (_02415_, _02413_);
  and (_02416_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_22666_, _02416_, _02414_);
  and (_02417_, _02413_, _24089_);
  and (_02418_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_27149_, _02418_, _02417_);
  and (_02419_, _02413_, _23887_);
  and (_02420_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_27148_, _02420_, _02419_);
  and (_02421_, _24497_, _24134_);
  and (_02422_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  or (_27245_, _02422_, _02421_);
  or (_02423_, _02386_, _02021_);
  or (_02424_, _02423_, _02389_);
  or (_02425_, _02424_, _02383_);
  and (_02426_, _02425_, _22737_);
  and (_02427_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02428_, _02427_, _02400_);
  or (_02429_, _02428_, _02426_);
  and (_26848_[0], _02429_, _22731_);
  and (_02430_, _24497_, _24051_);
  and (_02431_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  or (_22667_, _02431_, _02430_);
  and (_02432_, _25413_, _24016_);
  and (_02433_, _02432_, _23996_);
  not (_02434_, _02432_);
  and (_02435_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  or (_22668_, _02435_, _02433_);
  and (_02436_, _02413_, _23548_);
  and (_02437_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_22669_, _02437_, _02436_);
  and (_02438_, _24188_, _22868_);
  and (_02439_, _02438_, _24533_);
  and (_02440_, _02439_, _22731_);
  and (_02441_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_02442_, _02273_, _02253_);
  and (_02443_, _02442_, _02271_);
  and (_02444_, _02266_, _02237_);
  nor (_02445_, _02444_, _02443_);
  and (_02446_, _02445_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_02447_, _02445_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_02448_, _02447_, _02446_);
  nor (_02449_, _02448_, _02292_);
  not (_02450_, _24126_);
  and (_02451_, _02292_, _02450_);
  or (_02452_, _02451_, _02449_);
  and (_02453_, _02452_, _02295_);
  or (_22670_, _02453_, _02441_);
  and (_02455_, _24408_, _24016_);
  and (_02456_, _02455_, _24134_);
  not (_02458_, _02455_);
  and (_02459_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_22671_, _02459_, _02456_);
  and (_02460_, _02455_, _24089_);
  and (_02461_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_22672_, _02461_, _02460_);
  and (_02462_, _02232_, _23583_);
  and (_02463_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  or (_22673_, _02463_, _02462_);
  and (_02465_, _02232_, _23887_);
  and (_02467_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  or (_22674_, _02467_, _02465_);
  and (_02468_, _02232_, _23548_);
  and (_02469_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  or (_27019_, _02469_, _02468_);
  and (_02470_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  and (_02471_, _02338_, _23887_);
  or (_22675_, _02471_, _02470_);
  and (_02472_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  and (_02473_, _02338_, _23548_);
  or (_27025_, _02473_, _02472_);
  nand (_02474_, _26406_, _23531_);
  or (_02475_, _23531_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_02476_, _02475_, _22731_);
  and (_22676_, _02476_, _02474_);
  and (_02478_, _24899_, _24496_);
  and (_02479_, _02478_, _24134_);
  not (_02480_, _02478_);
  and (_02481_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_22677_, _02481_, _02479_);
  and (_02483_, _02455_, _23887_);
  and (_02484_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_22678_, _02484_, _02483_);
  and (_02485_, _02478_, _23996_);
  and (_02486_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or (_22679_, _02486_, _02485_);
  and (_02488_, _24349_, _24006_);
  and (_02489_, _02488_, _24089_);
  not (_02490_, _02488_);
  and (_02491_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  or (_22680_, _02491_, _02489_);
  and (_02492_, _02364_, _24089_);
  and (_02494_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_22681_, _02494_, _02492_);
  nand (_02495_, _24299_, _22847_);
  and (_02497_, _02495_, _24003_);
  and (_02498_, _02497_, _24159_);
  and (_02499_, _02498_, _24089_);
  not (_02500_, _02498_);
  and (_02501_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_22682_, _02501_, _02499_);
  and (_02502_, _24496_, _23941_);
  and (_02503_, _02502_, _24219_);
  not (_02504_, _02502_);
  and (_02505_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or (_27248_, _02505_, _02503_);
  and (_02507_, _02455_, _23548_);
  and (_02508_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_27145_, _02508_, _02507_);
  and (_02509_, _02498_, _23583_);
  and (_02511_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_22683_, _02511_, _02509_);
  and (_02512_, _24004_, _22977_);
  and (_02513_, _02512_, _24146_);
  not (_02514_, _02513_);
  and (_02515_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  and (_02516_, _02513_, _24089_);
  or (_22684_, _02516_, _02515_);
  and (_02517_, _24408_, _24236_);
  and (_02518_, _02517_, _23996_);
  not (_02519_, _02517_);
  and (_02520_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  or (_27143_, _02520_, _02518_);
  and (_02521_, _02517_, _24051_);
  and (_02522_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  or (_22685_, _02522_, _02521_);
  and (_02523_, _02517_, _23583_);
  and (_02524_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  or (_22686_, _02524_, _02523_);
  and (_02525_, _24889_, _23583_);
  and (_02526_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_22687_, _02526_, _02525_);
  and (_02527_, _24698_, _24543_);
  and (_02528_, _02527_, _24594_);
  nand (_02530_, _02528_, _23504_);
  or (_02531_, _02528_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_02532_, _25227_, _24628_);
  not (_02534_, _02532_);
  and (_02535_, _02534_, _02531_);
  and (_02536_, _02535_, _02530_);
  nor (_02537_, _02534_, _24126_);
  or (_02539_, _02537_, _02536_);
  and (_22690_, _02539_, _22731_);
  and (_02540_, _02527_, _24607_);
  nand (_02541_, _02540_, _23504_);
  or (_02542_, _02540_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_02543_, _02542_, _02534_);
  and (_02544_, _02543_, _02541_);
  nor (_02545_, _02534_, _24043_);
  or (_02546_, _02545_, _02544_);
  and (_22691_, _02546_, _22731_);
  and (_02548_, _24638_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_02549_, _02548_, _24637_);
  and (_02550_, _02549_, _02527_);
  not (_02551_, _02527_);
  or (_02552_, _02551_, _24643_);
  and (_02553_, _02552_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_02555_, _02553_, _02532_);
  or (_02556_, _02555_, _02550_);
  nand (_02557_, _02532_, _24082_);
  and (_02558_, _02557_, _22731_);
  and (_22692_, _02558_, _02556_);
  and (_02560_, _02527_, _24533_);
  nand (_02561_, _02560_, _23504_);
  or (_02562_, _02560_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_02563_, _02562_, _02534_);
  and (_02564_, _02563_, _02561_);
  and (_02565_, _02532_, _23577_);
  or (_02566_, _02565_, _02564_);
  and (_22693_, _02566_, _22731_);
  nor (_02568_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_02569_, _02568_);
  nor (_02570_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_02571_, _02570_, _02569_);
  and (_02572_, _02571_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not (_02573_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor (_02574_, _02571_, _02573_);
  or (_02576_, _02574_, _02572_);
  or (_02577_, _02576_, _02527_);
  not (_02578_, _24562_);
  nor (_02580_, _02578_, _23504_);
  or (_02581_, _24562_, _02573_);
  nand (_02582_, _02581_, _02527_);
  or (_02583_, _02582_, _02580_);
  and (_02584_, _02583_, _02577_);
  or (_02585_, _02584_, _02532_);
  or (_02586_, _02534_, _23880_);
  and (_02587_, _02586_, _22731_);
  and (_22694_, _02587_, _02585_);
  or (_02588_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_02589_, _02588_, _02527_);
  and (_02590_, _24177_, _24531_);
  not (_02591_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_02592_, _24177_, _02591_);
  nand (_02593_, _02592_, _02527_);
  or (_02594_, _02593_, _02590_);
  and (_02595_, _02594_, _02589_);
  or (_02596_, _02595_, _02532_);
  nand (_02597_, _02532_, _23542_);
  and (_02598_, _02597_, _22731_);
  and (_22695_, _02598_, _02596_);
  and (_02599_, _24577_, _24531_);
  not (_02600_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_02601_, _24577_, _02600_);
  nand (_02602_, _02601_, _02527_);
  or (_02603_, _02602_, _02599_);
  not (_02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_02605_, _02604_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_02606_, _02605_, _02568_);
  and (_02607_, _02606_, _02570_);
  or (_02608_, _02607_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_02609_, _02608_, _02527_);
  and (_02610_, _02609_, _02603_);
  or (_02611_, _02610_, _02532_);
  nand (_02612_, _02532_, _24210_);
  and (_02613_, _02612_, _22731_);
  and (_22696_, _02613_, _02611_);
  nand (_02614_, _02294_, _23989_);
  nor (_02615_, _02283_, _02237_);
  and (_02616_, _25557_, _24174_);
  or (_02617_, _02616_, _02615_);
  and (_02618_, _02617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or (_02619_, _02284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_02620_, _02263_, _02248_);
  nor (_02621_, _02620_, _02615_);
  and (_02622_, _02621_, _02619_);
  and (_02623_, _02620_, _02283_);
  and (_02624_, _02623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_02625_, _02624_, _02622_);
  nor (_02626_, _02625_, _02616_);
  or (_02627_, _02626_, _02618_);
  or (_02628_, _02627_, _02294_);
  and (_02629_, _02628_, _22731_);
  and (_22697_, _02629_, _02614_);
  or (_02630_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_02631_, _02630_, _22731_);
  nand (_02632_, _02071_, _24126_);
  and (_22698_, _02632_, _02631_);
  or (_02633_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_02634_, _02633_, _22731_);
  nand (_02635_, _02071_, _24043_);
  and (_22699_, _02635_, _02634_);
  or (_02636_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_02637_, _02636_, _22731_);
  or (_02638_, _02074_, _23577_);
  and (_22700_, _02638_, _02637_);
  or (_02639_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_02640_, _02639_, _22731_);
  nand (_02641_, _02071_, _23542_);
  and (_22701_, _02641_, _02640_);
  nand (_02642_, _02071_, _24210_);
  or (_02643_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_02644_, _02643_, _22731_);
  and (_22702_, _02644_, _02642_);
  not (_02645_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_02646_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_02647_, _02646_, _02568_);
  and (_02648_, _02569_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_02649_, _02648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_02650_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_02651_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_02652_, _02651_, _02650_);
  and (_02653_, _02652_, _02649_);
  nor (_02654_, _02653_, _02647_);
  nor (_02655_, _02654_, _02645_);
  and (_02656_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor (_02657_, _02656_, _02655_);
  and (_02658_, _25227_, _24182_);
  nor (_02659_, _02658_, _02657_);
  not (_02660_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_02661_, _02660_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_02662_, _02661_, _02569_);
  and (_02663_, _02662_, _02658_);
  or (_02664_, _02663_, _02659_);
  and (_22703_, _02664_, _22731_);
  and (_02665_, _02658_, _02569_);
  nand (_02666_, _02665_, _23989_);
  and (_02668_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  not (_02669_, _02654_);
  and (_02670_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_02671_, _02670_, _02668_);
  or (_02672_, _02671_, _02658_);
  and (_02673_, _02672_, _22731_);
  and (_22704_, _02673_, _02666_);
  not (_02674_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_02675_, _02658_, _02660_);
  and (_02676_, _02675_, _02674_);
  and (_02677_, _02676_, _25554_);
  and (_02678_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_02679_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_02680_, _02679_, _02678_);
  nor (_02681_, _02680_, _02658_);
  and (_02682_, _02665_, _02450_);
  or (_02683_, _02682_, _02681_);
  or (_02684_, _02683_, _02677_);
  and (_22705_, _02684_, _22731_);
  and (_02685_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_02686_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_02687_, _02686_, _02685_);
  nor (_02688_, _02687_, _02658_);
  not (_02689_, _24043_);
  and (_02690_, _02665_, _02689_);
  and (_02691_, _02658_, _02568_);
  and (_02692_, _02691_, _02450_);
  or (_02693_, _02692_, _02690_);
  or (_02694_, _02693_, _02688_);
  and (_22706_, _02694_, _22731_);
  and (_02695_, _02676_, _02689_);
  and (_02696_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_02697_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor (_02698_, _02697_, _02696_);
  nor (_02699_, _02698_, _02658_);
  not (_02700_, _24082_);
  and (_02701_, _02665_, _02700_);
  or (_02702_, _02701_, _02699_);
  or (_02703_, _02702_, _02695_);
  and (_22707_, _02703_, _22731_);
  and (_02704_, _02665_, _23577_);
  and (_02705_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_02706_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_02707_, _02706_, _02705_);
  nor (_02708_, _02707_, _02658_);
  and (_02709_, _02691_, _02700_);
  or (_02710_, _02709_, _02708_);
  or (_02711_, _02710_, _02704_);
  and (_22708_, _02711_, _22731_);
  and (_02712_, _02676_, _23577_);
  and (_02713_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_02714_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_02715_, _02714_, _02713_);
  nor (_02716_, _02715_, _02658_);
  and (_02717_, _02665_, _23880_);
  or (_02718_, _02717_, _02716_);
  or (_02720_, _02718_, _02712_);
  and (_22709_, _02720_, _22731_);
  and (_02722_, _02676_, _23880_);
  and (_02723_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_02724_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_02726_, _02724_, _02723_);
  nor (_02727_, _02726_, _02658_);
  not (_02728_, _23542_);
  and (_02729_, _02665_, _02728_);
  or (_02730_, _02729_, _02727_);
  or (_02731_, _02730_, _02722_);
  and (_22710_, _02731_, _22731_);
  and (_02732_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_02733_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_02734_, _02733_, _02732_);
  nor (_02735_, _02734_, _02658_);
  and (_02737_, _02665_, _24671_);
  or (_02738_, _02737_, _02735_);
  and (_02739_, _02691_, _02728_);
  or (_02740_, _02739_, _02738_);
  and (_22711_, _02740_, _22731_);
  or (_02742_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_02743_, _02647_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_02744_, _02743_, _02653_);
  and (_02745_, _02744_, _02742_);
  nor (_02746_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nor (_02748_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_02749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_02750_, _02749_, _02748_);
  and (_02752_, _02750_, _02746_);
  nor (_02753_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_02754_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_02755_, _02754_, _02753_);
  and (_02756_, _02755_, _02647_);
  and (_02757_, _02756_, _02752_);
  and (_02758_, _02757_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_02759_, _02758_, _02745_);
  nor (_02760_, _02759_, _02658_);
  and (_02761_, _02691_, _24671_);
  or (_02762_, _02761_, _02760_);
  and (_22712_, _02762_, _22731_);
  and (_02764_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  and (_02765_, _02338_, _24089_);
  or (_22713_, _02765_, _02764_);
  and (_02767_, _25413_, _24349_);
  and (_02768_, _02767_, _23996_);
  not (_02769_, _02767_);
  and (_02771_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_27175_, _02771_, _02768_);
  and (_02772_, _02488_, _23887_);
  and (_02774_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  or (_22714_, _02774_, _02772_);
  and (_02775_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  and (_02776_, _02338_, _23583_);
  or (_27026_, _02776_, _02775_);
  and (_02777_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_02778_, _02777_, _02569_);
  not (_02779_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_02780_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _02779_);
  not (_02782_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_02783_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _02782_);
  and (_02784_, _02783_, _02780_);
  and (_02785_, _02784_, _02778_);
  not (_02786_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_02787_, _02786_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_02789_, _02568_, _02600_);
  and (_02790_, _02789_, _02787_);
  and (_02792_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_02793_, _02792_, _02569_);
  nor (_02794_, _02793_, _02790_);
  nor (_02795_, _02794_, _02778_);
  or (_02796_, _02795_, _02785_);
  and (_02798_, _02568_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_02799_, _02798_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or (_02800_, _02799_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_02801_, _02800_, _02796_);
  nor (_02802_, _02799_, _02785_);
  or (_02803_, _02802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02804_, _02803_, _02080_);
  and (_02806_, _02804_, _02801_);
  or (_22715_, _02806_, _02079_);
  and (_22716_, t0_i, _22731_);
  and (_02807_, _02498_, _23996_);
  and (_02809_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_22717_, _02809_, _02807_);
  not (_02810_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not (_02811_, _02802_);
  nor (_02812_, _02811_, _02795_);
  nor (_02813_, _02812_, _02810_);
  or (_02814_, _02813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_02815_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _02810_);
  or (_02816_, _02815_, _02802_);
  and (_02817_, _02816_, _22731_);
  and (_22718_, _02817_, _02814_);
  and (_02818_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_02819_, _02811_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  not (_02820_, _02778_);
  nor (_02821_, _02784_, _02820_);
  and (_02823_, _02821_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nor (_02824_, _02778_, _02790_);
  or (_02825_, _02824_, _02823_);
  nor (_02826_, _02793_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nor (_02827_, _02826_, _02799_);
  and (_02829_, _02827_, _02825_);
  or (_02830_, _02829_, _02819_);
  and (_02831_, _02830_, _02080_);
  or (_22719_, _02831_, _02818_);
  and (_02832_, _02488_, _23548_);
  and (_02833_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  or (_22720_, _02833_, _02832_);
  and (_02834_, _02498_, _24134_);
  and (_02835_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_22721_, _02835_, _02834_);
  and (_02836_, _02039_, _24016_);
  not (_02837_, _02836_);
  and (_02838_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  and (_02839_, _02836_, _24134_);
  or (_27024_, _02839_, _02838_);
  not (_02840_, _02812_);
  or (_02841_, _02840_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_02842_, _02802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_02844_, _02842_, _02080_);
  and (_02845_, _02844_, _02841_);
  or (_22722_, _02845_, _02085_);
  and (_02846_, _02478_, _23583_);
  and (_02847_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  or (_27247_, _02847_, _02846_);
  and (_02848_, _02517_, _23887_);
  and (_02849_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  or (_22723_, _02849_, _02848_);
  and (_02851_, _02432_, _24051_);
  and (_02852_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  or (_22724_, _02852_, _02851_);
  and (_02854_, _02784_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_02855_, _02854_, _02794_);
  or (_02856_, _02855_, _02812_);
  and (_02857_, _02856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_02858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _02810_);
  nand (_02859_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_02860_, _02859_, _02802_);
  or (_02861_, _02860_, _02858_);
  or (_02862_, _02861_, _02857_);
  and (_22725_, _02862_, _22731_);
  nor (_02863_, _02793_, _02778_);
  or (_02865_, _02863_, _02810_);
  or (_02866_, _02865_, _02782_);
  and (_02867_, _02778_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02868_, _02867_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_02869_, _02868_, _22731_);
  and (_22726_, _02869_, _02866_);
  nand (_02870_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22731_);
  nor (_02871_, _02870_, _02813_);
  or (_02872_, _02855_, _02811_);
  and (_02873_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_02874_, _02873_, _02872_);
  or (_22727_, _02874_, _02871_);
  and (_02875_, _02865_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_02876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_02877_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_02879_, _02877_, _02876_);
  and (_02880_, _02879_, _02867_);
  or (_02881_, _02880_, _02875_);
  and (_22728_, _02881_, _22731_);
  and (_02882_, _02497_, _24297_);
  and (_02883_, _02882_, _24134_);
  not (_02884_, _02882_);
  and (_02885_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_22729_, _02885_, _02883_);
  or (_02886_, _02649_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_02887_, _02649_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_02888_, _02887_, rst);
  nand (_02889_, _02888_, _02886_);
  nor (_22730_, _02889_, _02658_);
  and (_02890_, _24408_, _24349_);
  and (_02891_, _02890_, _23996_);
  not (_02892_, _02890_);
  and (_02893_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  or (_22739_, _02893_, _02891_);
  and (_02894_, _02478_, _24089_);
  and (_02895_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or (_22743_, _02895_, _02894_);
  and (_02896_, _02876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02897_, _02896_, _02779_);
  and (_02898_, _02867_, _02897_);
  or (_02899_, _02898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not (_02900_, rxd_i);
  nand (_02901_, _02898_, _02900_);
  and (_02902_, _02901_, _22731_);
  and (_22748_, _02902_, _02899_);
  and (_02903_, _02882_, _24051_);
  and (_02904_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_26986_, _02904_, _02903_);
  or (_02905_, _02887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_02906_, _02887_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_02907_, _02906_, rst);
  nand (_02908_, _02907_, _02905_);
  nor (_22754_, _02908_, _02658_);
  nor (_02909_, _02906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_02910_, _02906_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_02911_, _02910_, _02909_);
  nand (_02912_, _02911_, _22731_);
  nor (_22756_, _02912_, _02658_);
  or (_02913_, _02813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_02914_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _02810_);
  or (_02915_, _02914_, _02802_);
  and (_02916_, _02915_, _22731_);
  and (_22765_, _02916_, _02913_);
  and (_02917_, _02882_, _24089_);
  and (_02918_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_22770_, _02918_, _02917_);
  and (_02919_, _02478_, _24051_);
  and (_02920_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_22787_, _02920_, _02919_);
  and (_02921_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  and (_02922_, _02836_, _23996_);
  or (_22798_, _02922_, _02921_);
  and (_02923_, _02865_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nor (_02925_, _02896_, _02820_);
  or (_02926_, _02925_, _02923_);
  and (_02927_, _02876_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02928_, _02927_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02929_, _02928_, _22731_);
  and (_22807_, _02929_, _02926_);
  and (_02930_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_22819_, _02930_, _02818_);
  and (_02931_, _02498_, _24219_);
  and (_02932_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  or (_27007_, _02932_, _02931_);
  and (_02934_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_02935_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_22842_, _02935_, _02934_);
  and (_02936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02937_, _02936_, _02858_);
  and (_22848_, _02937_, _22731_);
  and (_02938_, _02890_, _24134_);
  and (_02939_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  or (_22860_, _02939_, _02938_);
  and (_02940_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02941_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_22870_, _02941_, _02940_);
  and (_02942_, _02882_, _23996_);
  and (_02943_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_22873_, _02943_, _02942_);
  and (_02944_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  and (_02945_, _02836_, _23887_);
  or (_22879_, _02945_, _02944_);
  or (_02946_, _02813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_02947_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _02810_);
  or (_02948_, _02947_, _02802_);
  and (_02949_, _02948_, _22731_);
  and (_22883_, _02949_, _02946_);
  or (_02950_, _02840_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_02951_, _02802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_02952_, _02951_, _02080_);
  and (_02953_, _02952_, _02950_);
  or (_22889_, _02953_, _02083_);
  or (_02954_, _02813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_02955_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _02810_);
  or (_02956_, _02955_, _02802_);
  and (_02957_, _02956_, _22731_);
  and (_22892_, _02957_, _02954_);
  or (_02958_, _02813_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_02959_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _02810_);
  or (_02960_, _02959_, _02802_);
  and (_02961_, _02960_, _22731_);
  and (_22895_, _02961_, _02958_);
  and (_02962_, _02890_, _24089_);
  and (_02963_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  or (_22915_, _02963_, _02962_);
  and (_02964_, _24476_, _24236_);
  and (_02965_, _02964_, _23996_);
  not (_02966_, _02964_);
  and (_02967_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_27187_, _02967_, _02965_);
  and (_02968_, _02890_, _23887_);
  and (_02969_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  or (_22929_, _02969_, _02968_);
  and (_02970_, _24301_, _24016_);
  and (_02971_, _02970_, _23583_);
  not (_02972_, _02970_);
  and (_02973_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  or (_22939_, _02973_, _02971_);
  and (_02974_, _24497_, _23583_);
  and (_02975_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or (_22944_, _02975_, _02974_);
  and (_02976_, _02882_, _24219_);
  and (_02977_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_22955_, _02977_, _02976_);
  and (_02978_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  and (_02979_, _02836_, _24089_);
  or (_22959_, _02979_, _02978_);
  and (_02980_, _02497_, _24016_);
  and (_02981_, _02980_, _23996_);
  not (_02982_, _02980_);
  and (_02983_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_23014_, _02983_, _02981_);
  and (_02984_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  and (_02985_, _02836_, _23583_);
  or (_23021_, _02985_, _02984_);
  and (_02986_, _02882_, _23548_);
  and (_02987_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_23046_, _02987_, _02986_);
  and (_02988_, _02882_, _23887_);
  and (_02989_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_23077_, _02989_, _02988_);
  and (_02990_, _24899_, _23945_);
  and (_02991_, _02990_, _24089_);
  not (_02992_, _02990_);
  and (_02993_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  or (_27055_, _02993_, _02991_);
  and (_02994_, _02970_, _23887_);
  and (_02995_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  or (_23102_, _02995_, _02994_);
  and (_02996_, _24301_, _24140_);
  and (_02997_, _02996_, _23583_);
  not (_02998_, _02996_);
  and (_02999_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  or (_23110_, _02999_, _02997_);
  and (_03001_, _24372_, _24301_);
  and (_03002_, _03001_, _23548_);
  not (_03003_, _03001_);
  and (_03004_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_23135_, _03004_, _03002_);
  and (_03005_, _02980_, _23583_);
  and (_03006_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_23153_, _03006_, _03005_);
  and (_03007_, _02980_, _23887_);
  and (_03008_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_23165_, _03008_, _03007_);
  nor (_26867_[2], _00223_, rst);
  and (_03009_, _24518_, _24219_);
  and (_03010_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  or (_23171_, _03010_, _03009_);
  and (_03011_, _02512_, _24372_);
  not (_03013_, _03011_);
  and (_03014_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  and (_03015_, _03011_, _24219_);
  or (_23180_, _03015_, _03014_);
  nor (_26877_[4], _00676_, rst);
  and (_03016_, _02990_, _23548_);
  and (_03017_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  or (_23200_, _03017_, _03016_);
  and (_03018_, _02980_, _24051_);
  and (_03019_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_26971_, _03019_, _03018_);
  and (_03020_, _02497_, _24236_);
  and (_03021_, _03020_, _23996_);
  not (_03022_, _03020_);
  and (_03023_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_26952_, _03023_, _03021_);
  and (_03024_, _03020_, _24134_);
  and (_03025_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_23303_, _03025_, _03024_);
  and (_03026_, _24474_, _23945_);
  and (_03028_, _03026_, _24051_);
  not (_03029_, _03026_);
  and (_03030_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_23307_, _03030_, _03028_);
  and (_03031_, _24237_, _24051_);
  and (_03032_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_23315_, _03032_, _03031_);
  and (_03033_, _25413_, _24372_);
  and (_03034_, _03033_, _24089_);
  not (_03035_, _03033_);
  and (_03036_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or (_23326_, _03036_, _03034_);
  and (_03037_, _03026_, _23996_);
  and (_03038_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_23332_, _03038_, _03037_);
  and (_03039_, _02980_, _24219_);
  and (_03040_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_23339_, _03040_, _03039_);
  and (_03041_, _03026_, _24134_);
  and (_03042_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_27052_, _03042_, _03041_);
  and (_03043_, _24496_, _24236_);
  and (_03044_, _03043_, _24051_);
  not (_03045_, _03043_);
  and (_03046_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  or (_23365_, _03046_, _03044_);
  nor (_26877_[3], _00592_, rst);
  and (_03048_, _02497_, _24349_);
  and (_03049_, _03048_, _23996_);
  not (_03050_, _03048_);
  and (_03052_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  or (_26933_, _03052_, _03049_);
  and (_03054_, _24442_, _24089_);
  and (_03055_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  or (_23384_, _03055_, _03054_);
  and (_03057_, _03048_, _24134_);
  and (_03058_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_23389_, _03058_, _03057_);
  and (_03059_, _03048_, _24051_);
  and (_03060_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_23394_, _03060_, _03059_);
  and (_03061_, _03026_, _23583_);
  and (_03062_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_23428_, _03062_, _03061_);
  and (_03065_, _03020_, _24219_);
  and (_03066_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  or (_23431_, _03066_, _03065_);
  and (_03067_, _03020_, _23887_);
  and (_03068_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_23435_, _03068_, _03067_);
  and (_03070_, _02432_, _24134_);
  and (_03071_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  or (_23502_, _03071_, _03070_);
  and (_03072_, _24497_, _23887_);
  and (_03073_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or (_27244_, _03073_, _03072_);
  nor (_03074_, _00287_, _26581_);
  nor (_03075_, _03074_, _26601_);
  nor (_03077_, _00239_, _23893_);
  and (_03078_, _03077_, _23902_);
  and (_03080_, _03078_, _23931_);
  and (_03081_, _03080_, _02374_);
  nor (_03082_, _03081_, _24279_);
  nor (_03083_, _03082_, _03075_);
  nor (_26892_, _03083_, rst);
  and (_03084_, _24298_, _24173_);
  and (_03085_, _03084_, _25024_);
  and (_03086_, _03085_, _22978_);
  nand (_03087_, _03086_, _23989_);
  or (_03088_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_03089_, _03088_, _22731_);
  and (_26854_[7], _03089_, _03087_);
  and (_03090_, _03084_, _26779_);
  not (_03091_, _03090_);
  nor (_03093_, _03091_, _23989_);
  and (_03094_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_03096_, _03094_, _22979_);
  or (_03097_, _03096_, _03093_);
  or (_03098_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_03100_, _03098_, _22731_);
  and (_26855_[7], _03100_, _03097_);
  nor (_03101_, _03090_, _03085_);
  and (_03102_, _03084_, _24627_);
  not (_03104_, _03102_);
  and (_03105_, _03104_, _03101_);
  nor (_03106_, _03105_, _22979_);
  not (_03107_, _03106_);
  and (_03108_, _03107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_03109_, _03104_, _23989_);
  not (_03110_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_03111_, _03101_, _03110_);
  or (_03113_, _03111_, _03109_);
  and (_03114_, _03113_, _22978_);
  or (_03115_, _03114_, _03108_);
  and (_26856_[7], _03115_, _22731_);
  and (_03118_, _03084_, _24187_);
  and (_03119_, _03118_, _22978_);
  and (_03120_, _03119_, _25554_);
  nor (_03121_, _03118_, _03102_);
  and (_03122_, _03121_, _03101_);
  or (_03124_, _03122_, _22979_);
  or (_03126_, _03124_, _03106_);
  and (_03127_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_03128_, _03127_, _03120_);
  and (_26857_[7], _03128_, _22731_);
  nand (_03129_, _03121_, _03091_);
  and (_03131_, _03129_, _22978_);
  and (_03132_, _25226_, _24298_);
  and (_03133_, _03132_, _25024_);
  not (_03134_, _03133_);
  and (_03135_, _03134_, _03121_);
  and (_03136_, _03135_, _03091_);
  or (_03137_, _03085_, _22979_);
  or (_03138_, _03137_, _03136_);
  or (_03139_, _03138_, _03131_);
  and (_03140_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nand (_03141_, _03133_, _22978_);
  nor (_03142_, _03141_, _23989_);
  or (_03143_, _03142_, _03140_);
  and (_26858_[7], _03143_, _22731_);
  and (_03144_, _03132_, _26779_);
  and (_03145_, _03144_, _22978_);
  and (_03146_, _03145_, _25554_);
  nor (_03147_, _03144_, _03133_);
  and (_03148_, _03147_, _03122_);
  or (_03149_, _03137_, _03090_);
  nor (_03150_, _03149_, _03148_);
  nand (_03151_, _03150_, _03135_);
  and (_03152_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  or (_03153_, _03152_, _03146_);
  and (_26859_[7], _03153_, _22731_);
  and (_03155_, _03132_, _24627_);
  not (_03157_, _03155_);
  and (_03158_, _03157_, _03148_);
  or (_03159_, _03158_, _22979_);
  nor (_03161_, _03148_, _22979_);
  or (_03162_, _03161_, _03159_);
  and (_03164_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nand (_03165_, _03155_, _22978_);
  nor (_03166_, _03165_, _23989_);
  or (_03167_, _03166_, _03164_);
  and (_26860_[7], _03167_, _22731_);
  and (_03168_, _03132_, _24187_);
  and (_03169_, _03168_, _25554_);
  and (_03170_, _03168_, _22978_);
  not (_03171_, _03170_);
  and (_03172_, _03171_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or (_03173_, _03172_, _03169_);
  or (_03174_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_03175_, _03174_, _22731_);
  and (_26861_[7], _03175_, _03173_);
  nor (_26877_[2], _00496_, rst);
  and (_03176_, _03020_, _23548_);
  and (_03178_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_26951_, _03178_, _03176_);
  and (_03180_, _02497_, _23941_);
  and (_03181_, _03180_, _23996_);
  not (_03182_, _03180_);
  and (_03183_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_23678_, _03183_, _03181_);
  and (_03184_, _03048_, _24219_);
  and (_03185_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  or (_23725_, _03185_, _03184_);
  and (_03186_, _24056_, _23945_);
  and (_03187_, _03186_, _23583_);
  not (_03188_, _03186_);
  and (_03189_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  or (_27051_, _03189_, _03187_);
  nor (_26877_[1], _00415_, rst);
  and (_03190_, _03048_, _23583_);
  and (_03191_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_23849_, _03191_, _03190_);
  and (_03192_, _24330_, _23996_);
  and (_03193_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_23852_, _03193_, _03192_);
  and (_03194_, _03048_, _23887_);
  and (_03195_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_23866_, _03195_, _03194_);
  nor (_26877_[0], _26654_, rst);
  and (_03197_, _03180_, _23548_);
  and (_03198_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_23942_, _03198_, _03197_);
  and (_03199_, _03180_, _24219_);
  and (_03200_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_23956_, _03200_, _03199_);
  and (_03201_, _03186_, _24219_);
  and (_03202_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  or (_23961_, _03202_, _03201_);
  and (_03203_, _03186_, _24134_);
  and (_03204_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  or (_24007_, _03204_, _03203_);
  and (_03205_, _03180_, _23583_);
  and (_03207_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_24010_, _03207_, _03205_);
  and (_03208_, _03180_, _24051_);
  and (_03209_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_24012_, _03209_, _03208_);
  and (_03210_, _03180_, _24089_);
  and (_03211_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_24046_, _03211_, _03210_);
  and (_03212_, _03186_, _24051_);
  and (_03213_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  or (_24049_, _03213_, _03212_);
  and (_03214_, _03186_, _23996_);
  and (_03215_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  or (_24084_, _03215_, _03214_);
  and (_03217_, _02497_, _24899_);
  and (_03218_, _03217_, _23887_);
  not (_03219_, _03217_);
  and (_03220_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_24090_, _03220_, _03218_);
  and (_03221_, _02512_, _24319_);
  not (_03222_, _03221_);
  and (_03224_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  and (_03225_, _03221_, _23583_);
  or (_24103_, _03225_, _03224_);
  and (_03226_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  and (_03227_, _03221_, _23887_);
  or (_24128_, _03227_, _03226_);
  and (_03228_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  and (_03229_, _03221_, _23548_);
  or (_24135_, _03229_, _03228_);
  and (_03230_, _03217_, _24134_);
  and (_03231_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_24138_, _03231_, _03230_);
  and (_03232_, _03217_, _24051_);
  and (_03233_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_24168_, _03233_, _03232_);
  and (_03234_, _03217_, _24089_);
  and (_03235_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_27312_, _03235_, _03234_);
  and (_03236_, _24408_, _24095_);
  and (_03237_, _03236_, _23996_);
  not (_03238_, _03236_);
  and (_03239_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_24183_, _03239_, _03237_);
  and (_03241_, _25413_, _23941_);
  and (_03242_, _03241_, _24051_);
  not (_03243_, _03241_);
  and (_03244_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  or (_24191_, _03244_, _03242_);
  and (_03245_, _25413_, _24899_);
  and (_03246_, _03245_, _23996_);
  not (_03247_, _03245_);
  and (_03248_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  or (_24195_, _03248_, _03246_);
  and (_03249_, _03245_, _23548_);
  and (_03250_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  or (_24199_, _03250_, _03249_);
  and (_03251_, _02497_, _24474_);
  and (_03252_, _03251_, _24089_);
  not (_03253_, _03251_);
  and (_03254_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_24202_, _03254_, _03252_);
  and (_03255_, _25413_, _24474_);
  and (_03256_, _03255_, _23583_);
  not (_03257_, _03255_);
  and (_03258_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_24205_, _03258_, _03256_);
  and (_03259_, _03251_, _23583_);
  and (_03260_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_24211_, _03260_, _03259_);
  and (_03261_, _03236_, _24089_);
  and (_03263_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_24213_, _03263_, _03261_);
  and (_03264_, _03236_, _24134_);
  and (_03265_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_24215_, _03265_, _03264_);
  and (_03266_, _03251_, _23887_);
  and (_03267_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_27290_, _03267_, _03266_);
  and (_03269_, _25413_, _24056_);
  and (_03270_, _03269_, _24219_);
  not (_03271_, _03269_);
  and (_03272_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  or (_24222_, _03272_, _03270_);
  and (_03273_, _03251_, _23548_);
  and (_03274_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_27289_, _03274_, _03273_);
  and (_03275_, _25413_, _24223_);
  and (_03276_, _03275_, _24089_);
  not (_03277_, _03275_);
  and (_03278_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_24227_, _03278_, _03276_);
  and (_03279_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  and (_03280_, _02513_, _23996_);
  or (_24235_, _03280_, _03279_);
  and (_03281_, _25413_, _24319_);
  and (_03282_, _03281_, _24219_);
  not (_03283_, _03281_);
  and (_03284_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or (_24241_, _03284_, _03282_);
  and (_03285_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  and (_03286_, _03221_, _24134_);
  or (_24242_, _03286_, _03285_);
  and (_03287_, _25413_, _24095_);
  and (_03288_, _03287_, _24134_);
  not (_03289_, _03287_);
  and (_03290_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  or (_24252_, _03290_, _03288_);
  and (_03291_, _03251_, _23996_);
  and (_03292_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_24256_, _03292_, _03291_);
  and (_03293_, _03287_, _23887_);
  and (_03294_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  or (_24280_, _03294_, _03293_);
  and (_03295_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  and (_03296_, _03221_, _24051_);
  or (_24282_, _03296_, _03295_);
  and (_03298_, _03251_, _24134_);
  and (_03299_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_24285_, _03299_, _03298_);
  and (_03301_, _03251_, _24051_);
  and (_03302_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_24288_, _03302_, _03301_);
  and (_03303_, _03033_, _24051_);
  and (_03304_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or (_27162_, _03304_, _03303_);
  and (_03305_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  and (_03306_, _03221_, _24089_);
  or (_24316_, _03306_, _03305_);
  and (_03307_, _23944_, _22847_);
  and (_03308_, _24003_, _03307_);
  and (_03309_, _03308_, _24223_);
  and (_03310_, _03309_, _24219_);
  not (_03311_, _03309_);
  and (_03312_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  or (_26962_, _03312_, _03310_);
  and (_03313_, _25413_, _24297_);
  and (_03314_, _03313_, _23583_);
  not (_03315_, _03313_);
  and (_03316_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  or (_27177_, _03316_, _03314_);
  and (_03317_, _03313_, _24219_);
  and (_03318_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  or (_24326_, _03318_, _03317_);
  and (_03319_, _02512_, _22974_);
  not (_03320_, _03319_);
  and (_03322_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and (_03323_, _03319_, _23583_);
  or (_24329_, _03323_, _03322_);
  and (_03324_, _02497_, _24056_);
  and (_03325_, _03324_, _24134_);
  not (_03326_, _03324_);
  and (_03327_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_24335_, _03327_, _03325_);
  and (_03328_, _03324_, _24051_);
  and (_03329_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_24338_, _03329_, _03328_);
  and (_03330_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_03331_, _03319_, _24089_);
  or (_24344_, _03331_, _03330_);
  and (_03332_, _24518_, _23887_);
  and (_03333_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  or (_24346_, _03333_, _03332_);
  and (_03334_, _03324_, _23996_);
  and (_03335_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_24356_, _03335_, _03334_);
  and (_03337_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and (_03338_, _03319_, _24134_);
  or (_24359_, _03338_, _03337_);
  and (_03340_, _02488_, _24219_);
  and (_03341_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  or (_24363_, _03341_, _03340_);
  and (_03343_, _02497_, _24223_);
  and (_03344_, _03343_, _23996_);
  not (_03346_, _03343_);
  and (_03347_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_24366_, _03347_, _03344_);
  and (_03348_, _03324_, _24219_);
  and (_03349_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_27258_, _03349_, _03348_);
  and (_03350_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and (_03351_, _03319_, _23996_);
  or (_24370_, _03351_, _03350_);
  and (_03353_, _02767_, _24089_);
  and (_03354_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or (_24390_, _03354_, _03353_);
  and (_03355_, _24159_, _24141_);
  and (_03356_, _03355_, _23548_);
  not (_03357_, _03355_);
  and (_03358_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_24419_, _03358_, _03356_);
  and (_03360_, _25413_, _24236_);
  and (_03361_, _03360_, _24134_);
  not (_03362_, _03360_);
  and (_03363_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or (_24423_, _03363_, _03361_);
  and (_03364_, _03313_, _23996_);
  and (_03365_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  or (_24429_, _03365_, _03364_);
  and (_03366_, _03360_, _24089_);
  and (_03367_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_24432_, _03367_, _03366_);
  and (_03368_, _03324_, _23887_);
  and (_03369_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_24435_, _03369_, _03368_);
  and (_26840_[2], _23639_, _22731_);
  and (_03370_, _24408_, _22974_);
  and (_03371_, _03370_, _24219_);
  not (_03372_, _03370_);
  and (_03373_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_27117_, _03373_, _03371_);
  and (_03374_, _03370_, _23887_);
  and (_03375_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_24445_, _03375_, _03374_);
  and (_03376_, _03343_, _23887_);
  and (_03377_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_27243_, _03377_, _03376_);
  and (_03378_, _03343_, _23548_);
  and (_03379_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_24456_, _03379_, _03378_);
  and (_03380_, _03343_, _24219_);
  and (_03381_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_24463_, _03381_, _03380_);
  and (_03382_, _03287_, _23996_);
  and (_03383_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  or (_24466_, _03383_, _03382_);
  and (_03384_, _03355_, _24089_);
  and (_03385_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_24475_, _03385_, _03384_);
  and (_03386_, _03370_, _24051_);
  and (_03387_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_24477_, _03387_, _03386_);
  and (_03388_, _02432_, _23548_);
  and (_03390_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  or (_24483_, _03390_, _03388_);
  and (_03391_, _03370_, _24134_);
  and (_03392_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_24488_, _03392_, _03391_);
  and (_03393_, _02767_, _24051_);
  and (_03394_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_24498_, _03394_, _03393_);
  and (_03396_, _03343_, _24051_);
  and (_03397_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_24501_, _03397_, _03396_);
  and (_03398_, _03343_, _24089_);
  and (_03400_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or (_24506_, _03400_, _03398_);
  and (_03402_, _03343_, _23583_);
  and (_03403_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_24524_, _03403_, _03402_);
  not (_03404_, _03086_);
  and (_03405_, _03404_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_03406_, _03086_, _24671_);
  or (_03407_, _03406_, _03405_);
  and (_26854_[0], _03407_, _22731_);
  nand (_03408_, _03086_, _23542_);
  or (_03409_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_03410_, _03409_, _22731_);
  and (_26854_[1], _03410_, _03408_);
  or (_03411_, _03404_, _23880_);
  or (_03412_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_03413_, _03412_, _22731_);
  and (_26854_[2], _03413_, _03411_);
  or (_03414_, _03404_, _23577_);
  or (_03416_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_03417_, _03416_, _22731_);
  and (_26854_[3], _03417_, _03414_);
  nand (_03419_, _03086_, _24082_);
  or (_03420_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_03421_, _03420_, _22731_);
  and (_26854_[4], _03421_, _03419_);
  nand (_03423_, _03086_, _24043_);
  or (_03424_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_03425_, _03424_, _22731_);
  and (_26854_[5], _03425_, _03423_);
  nand (_03428_, _03086_, _24126_);
  or (_03429_, _03086_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_03430_, _03429_, _22731_);
  and (_26854_[6], _03430_, _03428_);
  and (_03431_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_03432_, _03090_, _24671_);
  or (_03433_, _03432_, _22979_);
  or (_03434_, _03433_, _03431_);
  or (_03435_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_03436_, _03435_, _22731_);
  and (_26855_[0], _03436_, _03434_);
  nor (_03437_, _03091_, _23542_);
  and (_03438_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  or (_03439_, _03438_, _22979_);
  or (_03441_, _03439_, _03437_);
  or (_03442_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_03444_, _03442_, _22731_);
  and (_26855_[1], _03444_, _03441_);
  and (_03445_, _03090_, _23880_);
  and (_03446_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_03447_, _03446_, _22979_);
  or (_03448_, _03447_, _03445_);
  or (_03449_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_03450_, _03449_, _22731_);
  and (_26855_[2], _03450_, _03448_);
  and (_03451_, _03090_, _23577_);
  and (_03452_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_03453_, _03452_, _22979_);
  or (_03454_, _03453_, _03451_);
  or (_03455_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_03457_, _03455_, _22731_);
  and (_26855_[3], _03457_, _03454_);
  nor (_03458_, _03091_, _24082_);
  and (_03459_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_03460_, _03459_, _22979_);
  or (_03461_, _03460_, _03458_);
  or (_03462_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_03463_, _03462_, _22731_);
  and (_26855_[4], _03463_, _03461_);
  nor (_03464_, _03091_, _24043_);
  and (_03465_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_03466_, _03465_, _22979_);
  or (_03468_, _03466_, _03464_);
  or (_03469_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_03470_, _03469_, _22731_);
  and (_26855_[5], _03470_, _03468_);
  nor (_03471_, _03091_, _24126_);
  and (_03473_, _03091_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_03474_, _03473_, _22979_);
  or (_03476_, _03474_, _03471_);
  or (_03478_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_03479_, _03478_, _22731_);
  and (_26855_[6], _03479_, _03476_);
  and (_03481_, _03107_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nand (_03482_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_03484_, _03482_, _03101_);
  nor (_03485_, _24210_, _22979_);
  and (_03487_, _03485_, _03102_);
  or (_03488_, _03487_, _03484_);
  or (_03489_, _03488_, _03481_);
  and (_26856_[0], _03489_, _22731_);
  or (_03490_, _03101_, _22979_);
  nand (_03491_, _03490_, _03106_);
  and (_03492_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nand (_03493_, _03102_, _22978_);
  nor (_03494_, _03493_, _23542_);
  or (_03495_, _03494_, _03492_);
  and (_26856_[1], _03495_, _22731_);
  and (_03496_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_03497_, _23880_, _22978_);
  and (_03499_, _03497_, _03102_);
  or (_03500_, _03499_, _03496_);
  and (_26856_[2], _03500_, _22731_);
  and (_03501_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_03502_, _23577_, _22978_);
  and (_03503_, _03502_, _03102_);
  or (_03504_, _03503_, _03501_);
  and (_26856_[3], _03504_, _22731_);
  and (_03505_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_03506_, _24082_, _22979_);
  and (_03508_, _03506_, _03102_);
  or (_03510_, _03508_, _03505_);
  and (_26856_[4], _03510_, _22731_);
  and (_03512_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_03513_, _24043_, _22979_);
  and (_03514_, _03513_, _03102_);
  or (_03515_, _03514_, _03512_);
  and (_26856_[5], _03515_, _22731_);
  and (_03516_, _03491_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_03517_, _24126_, _22979_);
  and (_03518_, _03517_, _03102_);
  or (_03520_, _03518_, _03516_);
  and (_26856_[6], _03520_, _22731_);
  and (_03521_, _03119_, _24671_);
  and (_03522_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or (_03523_, _03522_, _03521_);
  and (_26857_[0], _03523_, _22731_);
  and (_03524_, _03119_, _02728_);
  and (_03525_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_03526_, _03525_, _03524_);
  and (_26857_[1], _03526_, _22731_);
  and (_03527_, _03119_, _23880_);
  and (_03528_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_03530_, _03528_, _03527_);
  and (_26857_[2], _03530_, _22731_);
  and (_03531_, _03119_, _23577_);
  and (_03532_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_03534_, _03532_, _03531_);
  and (_26857_[3], _03534_, _22731_);
  and (_03535_, _03119_, _02700_);
  and (_03536_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or (_03537_, _03536_, _03535_);
  and (_26857_[4], _03537_, _22731_);
  and (_03538_, _03119_, _02689_);
  and (_03540_, _03126_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_03541_, _03540_, _03538_);
  and (_26857_[5], _03541_, _22731_);
  and (_03542_, _03119_, _02450_);
  and (_03543_, _03124_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nand (_03544_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_03545_, _03544_, _03105_);
  or (_03546_, _03545_, _03543_);
  or (_03547_, _03546_, _03542_);
  and (_26857_[6], _03547_, _22731_);
  and (_03549_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_03550_, _03485_, _03133_);
  or (_03551_, _03550_, _03549_);
  and (_26858_[0], _03551_, _22731_);
  and (_03552_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_03554_, _23542_, _22979_);
  and (_03555_, _03554_, _03133_);
  or (_03556_, _03555_, _03552_);
  and (_26858_[1], _03556_, _22731_);
  and (_03557_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_03558_, _03497_, _03133_);
  or (_03559_, _03558_, _03557_);
  and (_26858_[2], _03559_, _22731_);
  and (_03561_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_03562_, _03502_, _03133_);
  or (_03563_, _03562_, _03561_);
  and (_26858_[3], _03563_, _22731_);
  and (_03564_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_03565_, _03506_, _03133_);
  or (_03566_, _03565_, _03564_);
  and (_26858_[4], _03566_, _22731_);
  and (_03567_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_03568_, _03513_, _03133_);
  or (_03569_, _03568_, _03567_);
  and (_26858_[5], _03569_, _22731_);
  and (_03570_, _03139_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_03571_, _03517_, _03133_);
  or (_03572_, _03571_, _03570_);
  and (_26858_[6], _03572_, _22731_);
  and (_03574_, _03485_, _03144_);
  and (_03575_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  or (_03577_, _03575_, _03574_);
  and (_26859_[0], _03577_, _22731_);
  and (_03578_, _03145_, _02728_);
  and (_03579_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  or (_03580_, _03579_, _03578_);
  and (_26859_[1], _03580_, _22731_);
  and (_03581_, _03145_, _23880_);
  and (_03582_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  or (_03583_, _03582_, _03581_);
  and (_26859_[2], _03583_, _22731_);
  and (_03585_, _03145_, _23577_);
  and (_03586_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or (_03587_, _03586_, _03585_);
  and (_26859_[3], _03587_, _22731_);
  and (_03588_, _03145_, _02700_);
  and (_03589_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  or (_03590_, _03589_, _03588_);
  and (_26859_[4], _03590_, _22731_);
  and (_03591_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_03592_, _03145_, _02689_);
  or (_03593_, _03592_, _03591_);
  and (_26859_[5], _03593_, _22731_);
  and (_03594_, _03145_, _02450_);
  and (_03595_, _03151_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or (_03596_, _03595_, _03594_);
  and (_26859_[6], _03596_, _22731_);
  and (_03597_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_03599_, _03485_, _03155_);
  or (_03600_, _03599_, _03597_);
  and (_26860_[0], _03600_, _22731_);
  and (_03601_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_03602_, _03554_, _03155_);
  or (_03603_, _03602_, _03601_);
  and (_26860_[1], _03603_, _22731_);
  and (_03604_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_03606_, _03497_, _03155_);
  or (_03607_, _03606_, _03604_);
  and (_26860_[2], _03607_, _22731_);
  and (_03608_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_03610_, _03502_, _03155_);
  or (_03611_, _03610_, _03608_);
  and (_26860_[3], _03611_, _22731_);
  and (_03612_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_03613_, _03506_, _03155_);
  or (_03614_, _03613_, _03612_);
  and (_26860_[4], _03614_, _22731_);
  nor (_03615_, _03157_, _24043_);
  and (_03616_, _03157_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or (_03617_, _03616_, _22979_);
  or (_03618_, _03617_, _03615_);
  or (_03619_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_03620_, _03619_, _22731_);
  and (_26860_[5], _03620_, _03618_);
  and (_03621_, _03162_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_03622_, _03517_, _03155_);
  or (_03623_, _03622_, _03621_);
  and (_26860_[6], _03623_, _22731_);
  nand (_03624_, _03157_, _03147_);
  nor (_03625_, _03168_, _03624_);
  or (_03626_, _03625_, _22979_);
  and (_03628_, _03626_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_03629_, _03485_, _03168_);
  and (_03630_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_03632_, _03630_, _03624_);
  or (_03633_, _03632_, _03629_);
  or (_03634_, _03633_, _03628_);
  and (_26861_[0], _03634_, _22731_);
  and (_03635_, _03626_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_03636_, _03171_, _23542_);
  and (_03637_, _22978_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_03638_, _03637_, _03624_);
  or (_03639_, _03638_, _03636_);
  or (_03640_, _03639_, _03635_);
  and (_26861_[1], _03640_, _22731_);
  and (_03641_, _03170_, _23880_);
  or (_03642_, _03137_, _03129_);
  or (_03643_, _03642_, _03625_);
  and (_03644_, _03624_, _22978_);
  or (_03645_, _03644_, _03643_);
  and (_03646_, _03645_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or (_03647_, _03646_, _03641_);
  and (_26861_[2], _03647_, _22731_);
  and (_03649_, _03170_, _23577_);
  and (_03650_, _03645_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  or (_03651_, _03650_, _03649_);
  and (_26861_[3], _03651_, _22731_);
  nor (_03652_, _03171_, _24082_);
  and (_03653_, _03645_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or (_03654_, _03653_, _03652_);
  and (_26861_[4], _03654_, _22731_);
  and (_03655_, _03171_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_03656_, _03171_, _24043_);
  or (_03657_, _03656_, _03655_);
  and (_26861_[5], _03657_, _22731_);
  nor (_03658_, _03171_, _24126_);
  and (_03660_, _03645_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or (_03661_, _03660_, _03658_);
  and (_26861_[6], _03661_, _22731_);
  and (_03662_, _02512_, _24056_);
  not (_03663_, _03662_);
  and (_03665_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and (_03666_, _03662_, _23583_);
  or (_24958_, _03666_, _03665_);
  and (_03667_, _02497_, _24319_);
  and (_03668_, _03667_, _24089_);
  not (_03669_, _03667_);
  and (_03670_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  or (_25031_, _03670_, _03668_);
  and (_03672_, _02970_, _24051_);
  and (_03674_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  or (_25037_, _03674_, _03672_);
  and (_03676_, _02502_, _24051_);
  and (_03677_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or (_25076_, _03677_, _03676_);
  and (_03678_, _02890_, _24219_);
  and (_03679_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  or (_25079_, _03679_, _03678_);
  and (_03680_, _02502_, _24134_);
  and (_03681_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or (_25082_, _03681_, _03680_);
  and (_03682_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and (_03683_, _03662_, _23887_);
  or (_25087_, _03683_, _03682_);
  and (_03684_, _02970_, _23996_);
  and (_03685_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  or (_27229_, _03685_, _03684_);
  and (_03686_, _02970_, _24134_);
  and (_03687_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  or (_25170_, _03687_, _03686_);
  not (_03688_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_03689_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  and (_03690_, _03689_, _03688_);
  and (_03691_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _22731_);
  and (_27314_, _03691_, _03690_);
  nor (_03692_, _03690_, rst);
  nand (_03693_, _03689_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or (_03694_, _03689_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03696_, _03694_, _03693_);
  and (_27315_[3], _03696_, _03692_);
  not (_03698_, _00051_);
  nor (_03699_, _03698_, _00090_);
  not (_03700_, _00027_);
  and (_03702_, _03700_, _00143_);
  and (_03703_, _03702_, _26816_);
  and (_03705_, _03703_, _03699_);
  not (_03706_, _00325_);
  nand (_03707_, _00569_, _03706_);
  nor (_03708_, _24533_, _23195_);
  nor (_03709_, _03708_, _24534_);
  and (_03710_, _00329_, _00326_);
  not (_03711_, _03710_);
  nor (_03712_, _03711_, _03709_);
  and (_03713_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_03714_, _03713_, _00319_);
  nor (_03715_, _03714_, _03712_);
  nand (_03717_, _03715_, _03707_);
  and (_03719_, _01121_, _00319_);
  not (_03720_, _03719_);
  nand (_03721_, _03720_, _03717_);
  nand (_03722_, _00473_, _03706_);
  nor (_03723_, _24562_, _23210_);
  nor (_03724_, _03723_, _02580_);
  nor (_03725_, _03724_, _03711_);
  and (_03727_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_03728_, _03727_, _03725_);
  and (_03729_, _03728_, _00320_);
  and (_03730_, _03729_, _03722_);
  and (_03731_, _01061_, _00319_);
  nor (_03732_, _03731_, _03730_);
  nand (_03733_, _03732_, _03721_);
  or (_03734_, _03732_, _03721_);
  nand (_03735_, _03734_, _03733_);
  nand (_03736_, _26570_, _03706_);
  nor (_03737_, _24577_, _23291_);
  nor (_03738_, _03737_, _02599_);
  nor (_03739_, _03738_, _03711_);
  and (_03740_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03742_, _03740_, _00319_);
  nor (_03743_, _03742_, _03739_);
  nand (_03744_, _03743_, _03736_);
  or (_03745_, _00939_, _00320_);
  and (_03746_, _03745_, _03744_);
  nand (_03747_, _00393_, _03706_);
  nor (_03748_, _24177_, _23260_);
  nor (_03750_, _03748_, _02590_);
  nor (_03751_, _03750_, _03711_);
  and (_03752_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03754_, _03752_, _00319_);
  nor (_03755_, _03754_, _03751_);
  nand (_03756_, _03755_, _03747_);
  and (_03757_, _01009_, _00319_);
  not (_03758_, _03757_);
  nand (_03759_, _03758_, _03756_);
  nand (_03760_, _03759_, _03746_);
  or (_03762_, _03759_, _03746_);
  nand (_03763_, _03762_, _03760_);
  nand (_03764_, _03763_, _03735_);
  or (_03765_, _03763_, _03735_);
  nand (_03767_, _03765_, _03764_);
  nand (_03769_, _00654_, _03706_);
  nor (_03770_, _24636_, _23145_);
  nor (_03771_, _03770_, _24637_);
  nor (_03772_, _03771_, _03711_);
  and (_03773_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_03774_, _03773_, _00319_);
  nor (_03775_, _03774_, _03772_);
  nand (_03776_, _03775_, _03769_);
  and (_03777_, _01192_, _00319_);
  not (_03778_, _03777_);
  and (_03779_, _03778_, _03776_);
  nand (_03781_, _00747_, _03706_);
  nand (_03782_, _24607_, _23504_);
  or (_03783_, _24607_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_03784_, _03783_, _03710_);
  and (_03785_, _03784_, _03782_);
  and (_03786_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_03787_, _03786_, _00319_);
  nor (_03788_, _03787_, _03785_);
  nand (_03789_, _03788_, _03781_);
  and (_03790_, _01281_, _00319_);
  not (_03791_, _03790_);
  and (_03792_, _03791_, _03789_);
  or (_03793_, _03792_, _03779_);
  nand (_03794_, _03792_, _03779_);
  nand (_03795_, _03794_, _03793_);
  or (_03796_, _00813_, _00325_);
  not (_03797_, _24594_);
  nor (_03798_, _03797_, _23504_);
  nor (_03799_, _24594_, _23074_);
  nor (_03801_, _03799_, _03798_);
  nor (_03802_, _03801_, _03711_);
  and (_03803_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_03805_, _03803_, _00319_);
  nor (_03806_, _03805_, _03802_);
  and (_03807_, _03806_, _03796_);
  and (_03808_, _01353_, _00319_);
  or (_03809_, _03808_, _03807_);
  and (_03810_, _00883_, _03706_);
  nor (_03811_, _25481_, _23034_);
  or (_03813_, _03811_, _25482_);
  and (_03814_, _03813_, _03710_);
  and (_03815_, _00331_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_03816_, _03815_, _00319_);
  or (_03818_, _03816_, _03814_);
  or (_03819_, _03818_, _03810_);
  nor (_03821_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_03822_, _23003_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_03823_, _03822_, _03821_);
  nor (_03824_, _03823_, _01319_);
  and (_03825_, _03823_, _01319_);
  or (_03826_, _03825_, _03824_);
  and (_03828_, _03826_, _23390_);
  or (_03829_, _26539_, _26501_);
  and (_03830_, _03829_, _26540_);
  and (_03831_, _03830_, _23531_);
  and (_03832_, _01259_, _23120_);
  and (_03833_, _03832_, _23086_);
  nor (_03834_, _03833_, _01329_);
  or (_03835_, _03834_, _01341_);
  or (_03837_, _03835_, _23049_);
  nand (_03838_, _03835_, _23049_);
  and (_03839_, _03838_, _23514_);
  and (_03840_, _03839_, _03837_);
  and (_03841_, _23364_, _23050_);
  or (_03842_, _03841_, _23472_);
  and (_03843_, _03842_, _23506_);
  and (_03844_, _23488_, _23563_);
  and (_03845_, _23484_, _23050_);
  and (_03846_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  or (_03847_, _03846_, _03845_);
  or (_03849_, _03847_, _03844_);
  or (_03850_, _03849_, _03843_);
  or (_03851_, _03850_, _03840_);
  or (_03852_, _03851_, _03831_);
  or (_03853_, _03852_, _03828_);
  or (_03855_, _03853_, _00320_);
  and (_03857_, _03855_, _03819_);
  or (_03858_, _03857_, _03809_);
  nand (_03859_, _03857_, _03809_);
  and (_03860_, _03859_, _03858_);
  nand (_03861_, _03860_, _03795_);
  or (_03862_, _03860_, _03795_);
  nand (_03863_, _03862_, _03861_);
  nand (_03865_, _03863_, _03767_);
  or (_03866_, _03863_, _03767_);
  nand (_03868_, _03866_, _03865_);
  nand (_03869_, _03868_, _00228_);
  and (_03870_, _00191_, _00171_);
  or (_03871_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03872_, _03871_, _03870_);
  and (_03873_, _03872_, _03869_);
  not (_03874_, _00228_);
  not (_03875_, _00191_);
  and (_03876_, _03875_, _00171_);
  and (_03877_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor (_03878_, _00191_, _00171_);
  and (_03879_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_03880_, _03879_, _03877_);
  and (_03881_, _03880_, _03874_);
  not (_03882_, _00171_);
  and (_03883_, _00191_, _03882_);
  nor (_03884_, _00228_, _00546_);
  and (_03885_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03886_, _03885_, _03884_);
  and (_03887_, _03886_, _03883_);
  and (_03888_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03889_, _03878_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_03890_, _03889_, _03888_);
  and (_03891_, _03890_, _00228_);
  or (_03892_, _03891_, _03887_);
  or (_03893_, _03892_, _03881_);
  or (_03894_, _03893_, _03873_);
  and (_03895_, _03894_, _03705_);
  and (_03896_, _00051_, _00090_);
  and (_03897_, _00027_, _00143_);
  and (_03898_, _03897_, _26816_);
  and (_03899_, _23818_, _23824_);
  or (_03901_, _23815_, _26723_);
  nor (_03902_, _03901_, _03899_);
  not (_03903_, _26732_);
  not (_03904_, _23826_);
  not (_03905_, _26699_);
  and (_03906_, _23838_, _23810_);
  nor (_03908_, _03906_, _03905_);
  and (_03909_, _03908_, _03904_);
  and (_03910_, _03909_, _03903_);
  and (_03911_, _03910_, _03902_);
  and (_03912_, _26720_, _23834_);
  and (_03913_, _03912_, _03911_);
  or (_03914_, _23806_, _23801_);
  and (_03915_, _03914_, _23824_);
  not (_03916_, _03915_);
  nor (_03917_, _26757_, _23840_);
  not (_03919_, _03917_);
  nor (_03920_, _03919_, _26735_);
  and (_03922_, _03920_, _03916_);
  and (_03923_, _03922_, _26745_);
  and (_03925_, _03923_, _03913_);
  nor (_03926_, _03925_, _24279_);
  nor (_03927_, _03926_, p0_in[0]);
  and (_03928_, _03926_, _25360_);
  nor (_03929_, _03928_, _03927_);
  or (_03930_, _03929_, _03874_);
  nor (_03931_, _03926_, p0_in[4]);
  and (_03933_, _03926_, _25409_);
  nor (_03934_, _03933_, _03931_);
  or (_03935_, _03934_, _00228_);
  and (_03936_, _03935_, _03870_);
  and (_03937_, _03936_, _03930_);
  nor (_03938_, _03926_, p0_in[3]);
  not (_03939_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_03940_, _03926_, _03939_);
  nor (_03941_, _03940_, _03938_);
  or (_03942_, _03941_, _03874_);
  nor (_03943_, _03926_, p0_in[7]);
  not (_03944_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_03945_, _03926_, _03944_);
  nor (_03946_, _03945_, _03943_);
  or (_03947_, _03946_, _00228_);
  and (_03949_, _03947_, _03878_);
  and (_03950_, _03949_, _03942_);
  or (_03951_, _03950_, _03937_);
  nor (_03952_, _03926_, p0_in[1]);
  and (_03953_, _03926_, _25347_);
  nor (_03954_, _03953_, _03952_);
  or (_03955_, _03954_, _03874_);
  or (_03956_, _03926_, p0_in[5]);
  not (_03957_, _03926_);
  or (_03958_, _03957_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03959_, _03958_, _03956_);
  or (_03960_, _03959_, _00228_);
  and (_03962_, _03960_, _03876_);
  and (_03963_, _03962_, _03955_);
  nor (_03964_, _03926_, p0_in[2]);
  and (_03965_, _03926_, _25333_);
  nor (_03966_, _03965_, _03964_);
  or (_03967_, _03966_, _03874_);
  nor (_03968_, _03926_, p0_in[6]);
  and (_03970_, _03926_, _25392_);
  nor (_03972_, _03970_, _03968_);
  or (_03973_, _03972_, _00228_);
  and (_03975_, _03973_, _03883_);
  and (_03976_, _03975_, _03967_);
  or (_03977_, _03976_, _03963_);
  or (_03978_, _03977_, _03951_);
  and (_03979_, _03978_, _03898_);
  nor (_03980_, _03926_, p1_in[0]);
  and (_03981_, _03926_, _25277_);
  nor (_03982_, _03981_, _03980_);
  or (_03983_, _03982_, _03874_);
  nor (_03984_, _03926_, p1_in[4]);
  not (_03985_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03987_, _03926_, _03985_);
  nor (_03988_, _03987_, _03984_);
  or (_03990_, _03988_, _00228_);
  and (_03991_, _03990_, _03870_);
  and (_03993_, _03991_, _03983_);
  nor (_03995_, _03926_, p1_in[3]);
  and (_03996_, _03926_, _25234_);
  nor (_03997_, _03996_, _03995_);
  or (_03998_, _03997_, _03874_);
  nor (_04000_, _03926_, p1_in[7]);
  not (_04001_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_04003_, _03926_, _04001_);
  nor (_04004_, _04003_, _04000_);
  or (_04006_, _04004_, _00228_);
  and (_04008_, _04006_, _03878_);
  and (_04009_, _04008_, _03998_);
  or (_04011_, _04009_, _03993_);
  nor (_04012_, _03926_, p1_in[1]);
  and (_04014_, _03926_, _25263_);
  nor (_04016_, _04014_, _04012_);
  or (_04017_, _04016_, _03874_);
  or (_04018_, _03926_, p1_in[5]);
  or (_04019_, _03957_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_04020_, _04019_, _04018_);
  or (_04021_, _04020_, _00228_);
  and (_04022_, _04021_, _03876_);
  and (_04023_, _04022_, _04017_);
  nor (_04024_, _03926_, p1_in[2]);
  and (_04025_, _03926_, _25250_);
  nor (_04027_, _04025_, _04024_);
  or (_04028_, _04027_, _03874_);
  nor (_04029_, _03926_, p1_in[6]);
  and (_04030_, _03926_, _25295_);
  nor (_04031_, _04030_, _04029_);
  or (_04032_, _04031_, _00228_);
  and (_04033_, _04032_, _03883_);
  and (_04034_, _04033_, _04028_);
  or (_04035_, _04034_, _04023_);
  or (_04036_, _04035_, _04011_);
  and (_04038_, _04036_, _03703_);
  not (_04039_, _26816_);
  and (_04041_, _03702_, _04039_);
  and (_04042_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor (_04043_, _00228_, _02660_);
  or (_04045_, _04043_, _04042_);
  and (_04047_, _04045_, _03878_);
  nor (_04048_, _00228_, _02674_);
  and (_04049_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or (_04051_, _04049_, _04048_);
  and (_04052_, _04051_, _03883_);
  or (_04053_, _04052_, _04047_);
  and (_04054_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  not (_04056_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_04057_, _00228_, _04056_);
  or (_04058_, _04057_, _04054_);
  and (_04059_, _04058_, _03870_);
  and (_04060_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor (_04061_, _00228_, _02604_);
  or (_04062_, _04061_, _04060_);
  and (_04063_, _04062_, _03876_);
  or (_04064_, _04063_, _04059_);
  or (_04065_, _04064_, _04053_);
  and (_04066_, _04065_, _04041_);
  or (_04067_, _04066_, _04038_);
  or (_04069_, _04067_, _03979_);
  and (_04070_, _04069_, _03896_);
  and (_04071_, _03897_, _04039_);
  and (_04073_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_04074_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_04076_, _04074_, _04073_);
  and (_04078_, _04076_, _03878_);
  or (_04079_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or (_04080_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_04081_, _04080_, _03870_);
  and (_04082_, _04081_, _04079_);
  or (_04083_, _04082_, _04078_);
  nor (_04084_, _00228_, _02243_);
  and (_04085_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_04086_, _04085_, _04084_);
  and (_04088_, _04086_, _03883_);
  or (_04090_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  not (_04091_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand (_04093_, _00228_, _04091_);
  and (_04094_, _04093_, _03876_);
  and (_04095_, _04094_, _04090_);
  or (_04096_, _04095_, _04088_);
  or (_04098_, _04096_, _04083_);
  and (_04099_, _04098_, _03896_);
  and (_04100_, _03698_, _00090_);
  and (_04102_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_04103_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_04104_, _04103_, _04102_);
  and (_04105_, _04104_, _03878_);
  or (_04106_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_04108_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_04110_, _04108_, _03870_);
  and (_04111_, _04110_, _04106_);
  or (_04113_, _04111_, _04105_);
  and (_04114_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_04115_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_04117_, _04115_, _04114_);
  and (_04118_, _04117_, _03883_);
  or (_04119_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_04120_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_04121_, _04120_, _03876_);
  and (_04122_, _04121_, _04119_);
  or (_04123_, _04122_, _04118_);
  or (_04124_, _04123_, _04113_);
  and (_04125_, _04124_, _04100_);
  or (_04127_, _04125_, _04099_);
  and (_04128_, _04127_, _04071_);
  nor (_04129_, _03926_, p3_in[0]);
  and (_04130_, _03926_, _25074_);
  nor (_04131_, _04130_, _04129_);
  or (_04132_, _04131_, _03874_);
  nor (_04133_, _03926_, p3_in[4]);
  not (_04134_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_04135_, _03926_, _04134_);
  nor (_04136_, _04135_, _04133_);
  or (_04138_, _04136_, _00228_);
  and (_04139_, _04138_, _03870_);
  and (_04140_, _04139_, _04132_);
  nor (_04141_, _03926_, p3_in[3]);
  and (_04142_, _03926_, _25033_);
  nor (_04143_, _04142_, _04141_);
  or (_04144_, _04143_, _03874_);
  nor (_04145_, _03926_, p3_in[7]);
  not (_04146_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_04147_, _03926_, _04146_);
  nor (_04148_, _04147_, _04145_);
  or (_04149_, _04148_, _00228_);
  and (_04150_, _04149_, _03878_);
  and (_04151_, _04150_, _04144_);
  or (_04152_, _04151_, _04140_);
  nor (_04153_, _03926_, p3_in[1]);
  and (_04154_, _03926_, _25062_);
  nor (_04155_, _04154_, _04153_);
  or (_04156_, _04155_, _03874_);
  or (_04157_, _03926_, p3_in[5]);
  or (_04158_, _03957_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_04160_, _04158_, _04157_);
  or (_04161_, _04160_, _00228_);
  and (_04163_, _04161_, _03876_);
  and (_04164_, _04163_, _04156_);
  nor (_04166_, _03926_, p3_in[2]);
  and (_04167_, _03926_, _25049_);
  nor (_04169_, _04167_, _04166_);
  or (_04170_, _04169_, _03874_);
  nor (_04172_, _03926_, p3_in[6]);
  and (_04173_, _03926_, _25098_);
  nor (_04175_, _04173_, _04172_);
  or (_04176_, _04175_, _00228_);
  and (_04178_, _04176_, _03883_);
  and (_04179_, _04178_, _04170_);
  or (_04180_, _04179_, _04164_);
  or (_04181_, _04180_, _04152_);
  and (_04182_, _04181_, _03703_);
  nor (_04183_, _03926_, p2_in[0]);
  and (_04184_, _03926_, _25200_);
  nor (_04186_, _04184_, _04183_);
  or (_04188_, _04186_, _03874_);
  nor (_04190_, _03926_, p2_in[4]);
  and (_04192_, _03926_, _25160_);
  nor (_04193_, _04192_, _04190_);
  or (_04195_, _04193_, _00228_);
  and (_04196_, _04195_, _03870_);
  and (_04197_, _04196_, _04188_);
  nor (_04199_, _03926_, p2_in[3]);
  and (_04201_, _03926_, _25175_);
  nor (_04202_, _04201_, _04199_);
  or (_04203_, _04202_, _03874_);
  nor (_04204_, _03926_, p2_in[7]);
  not (_04206_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_04207_, _03926_, _04206_);
  nor (_04209_, _04207_, _04204_);
  or (_04210_, _04209_, _00228_);
  and (_04211_, _04210_, _03878_);
  and (_04212_, _04211_, _04203_);
  or (_04213_, _04212_, _04197_);
  nor (_04214_, _03926_, p2_in[1]);
  and (_04215_, _03926_, _25135_);
  nor (_04216_, _04215_, _04214_);
  or (_04217_, _04216_, _03874_);
  or (_04219_, _03926_, p2_in[5]);
  or (_04220_, _03957_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_04221_, _04220_, _04219_);
  or (_04222_, _04221_, _00228_);
  and (_04223_, _04222_, _03876_);
  and (_04224_, _04223_, _04217_);
  nor (_04225_, _03926_, p2_in[2]);
  and (_04226_, _03926_, _25188_);
  nor (_04227_, _04226_, _04225_);
  or (_04228_, _04227_, _03874_);
  nor (_04229_, _03926_, p2_in[6]);
  not (_04230_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_04231_, _03926_, _04230_);
  nor (_04232_, _04231_, _04229_);
  or (_04233_, _04232_, _00228_);
  and (_04234_, _04233_, _03883_);
  and (_04235_, _04234_, _04228_);
  or (_04236_, _04235_, _04224_);
  or (_04237_, _04236_, _04213_);
  and (_04238_, _04237_, _03898_);
  or (_04239_, _04238_, _04182_);
  and (_04240_, _04239_, _04100_);
  nor (_04241_, _00051_, _00090_);
  and (_04242_, _04241_, _03898_);
  and (_04243_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_04244_, _00228_, _23109_);
  or (_04245_, _04244_, _04243_);
  and (_04246_, _04245_, _03876_);
  nand (_04247_, _00228_, _23210_);
  or (_04248_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_04249_, _04248_, _03883_);
  and (_04250_, _04249_, _04247_);
  nor (_04251_, _00228_, _23034_);
  and (_04252_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_04253_, _04252_, _04251_);
  and (_04255_, _04253_, _03878_);
  or (_04256_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_04257_, _00228_, _23291_);
  and (_04258_, _04257_, _03870_);
  and (_04259_, _04258_, _04256_);
  or (_04260_, _04259_, _04255_);
  or (_04261_, _04260_, _04250_);
  or (_04263_, _04261_, _04246_);
  and (_04264_, _04263_, _04242_);
  nand (_04265_, _00143_, _00090_);
  or (_04266_, _04265_, _26816_);
  not (_04267_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_04268_, _03703_, _04267_);
  and (_04270_, _04268_, _04266_);
  and (_04272_, _04071_, _03699_);
  not (_04274_, _03699_);
  and (_04275_, _03898_, _04274_);
  nor (_04276_, _04275_, _04272_);
  and (_04277_, _04276_, _04270_);
  and (_04278_, _04100_, _04041_);
  or (_04280_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand (_04281_, _00228_, _24789_);
  and (_04283_, _04281_, _03878_);
  and (_04285_, _04283_, _04280_);
  and (_04286_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_04287_, _00228_, _24786_);
  or (_04288_, _04287_, _04286_);
  and (_04289_, _04288_, _03876_);
  or (_04290_, _04289_, _04285_);
  and (_04291_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor (_04292_, _00228_, _24784_);
  or (_04293_, _04292_, _04291_);
  and (_04295_, _04293_, _03870_);
  nand (_04297_, _00228_, _24800_);
  or (_04298_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_04300_, _04298_, _03883_);
  and (_04301_, _04300_, _04297_);
  or (_04302_, _04301_, _04295_);
  or (_04303_, _04302_, _04290_);
  and (_04304_, _04303_, _04278_);
  and (_04305_, _04241_, _03703_);
  and (_04306_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not (_04308_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor (_04309_, _00228_, _04308_);
  or (_04311_, _04309_, _04306_);
  and (_04312_, _04311_, _03878_);
  and (_04314_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  not (_04315_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor (_04317_, _00228_, _04315_);
  or (_04319_, _04317_, _04314_);
  and (_04320_, _04319_, _03876_);
  or (_04322_, _04320_, _04312_);
  and (_04323_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not (_04325_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor (_04326_, _00228_, _04325_);
  or (_04327_, _04326_, _04323_);
  and (_04328_, _04327_, _03870_);
  not (_04329_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor (_04330_, _00228_, _04329_);
  and (_04331_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_04332_, _04331_, _04330_);
  and (_04333_, _04332_, _03883_);
  or (_04334_, _04333_, _04328_);
  or (_04335_, _04334_, _04322_);
  and (_04336_, _04335_, _04305_);
  or (_04337_, _04336_, _04304_);
  or (_04338_, _04337_, _04277_);
  or (_04339_, _04338_, _04264_);
  and (_04340_, _00235_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_04341_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not (_04342_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_04343_, _00228_, _04342_);
  or (_04344_, _04343_, _04341_);
  and (_04345_, _04344_, _03876_);
  or (_04347_, _03874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_04348_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_04349_, _04348_, _03883_);
  and (_04350_, _04349_, _04347_);
  and (_04352_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_04353_, _00228_, _25483_);
  or (_04355_, _04353_, _04352_);
  and (_04356_, _04355_, _03878_);
  or (_04357_, _00228_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand (_04358_, _00228_, _25527_);
  and (_04360_, _04358_, _03870_);
  and (_04361_, _04360_, _04357_);
  or (_04362_, _04361_, _04356_);
  or (_04363_, _04362_, _04350_);
  or (_04364_, _04363_, _04345_);
  and (_04366_, _04364_, _04272_);
  or (_04367_, _04366_, _04340_);
  or (_04368_, _04367_, _04339_);
  or (_04370_, _04368_, _04240_);
  or (_04372_, _04370_, _04128_);
  or (_04373_, _04372_, _04070_);
  or (_04374_, _04373_, _03895_);
  and (_04375_, _04242_, _00322_);
  nor (_04376_, _04375_, _00151_);
  nand (_04377_, _04340_, _23504_);
  and (_04378_, _04377_, _04376_);
  and (_04379_, _04378_, _04374_);
  nor (_04380_, _00228_, _24043_);
  and (_04382_, _00228_, _02728_);
  or (_04383_, _04382_, _04380_);
  and (_04384_, _04383_, _03876_);
  or (_04385_, _00228_, _02450_);
  or (_04387_, _03874_, _23880_);
  and (_04388_, _04387_, _03883_);
  and (_04389_, _04388_, _04385_);
  nor (_04390_, _00228_, _23989_);
  and (_04392_, _00228_, _23577_);
  or (_04394_, _04392_, _04390_);
  and (_04395_, _04394_, _03878_);
  nand (_04396_, _00228_, _24210_);
  or (_04397_, _00228_, _02700_);
  and (_04399_, _04397_, _03870_);
  and (_04400_, _04399_, _04396_);
  or (_04401_, _04400_, _04395_);
  or (_04402_, _04401_, _04389_);
  nor (_04403_, _04402_, _04384_);
  nor (_04404_, _04403_, _04376_);
  or (_04405_, _04404_, _04379_);
  and (_27316_, _04405_, _22731_);
  and (_04406_, _24539_, _22844_);
  and (_04407_, _03878_, _03874_);
  not (_04409_, _04407_);
  and (_04410_, _04409_, _04406_);
  and (_04412_, _04410_, _00149_);
  not (_04413_, _00143_);
  nor (_04414_, _04413_, _00090_);
  and (_04416_, _00228_, _26816_);
  and (_04418_, _04416_, _03870_);
  nor (_04419_, _00051_, _03700_);
  and (_04420_, _04419_, _04418_);
  and (_04421_, _04420_, _04414_);
  and (_04423_, _04421_, _00322_);
  or (_04425_, _04423_, _00237_);
  or (_04426_, _04425_, _04412_);
  and (_04427_, _04421_, _00319_);
  and (_04428_, _00051_, _03700_);
  and (_04429_, _04428_, _04418_);
  and (_04430_, _04429_, _04414_);
  and (_04431_, _04430_, _00312_);
  and (_04433_, _00318_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_04434_, _03897_, _03896_);
  and (_04435_, _04434_, _03878_);
  and (_04436_, _04435_, _04416_);
  and (_04437_, _04436_, _04433_);
  or (_04438_, _04437_, _04431_);
  nor (_04439_, _04438_, _04427_);
  nor (_04440_, _04439_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_04441_, _04440_, _04426_);
  and (_04442_, _04434_, _03883_);
  and (_04443_, _04442_, _04416_);
  and (_04444_, _04443_, _04433_);
  nor (_04446_, _04444_, rst);
  and (_27317_, _04446_, _04441_);
  not (_04447_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_04448_, _03897_, _03699_);
  nor (_04449_, _00228_, _26816_);
  and (_04450_, _04449_, _03870_);
  and (_04451_, _04450_, _04448_);
  and (_04452_, _00228_, _04039_);
  and (_04454_, _04452_, _03870_);
  and (_04456_, _04454_, _04448_);
  nor (_04458_, _04456_, _04451_);
  and (_04459_, _04449_, _03876_);
  and (_04461_, _04459_, _04448_);
  and (_04462_, _04452_, _03883_);
  and (_04463_, _04462_, _04448_);
  nor (_04464_, _04463_, _04461_);
  and (_04465_, _04464_, _04458_);
  and (_04466_, _04454_, _04434_);
  and (_04467_, _04452_, _03878_);
  and (_04468_, _04467_, _04448_);
  nor (_04469_, _04468_, _04466_);
  and (_04470_, _04407_, _26816_);
  and (_04472_, _04100_, _03702_);
  and (_04474_, _04472_, _04470_);
  and (_04475_, _04100_, _03897_);
  and (_04476_, _04475_, _04454_);
  nor (_04477_, _04476_, _04474_);
  and (_04478_, _04477_, _04469_);
  and (_04479_, _04478_, _04465_);
  and (_04480_, _04467_, _04434_);
  and (_04481_, _04452_, _03876_);
  and (_04482_, _04481_, _04434_);
  nor (_04483_, _04482_, _04480_);
  and (_04484_, _04459_, _04434_);
  and (_04485_, _04462_, _04434_);
  nor (_04486_, _04485_, _04484_);
  and (_04488_, _04486_, _04483_);
  and (_04489_, _04470_, _04434_);
  and (_04491_, _04450_, _04434_);
  nor (_04493_, _04491_, _04489_);
  and (_04494_, _03896_, _03702_);
  and (_04495_, _04494_, _04454_);
  and (_04496_, _04481_, _04494_);
  nor (_04497_, _04496_, _04495_);
  and (_04498_, _04497_, _04493_);
  and (_04499_, _04498_, _04488_);
  and (_04500_, _04499_, _04479_);
  not (_04501_, _04418_);
  or (_04502_, _04501_, _04265_);
  and (_04503_, _04416_, _03878_);
  and (_04505_, _04503_, _04434_);
  nor (_04507_, _04443_, _04505_);
  and (_04508_, _04241_, _03702_);
  and (_04510_, _04508_, _04418_);
  and (_04512_, _04416_, _03876_);
  and (_04513_, _04512_, _04434_);
  nor (_04514_, _04513_, _04510_);
  and (_04516_, _04514_, _04507_);
  and (_04517_, _04516_, _04502_);
  nor (_04518_, _04430_, _04421_);
  and (_04519_, _04518_, _04517_);
  and (_04520_, _04519_, _04500_);
  nor (_04521_, _04520_, _04441_);
  nor (_04522_, _04521_, _04447_);
  not (_04523_, _04444_);
  nand (_04524_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_04526_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_04527_, _04526_, _04524_);
  nand (_04528_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nand (_04529_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_04530_, _04529_, _04528_);
  and (_04531_, _04530_, _04527_);
  nand (_04532_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand (_04533_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_04534_, _04533_, _04532_);
  nand (_04535_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nand (_04536_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_04537_, _04536_, _04535_);
  and (_04538_, _04537_, _04534_);
  and (_04539_, _04538_, _04531_);
  nand (_04540_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nand (_04541_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_04542_, _04541_, _04540_);
  nand (_04543_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_04544_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_04545_, _04544_, _04543_);
  and (_04547_, _04545_, _04542_);
  nand (_04548_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nand (_04549_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_04550_, _04549_, _04548_);
  nand (_04551_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_04552_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_04553_, _04552_, _04551_);
  and (_04554_, _04553_, _04550_);
  and (_04555_, _04554_, _04547_);
  and (_04556_, _04555_, _04539_);
  nand (_04557_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nand (_04558_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_04559_, _04558_, _04557_);
  nand (_04560_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_04561_, _04513_, _00105_);
  and (_04563_, _04561_, _04560_);
  and (_04564_, _04563_, _04559_);
  and (_04565_, _04475_, _04418_);
  nand (_04566_, _04565_, _04209_);
  and (_04567_, _04472_, _04418_);
  nand (_04568_, _04567_, _04148_);
  and (_04569_, _04568_, _04566_);
  and (_04570_, _04434_, _04418_);
  nand (_04572_, _04570_, _03946_);
  and (_04573_, _04494_, _04418_);
  nand (_04574_, _04573_, _04004_);
  and (_04575_, _04574_, _04572_);
  and (_04577_, _04575_, _04569_);
  and (_04578_, _04577_, _04564_);
  nand (_04579_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand (_04580_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_04581_, _04580_, _04579_);
  and (_04582_, _04581_, _04578_);
  and (_04583_, _04582_, _04556_);
  or (_04584_, _04583_, _04441_);
  nand (_04585_, _04584_, _04523_);
  or (_04586_, _04585_, _04522_);
  or (_04587_, _04523_, _00883_);
  and (_04589_, _04587_, _22731_);
  and (_27318_[7], _04589_, _04586_);
  and (_04590_, _03667_, _23583_);
  and (_04592_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_25237_, _04592_, _04590_);
  and (_04593_, _03667_, _23887_);
  and (_04594_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_25239_, _04594_, _04593_);
  and (_04595_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and (_04596_, _03662_, _23548_);
  or (_25245_, _04596_, _04595_);
  and (_04597_, _03667_, _23996_);
  and (_04598_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_25265_, _04598_, _04597_);
  and (_04599_, _03667_, _24134_);
  and (_04601_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_27228_, _04601_, _04599_);
  and (_04602_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and (_04603_, _03662_, _24134_);
  or (_25273_, _04603_, _04602_);
  and (_04604_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_04605_, _03662_, _24051_);
  or (_25282_, _04605_, _04604_);
  and (_04606_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and (_04607_, _03662_, _24089_);
  or (_27095_, _04607_, _04606_);
  and (_04608_, _02497_, _22974_);
  and (_04609_, _04608_, _23996_);
  not (_04610_, _04608_);
  and (_04611_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_25304_, _04611_, _04609_);
  and (_04612_, _04608_, _24134_);
  and (_04613_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_25317_, _04613_, _04612_);
  and (_04614_, _02512_, _24223_);
  not (_04615_, _04614_);
  and (_04616_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  and (_04617_, _04614_, _23887_);
  or (_25324_, _04617_, _04616_);
  and (_04619_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  and (_04620_, _04614_, _24089_);
  or (_25326_, _04620_, _04619_);
  and (_04622_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  and (_04623_, _04614_, _23583_);
  or (_25337_, _04623_, _04622_);
  and (_04625_, _03667_, _24219_);
  and (_04626_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_25348_, _04626_, _04625_);
  and (_04627_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  and (_04628_, _04614_, _24134_);
  or (_25373_, _04628_, _04627_);
  and (_04629_, _24219_, _24008_);
  and (_04630_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or (_25379_, _04630_, _04629_);
  and (_04631_, _04608_, _23548_);
  and (_04632_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_25389_, _04632_, _04631_);
  and (_04633_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  and (_04634_, _04614_, _23996_);
  or (_27094_, _04634_, _04633_);
  and (_04635_, _04608_, _24219_);
  and (_04636_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_25399_, _04636_, _04635_);
  and (_04637_, _04608_, _24089_);
  and (_04638_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_25427_, _04638_, _04637_);
  and (_04639_, _04608_, _23583_);
  and (_04640_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_27213_, _04640_, _04639_);
  and (_04641_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  and (_04642_, _04614_, _24219_);
  or (_25437_, _04642_, _04641_);
  and (_04643_, _04608_, _23887_);
  and (_04644_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_25439_, _04644_, _04643_);
  and (_04645_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  and (_04646_, _02836_, _23548_);
  or (_25452_, _04646_, _04645_);
  and (_04647_, _02497_, _24095_);
  and (_04648_, _04647_, _24134_);
  not (_04649_, _04647_);
  and (_04650_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_25464_, _04650_, _04648_);
  and (_04651_, _04647_, _24051_);
  and (_04652_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_25468_, _04652_, _04651_);
  and (_04653_, _02512_, _24095_);
  not (_04654_, _04653_);
  and (_04656_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_04657_, _04653_, _24219_);
  or (_25471_, _04657_, _04656_);
  and (_04658_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  and (_04659_, _03011_, _23996_);
  or (_25476_, _04659_, _04658_);
  and (_04660_, _04647_, _23996_);
  and (_04661_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_25498_, _04661_, _04660_);
  and (_04662_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and (_04663_, _04653_, _24089_);
  or (_27092_, _04663_, _04662_);
  and (_04665_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and (_04667_, _04653_, _23583_);
  or (_25525_, _04667_, _04665_);
  and (_04668_, _04647_, _23548_);
  and (_04669_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_25530_, _04669_, _04668_);
  and (_04670_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and (_04671_, _04653_, _23887_);
  or (_27091_, _04671_, _04670_);
  and (_04672_, _04647_, _24219_);
  and (_04673_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_25537_, _04673_, _04672_);
  and (_04674_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  and (_04675_, _03011_, _23583_);
  or (_25555_, _04675_, _04674_);
  and (_04676_, _04647_, _23583_);
  and (_04677_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_25559_, _04677_, _04676_);
  and (_04678_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  and (_04680_, _03011_, _23887_);
  or (_25562_, _04680_, _04678_);
  and (_04681_, _04647_, _23887_);
  and (_04682_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_25570_, _04682_, _04681_);
  not (_04683_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_04684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_04685_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor (_04686_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_04687_, _04686_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and (_04688_, _04687_, _04685_);
  and (_04689_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _02674_);
  or (_04690_, _04689_, _04688_);
  nor (_04691_, _04690_, _04684_);
  nand (_04692_, _04691_, _04683_);
  nor (_04693_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor (_04694_, _04693_, _04691_);
  nand (_04695_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_04696_, _04695_, _04694_);
  and (_04697_, _04696_, _22731_);
  and (_25638_, _04697_, _04692_);
  and (_04698_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  and (_04699_, _03011_, _24134_);
  or (_25641_, _04699_, _04698_);
  not (_04700_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and (_04701_, _02652_, _04700_);
  and (_04702_, _04701_, _02755_);
  and (_04703_, _04702_, _02752_);
  nand (_04704_, _04703_, _02648_);
  not (_04705_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_04706_, _02757_, _04705_);
  and (_04707_, _04706_, _04704_);
  or (_04708_, _04707_, _02658_);
  and (_25646_, _04708_, _22731_);
  and (_04709_, _02497_, _24372_);
  and (_04710_, _04709_, _24089_);
  not (_04711_, _04709_);
  and (_04712_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or (_25653_, _04712_, _04710_);
  and (_25655_, _04694_, _22731_);
  and (_04714_, _04709_, _23583_);
  and (_04715_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_25667_, _04715_, _04714_);
  and (_04716_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  and (_04718_, _03011_, _24051_);
  or (_25671_, _04718_, _04716_);
  and (_04719_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  and (_04721_, _03011_, _24089_);
  or (_25676_, _04721_, _04719_);
  and (_04722_, _02654_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  or (_04723_, _04722_, _02658_);
  nor (_04724_, _02675_, rst);
  and (_25678_, _04724_, _04723_);
  nand (_04725_, _02910_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or (_04726_, _02910_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_04727_, _04726_, _22731_);
  nand (_04729_, _04727_, _04725_);
  nor (_25680_, _04729_, _02658_);
  not (_04730_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_04732_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_04733_, _04687_, _04342_);
  or (_04735_, _04733_, _04689_);
  nor (_04736_, _04735_, _04732_);
  nand (_04737_, _04736_, _04730_);
  nor (_04738_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor (_04739_, _04738_, _04736_);
  nand (_04741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_04742_, _04741_, _04739_);
  and (_04743_, _04742_, _22731_);
  and (_25688_, _04743_, _04737_);
  and (_25690_, _04739_, _22731_);
  and (_04744_, _04709_, _23996_);
  and (_04745_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_27189_, _04745_, _04744_);
  and (_04747_, _04709_, _24134_);
  and (_04748_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_25702_, _04748_, _04747_);
  not (_04749_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor (_04750_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _04056_);
  not (_04751_, _04750_);
  nor (_04752_, _02568_, _02810_);
  and (_04753_, _04752_, _04751_);
  and (_04754_, _04753_, _02820_);
  nor (_04755_, _04754_, _04749_);
  and (_04756_, _04754_, rxd_i);
  or (_04757_, _04756_, rst);
  or (_25706_, _04757_, _04755_);
  or (_04758_, _02802_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_04759_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_04760_, _04759_, _02568_);
  or (_04761_, _04760_, _02778_);
  nand (_04762_, _04761_, _04758_);
  nand (_25708_, _04762_, _02080_);
  and (_04763_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and (_04764_, _04653_, _23996_);
  or (_25717_, _04764_, _04763_);
  and (_04766_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and (_04767_, _04653_, _24134_);
  or (_25725_, _04767_, _04766_);
  and (_04768_, _02497_, _24146_);
  and (_04769_, _04768_, _24134_);
  not (_04770_, _04768_);
  and (_04772_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_25731_, _04772_, _04769_);
  and (_04773_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and (_04774_, _04653_, _24051_);
  or (_25733_, _04774_, _04773_);
  and (_04775_, _04768_, _23996_);
  and (_04777_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_25742_, _04777_, _04775_);
  and (_04778_, _02502_, _23996_);
  and (_04779_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_25747_, _04779_, _04778_);
  and (_04781_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_04782_, _23687_);
  nor (_04783_, _26748_, _04782_);
  and (_04785_, _24257_, _23797_);
  or (_04786_, _04785_, _01985_);
  nor (_04787_, _23782_, _23749_);
  and (_04789_, _04787_, _23838_);
  or (_04790_, _04789_, _23897_);
  or (_04791_, _04790_, _04786_);
  or (_04792_, _04791_, _04783_);
  and (_04793_, _23784_, _23687_);
  or (_04794_, _01979_, _04793_);
  and (_04795_, _23911_, _23687_);
  or (_04796_, _03905_, _23841_);
  or (_04797_, _04796_, _04795_);
  nor (_04798_, _04797_, _04794_);
  nand (_04799_, _04798_, _26733_);
  and (_04800_, _23780_, _23772_);
  and (_04801_, _26730_, _23687_);
  or (_04802_, _04801_, _04800_);
  or (_04803_, _26757_, _24259_);
  and (_04804_, _04803_, _23791_);
  or (_04806_, _04804_, _04802_);
  or (_04807_, _04806_, _04799_);
  or (_04808_, _04807_, _04792_);
  and (_04809_, _04808_, _22737_);
  or (_04810_, _04809_, _04781_);
  and (_26847_[0], _04810_, _22731_);
  and (_04812_, _24408_, _23941_);
  and (_04813_, _04812_, _23996_);
  not (_04815_, _04812_);
  and (_04816_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_25762_, _04816_, _04813_);
  and (_04818_, _04812_, _24051_);
  and (_04819_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_25774_, _04819_, _04818_);
  and (_04820_, _04812_, _23583_);
  and (_04821_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_27138_, _04821_, _04820_);
  and (_04823_, _24134_, _22983_);
  and (_04824_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  or (_25847_, _04824_, _04823_);
  and (_04825_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and (_04826_, _03319_, _23548_);
  or (_25853_, _04826_, _04825_);
  and (_04827_, _04709_, _24219_);
  and (_04828_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_25857_, _04828_, _04827_);
  and (_04829_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and (_04830_, _03319_, _24219_);
  or (_25871_, _04830_, _04829_);
  and (_04831_, _24518_, _23583_);
  and (_04832_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  or (_25875_, _04832_, _04831_);
  and (_04833_, _02432_, _24219_);
  and (_04835_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  or (_25883_, _04835_, _04833_);
  and (_04837_, _04768_, _24219_);
  and (_04838_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_25887_, _04838_, _04837_);
  and (_04840_, _04768_, _23887_);
  and (_04841_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_25889_, _04841_, _04840_);
  and (_04843_, _04768_, _23548_);
  and (_04844_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_25904_, _04844_, _04843_);
  and (_04846_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_04847_, _03319_, _23887_);
  or (_25906_, _04847_, _04846_);
  and (_04848_, _03360_, _24219_);
  and (_04849_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or (_25927_, _04849_, _04848_);
  and (_04851_, _04768_, _23583_);
  and (_04852_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_27080_, _04852_, _04851_);
  and (_04853_, _02039_, _24140_);
  not (_04854_, _04853_);
  and (_04855_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  and (_04856_, _04853_, _23583_);
  or (_25939_, _04856_, _04855_);
  and (_04858_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  and (_04859_, _04853_, _23887_);
  or (_25946_, _04859_, _04858_);
  and (_04860_, _04768_, _24089_);
  and (_04861_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  or (_25949_, _04861_, _04860_);
  and (_04862_, _03360_, _23583_);
  and (_04864_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_25953_, _04864_, _04862_);
  and (_04865_, _03308_, _24056_);
  and (_04866_, _04865_, _24134_);
  not (_04867_, _04865_);
  and (_04868_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  or (_25957_, _04868_, _04866_);
  and (_04869_, _24518_, _24089_);
  and (_04871_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  or (_25960_, _04871_, _04869_);
  and (_04872_, _02432_, _24089_);
  and (_04874_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  or (_25966_, _04874_, _04872_);
  and (_04875_, _02432_, _23887_);
  and (_04876_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  or (_25972_, _04876_, _04875_);
  and (_04877_, _03360_, _24051_);
  and (_04878_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or (_25993_, _04878_, _04877_);
  and (_04879_, _02039_, _24319_);
  not (_04880_, _04879_);
  and (_04881_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_04882_, _04879_, _23548_);
  or (_25996_, _04882_, _04881_);
  and (_04884_, _03313_, _23887_);
  and (_04885_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  or (_26004_, _04885_, _04884_);
  and (_04886_, _03313_, _24134_);
  and (_04887_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  or (_26009_, _04887_, _04886_);
  and (_04888_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_04890_, _04879_, _23887_);
  or (_26012_, _04890_, _04888_);
  and (_04891_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_04892_, _04879_, _24089_);
  or (_26015_, _04892_, _04891_);
  and (_04893_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_04894_, _04879_, _24051_);
  or (_26019_, _04894_, _04893_);
  and (_04895_, _03313_, _24051_);
  and (_04896_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  or (_26026_, _04896_, _04895_);
  and (_04897_, _02039_, _24146_);
  not (_04898_, _04897_);
  and (_04899_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_04900_, _04897_, _24089_);
  or (_26029_, _04900_, _04899_);
  and (_04901_, _03033_, _23548_);
  and (_04902_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_26030_, _04902_, _04901_);
  and (_04903_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_04904_, _04897_, _24134_);
  or (_26033_, _04904_, _04903_);
  and (_04905_, _02039_, _24372_);
  not (_04907_, _04905_);
  and (_04908_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_04909_, _04905_, _23548_);
  or (_27010_, _04909_, _04908_);
  and (_04910_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_04912_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_04913_, _22740_, _04912_);
  or (_04915_, _04913_, _04910_);
  and (_26862_[15], _04915_, _22731_);
  and (_04916_, _03033_, _23583_);
  and (_04918_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or (_26046_, _04918_, _04916_);
  and (_04920_, _24301_, _24236_);
  and (_04921_, _04920_, _24051_);
  not (_04923_, _04920_);
  and (_04924_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_26052_, _04924_, _04921_);
  and (_04925_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_04926_, _04905_, _23583_);
  or (_26056_, _04926_, _04925_);
  and (_04928_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_04930_, _04905_, _24051_);
  or (_26062_, _04930_, _04928_);
  and (_04932_, _25672_, _23548_);
  and (_04933_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_26065_, _04933_, _04932_);
  and (_04935_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_04936_, _04905_, _23996_);
  or (_26069_, _04936_, _04935_);
  and (_04937_, _02039_, _24095_);
  not (_04938_, _04937_);
  and (_04939_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  and (_04940_, _04937_, _24219_);
  or (_27012_, _04940_, _04939_);
  and (_04941_, _03033_, _24219_);
  and (_04942_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_26075_, _04942_, _04941_);
  and (_04943_, _03001_, _24134_);
  and (_04944_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_26078_, _04944_, _04943_);
  and (_04946_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  and (_04947_, _04937_, _23887_);
  or (_26086_, _04947_, _04946_);
  and (_04948_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  and (_04949_, _04937_, _24089_);
  or (_26096_, _04949_, _04948_);
  and (_04950_, _25413_, _22974_);
  and (_04951_, _04950_, _24089_);
  not (_04952_, _04950_);
  and (_04953_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  or (_26105_, _04953_, _04951_);
  or (_04955_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_04956_, _04955_, _22731_);
  nand (_04957_, _02071_, _24082_);
  and (_26109_, _04957_, _04956_);
  nor (_27315_[0], \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_04959_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor (_04961_, _03689_, rst);
  and (_27315_[1], _04961_, _04959_);
  nor (_04964_, _03689_, _03688_);
  or (_04965_, _04964_, _03690_);
  and (_04967_, _03693_, _22731_);
  and (_27315_[2], _04967_, _04965_);
  and (_04969_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  and (_04970_, _04937_, _24134_);
  or (_26117_, _04970_, _04969_);
  nand (_04971_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_04973_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_04974_, _04973_, _04971_);
  nand (_04975_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_04976_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_04977_, _04976_, _04975_);
  and (_04978_, _04977_, _04974_);
  nand (_04979_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_04980_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_04981_, _04980_, _04979_);
  nand (_04982_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nand (_04983_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_04984_, _04983_, _04982_);
  and (_04985_, _04984_, _04981_);
  and (_04986_, _04985_, _04978_);
  nand (_04987_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand (_04988_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_04989_, _04988_, _04987_);
  nand (_04990_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_04991_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_04992_, _04991_, _04990_);
  and (_04993_, _04992_, _04989_);
  nand (_04994_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  nand (_04995_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_04996_, _04995_, _04994_);
  nand (_04997_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand (_04998_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_04999_, _04998_, _04997_);
  and (_05000_, _04999_, _04996_);
  and (_05001_, _05000_, _04993_);
  and (_05002_, _05001_, _04986_);
  nand (_05003_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand (_05004_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_05006_, _05004_, _05003_);
  nand (_05007_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not (_05008_, _00187_);
  nand (_05009_, _04513_, _05008_);
  and (_05010_, _05009_, _05007_);
  and (_05011_, _05010_, _05006_);
  nand (_05012_, _04565_, _04186_);
  nand (_05013_, _04567_, _04131_);
  and (_05014_, _05013_, _05012_);
  nand (_05015_, _04570_, _03929_);
  nand (_05016_, _04573_, _03982_);
  and (_05017_, _05016_, _05015_);
  and (_05018_, _05017_, _05014_);
  and (_05020_, _05018_, _05011_);
  not (_05021_, _04430_);
  or (_05022_, _05021_, _03868_);
  nand (_05023_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_05025_, _05023_, _05022_);
  and (_05026_, _05025_, _05020_);
  and (_05028_, _05026_, _05002_);
  nor (_05030_, _05028_, _04441_);
  not (_05031_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nor (_05032_, _04521_, _05031_);
  or (_05033_, _05032_, _04444_);
  or (_05034_, _05033_, _05030_);
  or (_05035_, _04523_, _26570_);
  and (_05036_, _05035_, _22731_);
  and (_27318_[0], _05036_, _05034_);
  not (_05037_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nor (_05038_, _04521_, _05037_);
  nand (_05039_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_05040_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_05041_, _05040_, _05039_);
  nand (_05042_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_05043_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_05044_, _05043_, _05042_);
  and (_05045_, _05044_, _05041_);
  nand (_05046_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_05047_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_05048_, _05047_, _05046_);
  nand (_05049_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_05050_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_05051_, _05050_, _05049_);
  and (_05053_, _05051_, _05048_);
  and (_05054_, _05053_, _05045_);
  nand (_05055_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand (_05056_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_05057_, _05056_, _05055_);
  nand (_05058_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nand (_05059_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_05060_, _05059_, _05058_);
  and (_05061_, _05060_, _05057_);
  nand (_05062_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  nand (_05063_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_05065_, _05063_, _05062_);
  nand (_05066_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_05067_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_05068_, _05067_, _05066_);
  and (_05069_, _05068_, _05065_);
  and (_05070_, _05069_, _05061_);
  and (_05071_, _05070_, _05054_);
  nand (_05072_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nand (_05073_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_05074_, _05073_, _05072_);
  nand (_05075_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_05076_, _04513_, _00167_);
  and (_05077_, _05076_, _05075_);
  and (_05078_, _05077_, _05074_);
  nand (_05079_, _04565_, _04216_);
  nand (_05080_, _04567_, _04155_);
  and (_05081_, _05080_, _05079_);
  nand (_05082_, _04570_, _03954_);
  nand (_05083_, _04573_, _04016_);
  and (_05084_, _05083_, _05082_);
  and (_05085_, _05084_, _05081_);
  and (_05086_, _05085_, _05078_);
  nand (_05087_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nand (_05088_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_05090_, _05088_, _05087_);
  and (_05092_, _05090_, _05086_);
  and (_05094_, _05092_, _05071_);
  nor (_05095_, _05094_, _04441_);
  or (_05096_, _05095_, _04444_);
  or (_05097_, _05096_, _05038_);
  or (_05098_, _04523_, _00393_);
  and (_05099_, _05098_, _22731_);
  and (_27318_[1], _05099_, _05097_);
  not (_05100_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nor (_05101_, _04521_, _05100_);
  nand (_05102_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nand (_05103_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and (_05104_, _05103_, _05102_);
  nand (_05105_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  nand (_05106_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_05107_, _05106_, _05105_);
  and (_05108_, _05107_, _05104_);
  nand (_05109_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand (_05110_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_05111_, _05110_, _05109_);
  nand (_05112_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand (_05114_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_05115_, _05114_, _05112_);
  and (_05117_, _05115_, _05111_);
  and (_05118_, _05117_, _05108_);
  nand (_05119_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand (_05120_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_05121_, _05120_, _05119_);
  nand (_05122_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nand (_05123_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_05124_, _05123_, _05122_);
  and (_05125_, _05124_, _05121_);
  nand (_05126_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand (_05127_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_05128_, _05127_, _05126_);
  nand (_05129_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand (_05130_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_05131_, _05130_, _05129_);
  and (_05132_, _05131_, _05128_);
  and (_05133_, _05132_, _05125_);
  and (_05134_, _05133_, _05118_);
  nand (_05136_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nand (_05137_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_05138_, _05137_, _05136_);
  nand (_05139_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_05140_, _04513_, _00205_);
  and (_05141_, _05140_, _05139_);
  and (_05142_, _05141_, _05138_);
  nand (_05144_, _04565_, _04227_);
  nand (_05145_, _04567_, _04169_);
  and (_05146_, _05145_, _05144_);
  nand (_05147_, _04573_, _04027_);
  nand (_05148_, _04570_, _03966_);
  and (_05149_, _05148_, _05147_);
  and (_05150_, _05149_, _05146_);
  and (_05151_, _05150_, _05142_);
  nand (_05152_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nand (_05153_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_05155_, _05153_, _05152_);
  and (_05156_, _05155_, _05151_);
  and (_05157_, _05156_, _05134_);
  or (_05158_, _05157_, _04441_);
  nand (_05159_, _05158_, _04523_);
  or (_05160_, _05159_, _05101_);
  or (_05161_, _04523_, _00473_);
  and (_05162_, _05161_, _22731_);
  and (_27318_[2], _05162_, _05160_);
  not (_05164_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nor (_05165_, _04521_, _05164_);
  nand (_05167_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  nand (_05169_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_05170_, _05169_, _05167_);
  nand (_05171_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_05173_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_05174_, _05173_, _05171_);
  and (_05176_, _05174_, _05170_);
  nand (_05177_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand (_05178_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_05179_, _05178_, _05177_);
  nand (_05180_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_05181_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_05182_, _05181_, _05180_);
  and (_05183_, _05182_, _05179_);
  and (_05184_, _05183_, _05176_);
  nand (_05185_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nand (_05186_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_05188_, _05186_, _05185_);
  nand (_05190_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nand (_05191_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_05192_, _05191_, _05190_);
  and (_05193_, _05192_, _05188_);
  nand (_05194_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand (_05195_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_05196_, _05195_, _05194_);
  nand (_05197_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nand (_05198_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_05199_, _05198_, _05197_);
  and (_05200_, _05199_, _05196_);
  and (_05201_, _05200_, _05193_);
  and (_05202_, _05201_, _05184_);
  nand (_05203_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nand (_05204_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_05205_, _05204_, _05203_);
  nand (_05207_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_05208_, _04513_, _26805_);
  and (_05209_, _05208_, _05207_);
  and (_05210_, _05209_, _05205_);
  nand (_05211_, _04565_, _04202_);
  nand (_05212_, _04567_, _04143_);
  and (_05213_, _05212_, _05211_);
  nand (_05214_, _04573_, _03997_);
  nand (_05215_, _04570_, _03941_);
  and (_05216_, _05215_, _05214_);
  and (_05218_, _05216_, _05213_);
  and (_05219_, _05218_, _05210_);
  nand (_05221_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand (_05223_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_05224_, _05223_, _05221_);
  and (_05225_, _05224_, _05219_);
  and (_05226_, _05225_, _05202_);
  or (_05227_, _05226_, _04441_);
  nand (_05228_, _05227_, _04523_);
  or (_05229_, _05228_, _05165_);
  or (_05230_, _04523_, _00569_);
  and (_05231_, _05230_, _22731_);
  and (_27318_[3], _05231_, _05229_);
  not (_05232_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nor (_05233_, _04521_, _05232_);
  nand (_05234_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  nand (_05235_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_05236_, _05235_, _05234_);
  nand (_05237_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  nand (_05239_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_05240_, _05239_, _05237_);
  and (_05242_, _05240_, _05236_);
  nand (_05243_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nand (_05244_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_05246_, _05244_, _05243_);
  nand (_05247_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_05248_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_05249_, _05248_, _05247_);
  and (_05250_, _05249_, _05246_);
  and (_05251_, _05250_, _05242_);
  nand (_05253_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nand (_05254_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_05255_, _05254_, _05253_);
  nand (_05256_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand (_05257_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_05258_, _05257_, _05256_);
  and (_05259_, _05258_, _05255_);
  nand (_05260_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand (_05261_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_05262_, _05261_, _05260_);
  nand (_05263_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand (_05264_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_05265_, _05264_, _05263_);
  and (_05266_, _05265_, _05262_);
  and (_05267_, _05266_, _05259_);
  and (_05268_, _05267_, _05251_);
  nand (_05269_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_05270_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_05271_, _05270_, _05269_);
  nand (_05273_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_05274_, _00014_);
  nand (_05275_, _04513_, _05274_);
  and (_05276_, _05275_, _05273_);
  and (_05277_, _05276_, _05271_);
  nand (_05278_, _04565_, _04193_);
  nand (_05279_, _04567_, _04136_);
  and (_05280_, _05279_, _05278_);
  nand (_05281_, _04573_, _03988_);
  nand (_05282_, _04570_, _03934_);
  and (_05284_, _05282_, _05281_);
  and (_05285_, _05284_, _05280_);
  and (_05286_, _05285_, _05277_);
  nand (_05287_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nand (_05288_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_05289_, _05288_, _05287_);
  and (_05291_, _05289_, _05286_);
  and (_05292_, _05291_, _05268_);
  or (_05293_, _05292_, _04441_);
  nand (_05294_, _05293_, _04523_);
  or (_05295_, _05294_, _05233_);
  or (_05296_, _04523_, _00654_);
  and (_05297_, _05296_, _22731_);
  and (_27318_[4], _05297_, _05295_);
  not (_05298_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_05299_, _04426_, _05298_);
  and (_05300_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_05301_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_05302_, _05301_, _05300_);
  and (_05304_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_05305_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or (_05306_, _05305_, _05304_);
  or (_05307_, _05306_, _05302_);
  and (_05308_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_05309_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_05310_, _05309_, _05308_);
  and (_05311_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_05312_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_05313_, _05312_, _05311_);
  or (_05314_, _05313_, _05310_);
  or (_05315_, _05314_, _05307_);
  and (_05316_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_05317_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_05318_, _05317_, _05316_);
  and (_05319_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_05321_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_05322_, _05321_, _05319_);
  or (_05323_, _05322_, _05318_);
  and (_05324_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_05326_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_05327_, _05326_, _05324_);
  and (_05328_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_05329_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_05331_, _05329_, _05328_);
  or (_05332_, _05331_, _05327_);
  or (_05333_, _05332_, _05323_);
  or (_05334_, _05333_, _05315_);
  and (_05335_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_05337_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_05338_, _05337_, _05335_);
  and (_05339_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_05340_, _00046_);
  and (_05341_, _04513_, _05340_);
  or (_05342_, _05341_, _05339_);
  or (_05343_, _05342_, _05338_);
  and (_05344_, _04565_, _04221_);
  and (_05345_, _04567_, _04160_);
  or (_05347_, _05345_, _05344_);
  and (_05348_, _04570_, _03959_);
  and (_05349_, _04573_, _04020_);
  or (_05350_, _05349_, _05348_);
  or (_05351_, _05350_, _05347_);
  or (_05352_, _05351_, _05343_);
  and (_05353_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_05355_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_05356_, _05355_, _05353_);
  or (_05358_, _05356_, _05352_);
  nor (_05359_, _05358_, _05334_);
  nor (_05360_, _05359_, _04440_);
  nor (_05361_, _04521_, _05298_);
  or (_05362_, _05361_, _05360_);
  and (_05363_, _05362_, _05299_);
  or (_05364_, _05363_, _04444_);
  or (_05365_, _04523_, _00747_);
  and (_05366_, _05365_, _22731_);
  and (_27318_[5], _05366_, _05364_);
  not (_05367_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nor (_05368_, _04521_, _05367_);
  nand (_05370_, _04468_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nand (_05371_, _04466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_05372_, _05371_, _05370_);
  nand (_05373_, _04474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nand (_05374_, _04476_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_05375_, _05374_, _05373_);
  and (_05376_, _05375_, _05372_);
  nand (_05377_, _04451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand (_05378_, _04456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_05380_, _05378_, _05377_);
  nand (_05381_, _04461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nand (_05382_, _04463_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_05384_, _05382_, _05381_);
  and (_05385_, _05384_, _05380_);
  and (_05386_, _05385_, _05376_);
  nand (_05387_, _04489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  nand (_05388_, _04491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_05389_, _05388_, _05387_);
  nand (_05391_, _04496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  nand (_05392_, _04495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_05393_, _05392_, _05391_);
  and (_05394_, _05393_, _05389_);
  nand (_05395_, _04480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_05396_, _04482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_05397_, _05396_, _05395_);
  nand (_05398_, _04484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_05399_, _04485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_05400_, _05399_, _05398_);
  and (_05401_, _05400_, _05397_);
  and (_05402_, _05401_, _05394_);
  and (_05403_, _05402_, _05386_);
  nand (_05404_, _04505_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  nand (_05405_, _04443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_05406_, _05405_, _05404_);
  nand (_05407_, _04510_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  not (_05408_, _00084_);
  nand (_05409_, _04513_, _05408_);
  and (_05410_, _05409_, _05407_);
  and (_05411_, _05410_, _05406_);
  nand (_05412_, _04565_, _04232_);
  nand (_05413_, _04567_, _04175_);
  and (_05414_, _05413_, _05412_);
  nand (_05415_, _04570_, _03972_);
  nand (_05416_, _04573_, _04031_);
  and (_05417_, _05416_, _05415_);
  and (_05418_, _05417_, _05414_);
  and (_05419_, _05418_, _05411_);
  nand (_05420_, _04421_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand (_05421_, _04430_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_05422_, _05421_, _05420_);
  and (_05424_, _05422_, _05419_);
  and (_05425_, _05424_, _05403_);
  or (_05426_, _05425_, _04441_);
  nand (_05427_, _05426_, _04523_);
  or (_05428_, _05427_, _05368_);
  nand (_05429_, _04444_, _00813_);
  and (_05430_, _05429_, _22731_);
  and (_27318_[6], _05430_, _05428_);
  and (_05431_, _24474_, _24408_);
  and (_05432_, _05431_, _23583_);
  not (_05434_, _05431_);
  and (_05435_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  or (_26604_, _05435_, _05432_);
  and (_05436_, _05431_, _23548_);
  and (_05437_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  or (_26621_, _05437_, _05436_);
  and (_05438_, _24476_, _24349_);
  and (_05439_, _05438_, _24219_);
  not (_05440_, _05438_);
  and (_05441_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_27185_, _05441_, _05439_);
  and (_05442_, _24476_, _24159_);
  and (_05443_, _05442_, _23548_);
  not (_05444_, _05442_);
  and (_05446_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_26661_, _05446_, _05443_);
  and (_05448_, _02502_, _23583_);
  and (_05449_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  or (_26685_, _05449_, _05448_);
  and (_05451_, _02502_, _24089_);
  and (_05453_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or (_26725_, _05453_, _05451_);
  and (_05454_, _02502_, _23887_);
  and (_05455_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  or (_26728_, _05455_, _05454_);
  and (_05456_, _24408_, _24056_);
  and (_05457_, _05456_, _24134_);
  not (_05458_, _05456_);
  and (_05459_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_26746_, _05459_, _05457_);
  and (_05460_, _24140_, _24006_);
  and (_05461_, _05460_, _24219_);
  not (_05462_, _05460_);
  and (_05464_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or (_26771_, _05464_, _05461_);
  and (_05465_, _24297_, _23945_);
  and (_05467_, _05465_, _23887_);
  not (_05468_, _05465_);
  and (_05469_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  or (_26774_, _05469_, _05467_);
  and (_05471_, _05456_, _24089_);
  and (_05472_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_27126_, _05472_, _05471_);
  and (_05473_, _05456_, _23887_);
  and (_05475_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_26785_, _05475_, _05473_);
  and (_05478_, _24496_, _24349_);
  and (_05479_, _05478_, _24051_);
  not (_05480_, _05478_);
  and (_05481_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  or (_26817_, _05481_, _05479_);
  and (_05482_, _05456_, _24219_);
  and (_05484_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_00007_, _05484_, _05482_);
  and (_05485_, _24899_, _24408_);
  and (_05486_, _05485_, _24051_);
  not (_05487_, _05485_);
  and (_05488_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_00019_, _05488_, _05486_);
  and (_05489_, _05478_, _24134_);
  and (_05490_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  or (_00022_, _05490_, _05489_);
  and (_05491_, _24408_, _24223_);
  and (_05492_, _05491_, _23996_);
  not (_05493_, _05491_);
  and (_05494_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  or (_00032_, _05494_, _05492_);
  and (_05495_, _05460_, _23548_);
  and (_05496_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_00044_, _05496_, _05495_);
  and (_05497_, _02045_, _23548_);
  and (_05498_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_00074_, _05498_, _05497_);
  and (_05499_, _05460_, _23887_);
  and (_05500_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_00079_, _05500_, _05499_);
  and (_05501_, _05478_, _23996_);
  and (_05502_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  or (_00082_, _05502_, _05501_);
  and (_05504_, _05491_, _24089_);
  and (_05505_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  or (_00087_, _05505_, _05504_);
  and (_05506_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  and (_05507_, _04937_, _23996_);
  or (_00103_, _05507_, _05506_);
  and (_05508_, _05465_, _24219_);
  and (_05509_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  or (_00172_, _05509_, _05508_);
  or (_05510_, _03083_, _00143_);
  or (_05511_, _05510_, _26816_);
  not (_05512_, _03083_);
  or (_05513_, _05512_, _00191_);
  nand (_05514_, _05513_, _05511_);
  and (_05515_, _05514_, _22888_);
  nor (_05516_, _05514_, _22888_);
  nor (_05517_, _05516_, _05515_);
  and (_05518_, _05510_, _03700_);
  nor (_05519_, _05518_, _24096_);
  and (_05520_, _05510_, _00051_);
  nor (_05521_, _05520_, _24001_);
  nor (_05522_, _05521_, _05519_);
  nor (_05523_, _22968_, _22871_);
  not (_05524_, _05523_);
  not (_05525_, _05510_);
  nor (_05526_, _05525_, _00090_);
  nor (_05527_, _05526_, _05524_);
  and (_05528_, _05526_, _05524_);
  nor (_05529_, _05528_, _05527_);
  and (_05530_, _05529_, _05522_);
  and (_05531_, _05530_, _05517_);
  not (_05532_, _22953_);
  nor (_05533_, _05510_, _00051_);
  nor (_05534_, _05512_, _00228_);
  nor (_05535_, _05534_, _05533_);
  nor (_05536_, _05535_, _05532_);
  and (_05537_, _05535_, _05532_);
  nor (_05538_, _05537_, _05536_);
  not (_05539_, _05538_);
  and (_05540_, _05510_, _26816_);
  and (_05541_, _05525_, _00090_);
  nor (_05542_, _05541_, _05540_);
  and (_05543_, _05542_, _22972_);
  nor (_05544_, _05542_, _22972_);
  or (_05545_, _05544_, _05543_);
  nor (_05546_, _05545_, _05539_);
  or (_05547_, _05510_, _00027_);
  or (_05548_, _05512_, _00171_);
  nand (_05549_, _05548_, _05547_);
  and (_05550_, _05549_, _22921_);
  nor (_05551_, _05549_, _22921_);
  nor (_05552_, _05551_, _05550_);
  and (_05553_, _05520_, _24001_);
  not (_05554_, _05553_);
  and (_05555_, _05518_, _24096_);
  not (_05556_, _05555_);
  nor (_05558_, _00146_, _22849_);
  and (_05559_, _05558_, _05556_);
  and (_05560_, _05559_, _05554_);
  and (_05561_, _05560_, _05552_);
  and (_05562_, _05561_, _05546_);
  and (_05563_, _05562_, _05531_);
  and (_26890_, _05563_, _22731_);
  and (_26891_[7], _23995_, _22731_);
  nor (_26893_[2], _00228_, rst);
  and (_05565_, _04865_, _24051_);
  and (_05566_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or (_00184_, _05566_, _05565_);
  and (_05567_, _02039_, _22974_);
  not (_05568_, _05567_);
  and (_05569_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  and (_05570_, _05567_, _23548_);
  or (_00203_, _05570_, _05569_);
  and (_05571_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  and (_05572_, _05567_, _23583_);
  or (_00209_, _05572_, _05571_);
  and (_05573_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  and (_05574_, _05567_, _24051_);
  or (_00212_, _05574_, _05573_);
  and (_05576_, _03281_, _23996_);
  and (_05577_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or (_00215_, _05577_, _05576_);
  and (_05578_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  and (_05579_, _05567_, _24134_);
  or (_00262_, _05579_, _05578_);
  and (_05580_, _02039_, _24223_);
  not (_05582_, _05580_);
  and (_05583_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_05584_, _05580_, _23548_);
  or (_00270_, _05584_, _05583_);
  and (_05585_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_05587_, _05580_, _23583_);
  or (_00276_, _05587_, _05585_);
  and (_05589_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_05591_, _05580_, _24051_);
  or (_00280_, _05591_, _05589_);
  and (_05592_, _04920_, _23996_);
  and (_05593_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_00289_, _05593_, _05592_);
  and (_05594_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_05595_, _05580_, _24134_);
  or (_00291_, _05595_, _05594_);
  and (_05596_, _02039_, _24056_);
  not (_05597_, _05596_);
  and (_05598_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  and (_05599_, _05596_, _24219_);
  or (_00299_, _05599_, _05598_);
  and (_05600_, _03275_, _23887_);
  and (_05601_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or (_00302_, _05601_, _05600_);
  and (_05603_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  and (_05604_, _05596_, _23887_);
  or (_00305_, _05604_, _05603_);
  and (_05605_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  and (_05606_, _05596_, _24089_);
  or (_00310_, _05606_, _05605_);
  and (_26891_[0], _24218_, _22731_);
  and (_26891_[1], _23547_, _22731_);
  and (_26891_[2], _23886_, _22731_);
  and (_26891_[3], _23582_, _22731_);
  and (_26891_[4], _24088_, _22731_);
  and (_26891_[5], _24050_, _22731_);
  and (_26891_[6], _24133_, _22731_);
  nor (_26893_[0], _00191_, rst);
  nor (_26893_[1], _00171_, rst);
  and (_05609_, _05491_, _23548_);
  and (_05610_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  or (_00515_, _05610_, _05609_);
  nor (_05611_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_05612_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01836_);
  nor (_05613_, _05612_, _05611_);
  not (_05614_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_05615_, _00613_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_05616_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01836_);
  nor (_05617_, _05616_, _05615_);
  nor (_05618_, _05617_, _05614_);
  and (_05619_, _05617_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_05620_, _05619_, _05618_);
  not (_05621_, _05620_);
  nor (_05622_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_05623_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01836_);
  nor (_05624_, _05623_, _05622_);
  not (_05625_, _05624_);
  nor (_05626_, _00517_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_05627_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01836_);
  nor (_05628_, _05627_, _05626_);
  and (_05629_, _05628_, _05625_);
  nand (_05630_, _05629_, _05621_);
  and (_05631_, _05630_, _05613_);
  nor (_05632_, _05628_, _05625_);
  not (_05633_, _05632_);
  not (_05634_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_05635_, _05617_, _05634_);
  and (_05636_, _05617_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05637_, _05636_, _05635_);
  nor (_05638_, _05637_, _05633_);
  and (_05639_, _05628_, _05624_);
  not (_05640_, _05639_);
  not (_05641_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_05642_, _05617_, _05641_);
  and (_05643_, _05617_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_05645_, _05643_, _05642_);
  nor (_05646_, _05645_, _05640_);
  nor (_05647_, _05646_, _05638_);
  nor (_05649_, _05628_, _05624_);
  not (_05651_, _05649_);
  and (_05652_, _05617_, \oc8051_symbolic_cxrom1.regvalid [9]);
  not (_05653_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_05654_, _05617_, _05653_);
  nor (_05655_, _05654_, _05652_);
  or (_05656_, _05655_, _05651_);
  and (_05657_, _05656_, _05647_);
  and (_05658_, _05657_, _05631_);
  not (_05659_, _05628_);
  not (_05660_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_05661_, _05617_, _05660_);
  and (_05662_, _05617_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_05663_, _05662_, _05661_);
  nor (_05664_, _05663_, _05659_);
  not (_05665_, _05664_);
  nor (_05667_, _05628_, _05617_);
  and (_05668_, _05667_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05669_, _05659_, _05617_);
  and (_05670_, _05669_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_05671_, _05670_, _05668_);
  and (_05672_, _05671_, _05665_);
  nor (_05673_, _05672_, _05624_);
  and (_05674_, _05667_, _05624_);
  and (_05675_, _05674_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not (_05677_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_05678_, _05617_, _05677_);
  nor (_05679_, _05617_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_05680_, _05679_, _05678_);
  nor (_05681_, _05680_, _05640_);
  and (_05682_, _05617_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_05683_, _05682_, _05632_);
  or (_05684_, _05683_, _05613_);
  or (_05685_, _05684_, _05681_);
  or (_05686_, _05685_, _05675_);
  nor (_05687_, _05686_, _05673_);
  nor (_05688_, _05687_, _05658_);
  not (_05689_, _05688_);
  and (_05690_, _05689_, word_in[7]);
  not (_05691_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_05692_, _05613_, _05691_);
  or (_05693_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_05694_, _05693_, _05692_);
  and (_05696_, _05694_, _05639_);
  not (_05697_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_05698_, _05613_, _05697_);
  or (_05699_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_05700_, _05699_, _05698_);
  and (_05701_, _05700_, _05632_);
  or (_05702_, _05701_, _05696_);
  not (_05704_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_05705_, _05613_, _05704_);
  or (_05706_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_05707_, _05706_, _05705_);
  and (_05708_, _05707_, _05629_);
  not (_05709_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_05710_, _05613_, _05709_);
  or (_05711_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_05712_, _05711_, _05710_);
  and (_05713_, _05712_, _05649_);
  or (_05715_, _05713_, _05708_);
  or (_05716_, _05715_, _05702_);
  and (_05717_, _05716_, _05617_);
  not (_05719_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_05720_, _05613_, _05719_);
  or (_05721_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_05722_, _05721_, _05720_);
  and (_05723_, _05722_, _05674_);
  not (_05724_, _05617_);
  and (_05725_, _05639_, _05724_);
  not (_05726_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_05727_, _05613_, _05726_);
  or (_05728_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_05730_, _05728_, _05727_);
  and (_05731_, _05730_, _05725_);
  not (_05732_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_05733_, _05613_, _05732_);
  or (_05734_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_05735_, _05734_, _05733_);
  and (_05736_, _05735_, _05629_);
  not (_05737_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_05738_, _05613_, _05737_);
  or (_05739_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_05741_, _05739_, _05738_);
  and (_05742_, _05741_, _05649_);
  or (_05743_, _05742_, _05736_);
  and (_05744_, _05743_, _05724_);
  or (_05745_, _05744_, _05731_);
  or (_05746_, _05745_, _05723_);
  or (_05747_, _05746_, _05717_);
  and (_05748_, _05747_, _05688_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _05748_, _05690_);
  and (_05749_, _03275_, _24134_);
  and (_05750_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_00527_, _05750_, _05749_);
  and (_05751_, _05625_, _05613_);
  not (_05752_, _05751_);
  and (_05753_, _05624_, _05613_);
  and (_05754_, _05753_, _05628_);
  nor (_05755_, _05753_, _05628_);
  nor (_05756_, _05755_, _05754_);
  not (_05757_, _05756_);
  nor (_05758_, _05757_, _05680_);
  nor (_05759_, _05754_, _05724_);
  nor (_05760_, _05659_, _05617_);
  and (_05761_, _05760_, _05753_);
  nor (_05762_, _05761_, _05759_);
  nor (_05763_, _05762_, _05756_);
  and (_05765_, _05763_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_05766_, _05755_, _05617_);
  nor (_05767_, _05766_, _05759_);
  and (_05768_, _05767_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_05769_, _05768_, _05765_);
  nor (_05770_, _05769_, _05758_);
  nor (_05771_, _05770_, _05752_);
  not (_05772_, _05753_);
  nor (_05773_, _05757_, _05663_);
  and (_05774_, _05767_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_05775_, _05774_, _05773_);
  or (_05776_, _05775_, _05772_);
  nand (_05777_, _05761_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05779_, _05777_, _05776_);
  not (_05780_, _05779_);
  nor (_05782_, _05780_, _05771_);
  nor (_05784_, _05624_, _05613_);
  or (_05785_, _05753_, _05784_);
  not (_05787_, _05785_);
  nor (_05789_, _05757_, _05620_);
  and (_05790_, _05763_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05792_, _05767_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05793_, _05792_, _05790_);
  nor (_05795_, _05793_, _05789_);
  or (_05796_, _05795_, _05787_);
  and (_05797_, _05756_, _05724_);
  and (_05798_, _05797_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_05799_, _05763_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_05800_, _05756_, _05617_);
  and (_05801_, _05800_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_05802_, _05767_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_05803_, _05802_, _05801_);
  or (_05804_, _05803_, _05799_);
  nor (_05806_, _05804_, _05798_);
  or (_05807_, _05806_, _05785_);
  and (_05808_, _05807_, _05796_);
  or (_05809_, _05808_, _05613_);
  and (_05810_, _05809_, _05782_);
  not (_05811_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_05813_, _05613_, _05811_);
  or (_05814_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_05815_, _05814_, _05813_);
  and (_05817_, _05815_, _05787_);
  not (_05818_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_05819_, _05613_, _05818_);
  or (_05821_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_05822_, _05821_, _05819_);
  and (_05823_, _05822_, _05785_);
  or (_05824_, _05823_, _05817_);
  and (_05826_, _05824_, _05800_);
  not (_05827_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_05828_, _05613_, _05827_);
  or (_05829_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_05830_, _05829_, _05828_);
  and (_05831_, _05830_, _05787_);
  not (_05832_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_05834_, _05613_, _05832_);
  or (_05835_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_05836_, _05835_, _05834_);
  and (_05837_, _05836_, _05785_);
  or (_05838_, _05837_, _05831_);
  and (_05839_, _05838_, _05763_);
  or (_05841_, _05839_, _05826_);
  not (_05842_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_05844_, _05613_, _05842_);
  or (_05845_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_05846_, _05845_, _05844_);
  and (_05847_, _05846_, _05785_);
  not (_05848_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_05849_, _05613_, _05848_);
  or (_05850_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_05851_, _05850_, _05849_);
  and (_05852_, _05851_, _05787_);
  or (_05853_, _05852_, _05847_);
  and (_05854_, _05853_, _05767_);
  not (_05855_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_05856_, _05613_, _05855_);
  or (_05857_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_05858_, _05857_, _05856_);
  and (_05860_, _05858_, _05785_);
  not (_05862_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_05863_, _05613_, _05862_);
  or (_05864_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_05865_, _05864_, _05863_);
  and (_05867_, _05865_, _05787_);
  or (_05868_, _05867_, _05860_);
  and (_05869_, _05868_, _05797_);
  or (_05870_, _05869_, _05854_);
  nor (_05871_, _05870_, _05841_);
  nor (_05872_, _05871_, _05810_);
  and (_05873_, _05810_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _05873_, _05872_);
  and (_05874_, _05639_, _05617_);
  and (_05875_, _05649_, _05724_);
  or (_05876_, _05875_, _05874_);
  and (_05877_, _05876_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_05878_, _05877_);
  nor (_05879_, _05639_, _05649_);
  not (_05880_, _05879_);
  nor (_05881_, _05880_, _05620_);
  or (_05883_, _05639_, _05617_);
  or (_05884_, _05649_, _05724_);
  and (_05885_, _05884_, _05883_);
  and (_05886_, _05885_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_05887_, _05886_, _05881_);
  and (_05888_, _05887_, _05878_);
  nor (_05889_, _05888_, _05772_);
  nor (_05890_, _05880_, _05645_);
  and (_05891_, _05876_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_05893_, _05885_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05894_, _05893_, _05891_);
  nor (_05895_, _05894_, _05890_);
  nor (_05896_, _05895_, _05752_);
  nor (_05897_, _05896_, _05889_);
  not (_05898_, _05784_);
  nor (_05899_, _05880_, _05680_);
  and (_05900_, _05876_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_05901_, _05885_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05902_, _05901_, _05900_);
  nor (_05903_, _05902_, _05899_);
  nor (_05904_, _05903_, _05898_);
  not (_05905_, _05613_);
  and (_05906_, _05624_, _05905_);
  not (_05907_, _05906_);
  nor (_05908_, _05880_, _05663_);
  and (_05910_, _05876_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05911_, _05885_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05912_, _05911_, _05910_);
  nor (_05914_, _05912_, _05908_);
  nor (_05915_, _05914_, _05907_);
  nor (_05916_, _05915_, _05904_);
  and (_05918_, _05916_, _05897_);
  and (_05919_, _05918_, word_in[23]);
  and (_05920_, _05640_, _05617_);
  or (_05921_, _05920_, _05725_);
  and (_05922_, _05730_, _05629_);
  and (_05923_, _05722_, _05649_);
  or (_05924_, _05923_, _05922_);
  and (_05925_, _05735_, _05632_);
  and (_05926_, _05741_, _05639_);
  or (_05927_, _05926_, _05925_);
  or (_05929_, _05927_, _05924_);
  or (_05930_, _05929_, _05921_);
  and (_05931_, _05707_, _05632_);
  and (_05933_, _05700_, _05649_);
  or (_05934_, _05933_, _05931_);
  and (_05936_, _05694_, _05629_);
  and (_05937_, _05712_, _05639_);
  or (_05938_, _05937_, _05936_);
  nor (_05939_, _05938_, _05934_);
  nand (_05941_, _05939_, _05921_);
  nand (_05942_, _05941_, _05930_);
  nor (_05943_, _05942_, _05918_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _05943_, _05919_);
  and (_05944_, _03269_, _24089_);
  and (_05946_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  or (_00541_, _05946_, _05944_);
  and (_05947_, _05898_, _05628_);
  nor (_05948_, _05898_, _05628_);
  nor (_05949_, _05948_, _05947_);
  not (_05950_, _05949_);
  or (_05952_, _05950_, _05663_);
  and (_05953_, _05947_, _05617_);
  nor (_05955_, _05947_, _05617_);
  nor (_05956_, _05955_, _05953_);
  and (_05957_, _05956_, _05950_);
  nand (_05958_, _05957_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05959_, _05958_, _05952_);
  or (_05961_, _05959_, _05752_);
  and (_05962_, _05628_, _05617_);
  and (_05963_, _05751_, _05962_);
  and (_05964_, _05963_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05965_, _05754_, _05617_);
  and (_05966_, _05965_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_05967_, _05680_, _05950_);
  and (_05968_, _05957_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05969_, _05968_, _05967_);
  and (_05970_, _05969_, _05753_);
  or (_05971_, _05970_, _05966_);
  nor (_05972_, _05971_, _05964_);
  and (_05973_, _05972_, _05961_);
  or (_05975_, _05950_, _05620_);
  nand (_05976_, _05957_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05977_, _05976_, _05975_);
  or (_05979_, _05977_, _05907_);
  and (_05980_, _05948_, _05635_);
  and (_05982_, _05874_, _05905_);
  and (_05983_, _05982_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_05984_, _05950_, _05645_);
  and (_05985_, _05957_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05986_, _05985_, _05984_);
  and (_05987_, _05986_, _05784_);
  or (_05988_, _05987_, _05983_);
  nor (_05989_, _05988_, _05980_);
  and (_05990_, _05989_, _05979_);
  and (_05991_, _05990_, _05973_);
  and (_05992_, _05836_, _05787_);
  and (_05993_, _05830_, _05785_);
  or (_05994_, _05993_, _05992_);
  and (_05995_, _05994_, _05957_);
  nor (_05996_, _05956_, _05949_);
  and (_05997_, _05846_, _05787_);
  and (_05999_, _05851_, _05785_);
  or (_06000_, _05999_, _05997_);
  and (_06001_, _06000_, _05996_);
  not (_06002_, _05948_);
  and (_06003_, _05955_, _06002_);
  and (_06004_, _05858_, _05787_);
  and (_06005_, _05865_, _05785_);
  or (_06006_, _06005_, _06004_);
  and (_06007_, _06006_, _06003_);
  and (_06008_, _05949_, _05617_);
  and (_06009_, _05822_, _05787_);
  and (_06010_, _05815_, _05785_);
  or (_06011_, _06010_, _06009_);
  and (_06012_, _06011_, _06008_);
  or (_06013_, _06012_, _06007_);
  or (_06014_, _06013_, _06001_);
  nor (_06015_, _06014_, _05995_);
  nor (_06016_, _06015_, _05991_);
  and (_06017_, _05991_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _06017_, _06016_);
  or (_06018_, _05962_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_26822_[15], _06018_, _22731_);
  and (_06019_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  and (_06020_, _05596_, _24051_);
  or (_00596_, _06020_, _06019_);
  and (_06022_, _05918_, _22731_);
  and (_06023_, _06022_, _05879_);
  and (_06024_, _06023_, _05921_);
  and (_06026_, _06024_, _05751_);
  not (_06027_, _06026_);
  and (_06028_, _05810_, _22731_);
  and (_06029_, _06028_, _05906_);
  and (_06030_, _06029_, _05800_);
  and (_06031_, _05658_, _22731_);
  and (_06032_, _06031_, _05624_);
  nor (_06033_, _05688_, rst);
  and (_06034_, _06033_, _05962_);
  and (_06035_, _06034_, _06032_);
  and (_06036_, _06035_, word_in[7]);
  nor (_06037_, _06035_, _05691_);
  nor (_06038_, _06037_, _06036_);
  nor (_06039_, _06038_, _06030_);
  and (_06040_, _06030_, word_in[15]);
  or (_06041_, _06040_, _06039_);
  and (_06042_, _06041_, _06027_);
  and (_06043_, _05991_, _22731_);
  and (_06044_, _06043_, _05784_);
  and (_06046_, _06044_, _05962_);
  and (_06047_, _06022_, word_in[23]);
  and (_06048_, _06047_, _06026_);
  or (_06049_, _06048_, _06046_);
  or (_06050_, _06049_, _06042_);
  not (_06051_, _06046_);
  and (_06052_, _06043_, word_in[31]);
  or (_06053_, _06052_, _06051_);
  and (_26829_[7], _06053_, _06050_);
  or (_06055_, _05996_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_26839_, _06055_, _22731_);
  and (_06057_, _04920_, _24134_);
  and (_06058_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_00657_, _06058_, _06057_);
  or (_06060_, _05965_, _05875_);
  or (_06061_, _05982_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_06062_, _06061_, _06060_);
  and (_26822_[1], _06062_, _22731_);
  and (_06063_, _03001_, _23887_);
  and (_06064_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_00674_, _06064_, _06063_);
  or (_06066_, _05617_, _05613_);
  nor (_06067_, _06066_, _05633_);
  or (_06069_, _06067_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_06070_, _06060_, _06069_);
  and (_26822_[2], _06070_, _22731_);
  or (_06072_, _05667_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_26822_[3], _06072_, _22731_);
  and (_06073_, _05753_, _05667_);
  and (_06074_, _05751_, _06003_);
  and (_06075_, _05948_, _05724_);
  and (_06077_, _06075_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_06078_, _06077_, _06074_);
  not (_06079_, _05667_);
  and (_06080_, _05760_, _05784_);
  or (_06081_, _06080_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_06082_, _06081_, _06079_);
  or (_06083_, _06082_, _06078_);
  or (_06084_, _06083_, _06073_);
  or (_06085_, _06084_, _06067_);
  and (_26822_[4], _06085_, _22731_);
  or (_06087_, _06080_, _06073_);
  or (_06089_, _06087_, _05883_);
  and (_06090_, _06089_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_06091_, _05760_, _05751_);
  and (_06092_, _06067_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_06093_, _06092_, _06091_);
  nor (_06094_, _06093_, _06090_);
  nor (_06096_, _06094_, _05955_);
  and (_06097_, _05649_, _05618_);
  or (_06098_, _06097_, _06067_);
  or (_06099_, _06098_, _06080_);
  or (_06100_, _06099_, _06073_);
  or (_06101_, _06100_, _06096_);
  and (_26822_[5], _06101_, _22731_);
  and (_06102_, _05947_, _05724_);
  or (_06103_, _05759_, _06102_);
  or (_06104_, _05759_, _05725_);
  nor (_06105_, _06066_, _05640_);
  not (_06106_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_06108_, _05667_, _06106_);
  and (_06109_, _06108_, _06066_);
  or (_06110_, _06109_, _06105_);
  and (_06111_, _06110_, _06104_);
  and (_06112_, _06087_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_06113_, _06112_, _06091_);
  or (_06114_, _06113_, _06111_);
  and (_06115_, _06114_, _06103_);
  or (_06116_, _06112_, _06110_);
  and (_06117_, _06116_, _05965_);
  and (_06118_, _06067_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_06119_, _05875_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_06121_, _06119_, _06073_);
  or (_06122_, _06121_, _06118_);
  or (_06124_, _06122_, _06080_);
  or (_06125_, _06124_, _06117_);
  or (_06126_, _06125_, _06115_);
  and (_26822_[6], _06126_, _22731_);
  and (_06127_, _24320_, _24219_);
  and (_06128_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_00972_, _06128_, _06127_);
  and (_06129_, _24496_, _24223_);
  and (_06130_, _06129_, _23996_);
  not (_06131_, _06129_);
  and (_06132_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  or (_00985_, _06132_, _06130_);
  and (_06133_, _25658_, _24219_);
  and (_06134_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or (_00994_, _06134_, _06133_);
  or (_06135_, _05754_, _05617_);
  or (_06136_, _06105_, _05617_);
  and (_06137_, _06136_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_06138_, _05642_, _05640_);
  or (_06139_, _06138_, _05761_);
  or (_06140_, _06139_, _06137_);
  and (_06141_, _06140_, _06135_);
  and (_06142_, _05667_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_06143_, _06142_, _06080_);
  or (_06144_, _06143_, _06091_);
  or (_06145_, _06144_, _06105_);
  or (_06146_, _06145_, _06141_);
  and (_26822_[7], _06146_, _22731_);
  or (_06148_, _05957_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_26822_[8], _06148_, _22731_);
  and (_06150_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  and (_06152_, _02513_, _24219_);
  or (_01070_, _06152_, _06150_);
  nand (_06153_, _02294_, _24082_);
  or (_06154_, _02616_, _02281_);
  and (_06155_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_06156_, _02283_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_06157_, _06156_, _02285_);
  not (_06158_, _02281_);
  nor (_06159_, _02258_, _02249_);
  nor (_06160_, _06159_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_06162_, _02259_, _02248_);
  nor (_06163_, _06162_, _06160_);
  and (_06164_, _06163_, _06158_);
  nor (_06165_, _06164_, _06157_);
  nor (_06166_, _06165_, _02616_);
  or (_06167_, _06166_, _06155_);
  or (_06168_, _06167_, _02294_);
  and (_06170_, _06168_, _22731_);
  and (_01093_, _06170_, _06153_);
  and (_06171_, _05759_, _06002_);
  and (_06172_, _05725_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_06173_, _05751_, _06008_);
  or (_06174_, _06173_, _05652_);
  or (_06175_, _06174_, _06172_);
  and (_06176_, _06175_, _06171_);
  and (_06177_, _05948_, _05617_);
  or (_06178_, _06172_, _06177_);
  or (_06180_, _06178_, _06176_);
  and (_06181_, _06180_, _05759_);
  and (_06182_, _06175_, _05965_);
  or (_06183_, _06091_, _06003_);
  and (_06184_, _06183_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_06185_, _06075_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_06186_, _06185_, _05725_);
  or (_06187_, _06186_, _06184_);
  or (_06188_, _06187_, _06182_);
  or (_06189_, _06188_, _06181_);
  and (_26822_[9], _06189_, _22731_);
  and (_06190_, _05906_, _06008_);
  not (_06191_, _05755_);
  and (_06192_, _06191_, _05682_);
  or (_06193_, _06192_, _06190_);
  and (_06194_, _05879_, _05724_);
  and (_06195_, _06194_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_06196_, _06105_, _05875_);
  and (_06197_, _06196_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_06198_, _06197_, _05761_);
  or (_06199_, _06198_, _06195_);
  or (_06200_, _06199_, _06177_);
  or (_06201_, _06200_, _06173_);
  or (_06202_, _06201_, _06193_);
  and (_26822_[10], _06202_, _22731_);
  and (_06203_, _02512_, _24140_);
  not (_06204_, _06203_);
  and (_06205_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_06206_, _06203_, _23996_);
  or (_01196_, _06206_, _06205_);
  and (_06208_, _24474_, _24301_);
  and (_06209_, _06208_, _23887_);
  not (_06210_, _06208_);
  and (_06211_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_01224_, _06211_, _06209_);
  and (_06212_, _25658_, _23583_);
  and (_06213_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  or (_01235_, _06213_, _06212_);
  and (_06215_, _25658_, _23887_);
  and (_06216_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  or (_01254_, _06216_, _06215_);
  and (_06217_, _05787_, _05667_);
  or (_06218_, _06217_, _05766_);
  or (_06219_, _06218_, _05962_);
  and (_06220_, _06219_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_06221_, _05753_, _06008_);
  and (_06222_, _06075_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_06223_, _06222_, _06177_);
  or (_06224_, _06223_, _06173_);
  or (_06226_, _06224_, _06190_);
  or (_06227_, _06226_, _06221_);
  or (_06228_, _06227_, _06220_);
  and (_26822_[11], _06228_, _22731_);
  and (_06230_, _25637_, _24051_);
  and (_06231_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_01301_, _06231_, _06230_);
  and (_06233_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  and (_06234_, _02513_, _23548_);
  or (_01307_, _06234_, _06233_);
  and (_06236_, _02527_, _25481_);
  nand (_06237_, _06236_, _23504_);
  or (_06238_, _06236_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_06240_, _06238_, _02534_);
  and (_06241_, _06240_, _06237_);
  nor (_06242_, _02534_, _23989_);
  or (_06244_, _06242_, _06241_);
  and (_01332_, _06244_, _22731_);
  or (_06245_, _02925_, _02865_);
  and (_06246_, _06245_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_06247_, _06246_, _02898_);
  and (_01334_, _06247_, _22731_);
  nor (_01336_, _04686_, rst);
  and (_06249_, _24008_, _23583_);
  and (_06250_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_27083_, _06250_, _06249_);
  or (_06251_, _05957_, _05724_);
  and (_06252_, _06251_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_06253_, _05953_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_06254_, _06253_, _06008_);
  or (_06255_, _06254_, _06252_);
  and (_26822_[12], _06255_, _22731_);
  and (_06256_, _02078_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_06257_, _02080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_01355_, _06257_, _06256_);
  or (_06258_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_06259_, _06258_, _22731_);
  and (_06260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or (_06261_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_06262_, _06261_, rxd_i);
  or (_06263_, _06262_, _06260_);
  and (_06264_, _06263_, _02785_);
  and (_06265_, _02812_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_06267_, _06265_, _06264_);
  and (_06269_, _02799_, rxd_i);
  or (_06270_, _06269_, _02810_);
  or (_06271_, _06270_, _06267_);
  and (_01368_, _06271_, _06259_);
  and (_06272_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  and (_06273_, _02513_, _23887_);
  or (_01379_, _06273_, _06272_);
  and (_06274_, _04865_, _24219_);
  and (_06276_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_01388_, _06276_, _06274_);
  and (_06278_, _06129_, _23887_);
  and (_06279_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or (_01392_, _06279_, _06278_);
  and (_06281_, _02970_, _23548_);
  and (_06283_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  or (_01404_, _06283_, _06281_);
  and (_06284_, _06129_, _23548_);
  and (_06286_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  or (_01407_, _06286_, _06284_);
  and (_06287_, _02877_, _02780_);
  and (_06289_, _02867_, _06287_);
  nand (_06290_, _06289_, _02900_);
  or (_06291_, _06289_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_06292_, _06291_, _22731_);
  and (_01409_, _06292_, _06290_);
  and (_06293_, _05632_, _05617_);
  or (_06294_, _05963_, _06293_);
  and (_06295_, _05962_, _05784_);
  and (_06296_, _05874_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_06298_, _05884_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or (_06299_, _06298_, _06296_);
  or (_06300_, _06299_, _06295_);
  or (_06301_, _06300_, _06294_);
  and (_26822_[13], _06301_, _22731_);
  nor (_06302_, _02792_, _02786_);
  and (_06303_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _02900_);
  and (_06305_, _06303_, _02792_);
  or (_06306_, _06305_, _06302_);
  and (_06307_, _06306_, _02569_);
  not (_06308_, _02798_);
  nand (_06310_, _02824_, _06308_);
  or (_06311_, _06310_, _06307_);
  and (_01421_, _06311_, _02080_);
  or (_06312_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_06313_, _06312_, _22731_);
  nand (_06315_, _02071_, _23989_);
  and (_01423_, _06315_, _06313_);
  not (_06316_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_06317_, _02652_, _06316_);
  or (_06318_, _06317_, _04703_);
  and (_06319_, _06318_, _02649_);
  nand (_06320_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_06321_, _06320_, _02648_);
  nor (_06322_, _06321_, _06319_);
  nor (_06323_, _06322_, _02647_);
  or (_06324_, _06323_, _02757_);
  nand (_06325_, _06324_, _22731_);
  nor (_01426_, _06325_, _02658_);
  or (_06326_, _05800_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_26822_[14], _06326_, _22731_);
  and (_06328_, _06129_, _24051_);
  and (_06329_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  or (_01495_, _06329_, _06328_);
  and (_06330_, _24008_, _23887_);
  and (_06331_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_01500_, _06331_, _06330_);
  and (_06332_, _02970_, _24219_);
  and (_06334_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  or (_01504_, _06334_, _06332_);
  and (_06335_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  and (_06337_, _05596_, _23996_);
  or (_01600_, _06337_, _06335_);
  and (_06339_, _02039_, _24474_);
  not (_06341_, _06339_);
  and (_06342_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_06343_, _06339_, _24219_);
  or (_01604_, _06343_, _06342_);
  and (_06344_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_06345_, _06339_, _23887_);
  or (_01606_, _06345_, _06344_);
  and (_06347_, _03245_, _24089_);
  and (_06348_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  or (_27170_, _06348_, _06347_);
  and (_06351_, _02767_, _23583_);
  and (_06352_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or (_01662_, _06352_, _06351_);
  and (_06353_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_06354_, _06339_, _23583_);
  or (_27015_, _06354_, _06353_);
  and (_06356_, _25413_, _24159_);
  and (_06357_, _06356_, _24089_);
  not (_06358_, _06356_);
  and (_06359_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_01688_, _06359_, _06357_);
  and (_06360_, _06356_, _23887_);
  and (_06361_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_01698_, _06361_, _06360_);
  and (_06362_, _06356_, _23996_);
  and (_06363_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_01729_, _06363_, _06362_);
  and (_06364_, _06043_, word_in[24]);
  and (_06365_, _06364_, _05963_);
  and (_06366_, _06022_, _05982_);
  and (_06367_, _06028_, _05965_);
  not (_06368_, _06367_);
  and (_06369_, _06033_, _05624_);
  nor (_06370_, _06369_, _06031_);
  and (_06371_, _06033_, _05667_);
  and (_06372_, _06371_, _06370_);
  and (_06374_, _06372_, word_in[0]);
  not (_06375_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_06376_, _06372_, _06375_);
  or (_06377_, _06376_, _06374_);
  and (_06378_, _06377_, _06368_);
  and (_06379_, _06367_, word_in[8]);
  or (_06381_, _06379_, _06378_);
  or (_06383_, _06381_, _06366_);
  and (_06384_, _06043_, _05963_);
  not (_06385_, _06384_);
  not (_06386_, _06366_);
  or (_06387_, _06386_, word_in[16]);
  and (_06388_, _06387_, _06385_);
  and (_06389_, _06388_, _06383_);
  or (_26823_[0], _06389_, _06365_);
  and (_06391_, _06022_, word_in[17]);
  and (_06392_, _06391_, _05982_);
  not (_06393_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_06394_, _06372_, _06393_);
  and (_06395_, _06372_, word_in[1]);
  or (_06397_, _06395_, _06394_);
  and (_06398_, _06397_, _06368_);
  and (_06399_, _06367_, word_in[9]);
  or (_06400_, _06399_, _06398_);
  and (_06402_, _06400_, _06386_);
  or (_06404_, _06402_, _06392_);
  and (_06405_, _06404_, _06385_);
  and (_06406_, _06384_, word_in[25]);
  or (_26823_[1], _06406_, _06405_);
  and (_06407_, _06043_, word_in[26]);
  and (_06409_, _06407_, _05963_);
  not (_06410_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_06411_, _06372_, _06410_);
  and (_06412_, _06033_, word_in[2]);
  and (_06413_, _06412_, _06372_);
  or (_06415_, _06413_, _06411_);
  or (_06417_, _06415_, _06367_);
  or (_06418_, _06368_, word_in[10]);
  and (_06419_, _06418_, _06417_);
  or (_06421_, _06419_, _06366_);
  or (_06422_, _06386_, word_in[18]);
  and (_06423_, _06422_, _06385_);
  and (_06424_, _06423_, _06421_);
  or (_26823_[2], _06424_, _06409_);
  not (_06425_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_06426_, _06372_, _06425_);
  and (_06427_, _06033_, word_in[3]);
  and (_06429_, _06427_, _06372_);
  or (_06430_, _06429_, _06426_);
  or (_06431_, _06430_, _06367_);
  or (_06432_, _06368_, word_in[11]);
  and (_06433_, _06432_, _06431_);
  or (_06435_, _06433_, _06366_);
  or (_06437_, _06386_, word_in[19]);
  and (_06438_, _06437_, _06385_);
  and (_06440_, _06438_, _06435_);
  and (_06441_, _06043_, word_in[27]);
  and (_06443_, _06441_, _05963_);
  or (_26823_[3], _06443_, _06440_);
  and (_06446_, _06043_, word_in[28]);
  and (_06447_, _06446_, _05963_);
  not (_06448_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_06449_, _06372_, _06448_);
  and (_06450_, _06033_, word_in[4]);
  and (_06451_, _06450_, _06372_);
  or (_06452_, _06451_, _06449_);
  or (_06453_, _06452_, _06367_);
  or (_06454_, _06368_, word_in[12]);
  and (_06455_, _06454_, _06453_);
  or (_06456_, _06455_, _06366_);
  or (_06458_, _06386_, word_in[20]);
  and (_06460_, _06458_, _06385_);
  and (_06461_, _06460_, _06456_);
  or (_26823_[4], _06461_, _06447_);
  and (_06463_, _06043_, word_in[29]);
  and (_06464_, _06463_, _05963_);
  not (_06466_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_06468_, _06372_, _06466_);
  and (_06469_, _06033_, word_in[5]);
  and (_06470_, _06469_, _06372_);
  or (_06471_, _06470_, _06468_);
  or (_06472_, _06471_, _06367_);
  or (_06473_, _06368_, word_in[13]);
  and (_06474_, _06473_, _06472_);
  or (_06475_, _06474_, _06366_);
  or (_06476_, _06386_, word_in[21]);
  and (_06478_, _06476_, _06385_);
  and (_06479_, _06478_, _06475_);
  or (_26823_[5], _06479_, _06464_);
  and (_06480_, _06384_, word_in[30]);
  not (_06481_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_06482_, _06372_, _06481_);
  and (_06483_, _06372_, word_in[6]);
  or (_06484_, _06483_, _06482_);
  and (_06486_, _06484_, _06368_);
  and (_06487_, _06367_, word_in[14]);
  or (_06488_, _06487_, _06486_);
  or (_06489_, _06488_, _06366_);
  or (_06490_, _06386_, word_in[22]);
  and (_06491_, _06490_, _06385_);
  and (_06492_, _06491_, _06489_);
  or (_26823_[6], _06492_, _06480_);
  and (_06493_, _24442_, _23583_);
  and (_06494_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  or (_01799_, _06494_, _06493_);
  nor (_06495_, _06372_, _05842_);
  and (_06496_, _06033_, word_in[7]);
  and (_06497_, _06372_, _06496_);
  or (_06498_, _06497_, _06495_);
  or (_06499_, _06498_, _06367_);
  or (_06500_, _06368_, word_in[15]);
  and (_06502_, _06500_, _06499_);
  or (_06503_, _06502_, _06366_);
  or (_06505_, _06386_, word_in[23]);
  and (_06507_, _06505_, _06385_);
  and (_06508_, _06507_, _06503_);
  and (_06509_, _06384_, word_in[31]);
  or (_26823_[7], _06509_, _06508_);
  and (_06512_, _06022_, _05753_);
  and (_06513_, _06512_, _05876_);
  and (_06515_, _06028_, _05784_);
  and (_06516_, _06515_, _05767_);
  not (_06518_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_06520_, _06033_, _06079_);
  and (_06521_, _06031_, _05625_);
  not (_06522_, _06521_);
  nor (_06523_, _06522_, _06520_);
  nor (_06524_, _06523_, _06518_);
  and (_06525_, _06033_, word_in[0]);
  and (_06527_, _06523_, _06525_);
  or (_06528_, _06527_, _06524_);
  or (_06529_, _06528_, _06516_);
  not (_06531_, _06516_);
  or (_06532_, _06531_, word_in[8]);
  and (_06533_, _06532_, _06529_);
  or (_06534_, _06533_, _06513_);
  and (_06535_, _06043_, _05982_);
  not (_06537_, _06535_);
  and (_06538_, _06022_, word_in[16]);
  not (_06539_, _06513_);
  or (_06540_, _06539_, _06538_);
  and (_06542_, _06540_, _06537_);
  and (_06543_, _06542_, _06534_);
  and (_06544_, _06535_, word_in[24]);
  or (_26830_[0], _06544_, _06543_);
  not (_06545_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_06546_, _06523_, _06545_);
  and (_06548_, _06033_, word_in[1]);
  and (_06549_, _06523_, _06548_);
  or (_06550_, _06549_, _06546_);
  or (_06551_, _06550_, _06516_);
  or (_06552_, _06531_, word_in[9]);
  and (_06553_, _06552_, _06551_);
  or (_06554_, _06553_, _06513_);
  or (_06556_, _06539_, _06391_);
  and (_06557_, _06556_, _06537_);
  and (_06559_, _06557_, _06554_);
  and (_06561_, _06535_, word_in[25]);
  or (_26830_[1], _06561_, _06559_);
  not (_06562_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_06563_, _06523_, _06562_);
  and (_06565_, _06523_, _06412_);
  or (_06566_, _06565_, _06563_);
  or (_06567_, _06566_, _06516_);
  or (_06568_, _06531_, word_in[10]);
  and (_06570_, _06568_, _06567_);
  or (_06571_, _06570_, _06513_);
  and (_06572_, _06022_, word_in[18]);
  or (_06573_, _06539_, _06572_);
  and (_06575_, _06573_, _06537_);
  and (_06576_, _06575_, _06571_);
  and (_06577_, _06535_, word_in[26]);
  or (_26830_[2], _06577_, _06576_);
  not (_06578_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_06579_, _06523_, _06578_);
  and (_06580_, _06523_, _06427_);
  or (_06581_, _06580_, _06579_);
  or (_06582_, _06581_, _06516_);
  or (_06583_, _06531_, word_in[11]);
  and (_06584_, _06583_, _06582_);
  or (_06585_, _06584_, _06513_);
  and (_06586_, _06022_, word_in[19]);
  or (_06587_, _06539_, _06586_);
  and (_06588_, _06587_, _06537_);
  and (_06589_, _06588_, _06585_);
  and (_06590_, _06535_, word_in[27]);
  or (_26830_[3], _06590_, _06589_);
  and (_06591_, _06022_, word_in[20]);
  and (_06592_, _06513_, _06591_);
  and (_06593_, _06523_, _06450_);
  not (_06594_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_06595_, _06523_, _06594_);
  nor (_06596_, _06595_, _06593_);
  nor (_06597_, _06596_, _06516_);
  and (_06598_, _06516_, word_in[12]);
  or (_06599_, _06598_, _06597_);
  and (_06600_, _06599_, _06539_);
  or (_06602_, _06600_, _06592_);
  and (_06603_, _06602_, _06537_);
  and (_06605_, _06535_, word_in[28]);
  or (_26830_[4], _06605_, _06603_);
  and (_06606_, _06022_, word_in[21]);
  and (_06607_, _06513_, _06606_);
  and (_06608_, _06523_, _06469_);
  not (_06609_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_06610_, _06523_, _06609_);
  nor (_06611_, _06610_, _06608_);
  nor (_06612_, _06611_, _06516_);
  and (_06613_, _06516_, word_in[13]);
  or (_06615_, _06613_, _06612_);
  and (_06616_, _06615_, _06539_);
  or (_06617_, _06616_, _06607_);
  and (_06618_, _06617_, _06537_);
  and (_06619_, _06535_, word_in[29]);
  or (_26830_[5], _06619_, _06618_);
  and (_06620_, _06022_, word_in[22]);
  and (_06621_, _06513_, _06620_);
  and (_06623_, _06033_, word_in[6]);
  and (_06624_, _06523_, _06623_);
  not (_06625_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_06626_, _06523_, _06625_);
  nor (_06628_, _06626_, _06624_);
  nor (_06629_, _06628_, _06516_);
  and (_06630_, _06516_, word_in[14]);
  or (_06631_, _06630_, _06629_);
  and (_06632_, _06631_, _06539_);
  or (_06633_, _06632_, _06621_);
  and (_06634_, _06633_, _06537_);
  and (_06635_, _06535_, word_in[30]);
  or (_26830_[6], _06635_, _06634_);
  and (_06636_, _06513_, _06047_);
  and (_06637_, _06523_, _06496_);
  nor (_06638_, _06523_, _05737_);
  nor (_06639_, _06638_, _06637_);
  nor (_06640_, _06639_, _06516_);
  and (_06641_, _06516_, word_in[15]);
  or (_06642_, _06641_, _06640_);
  and (_06643_, _06642_, _06539_);
  or (_06644_, _06643_, _06636_);
  and (_06645_, _06644_, _06537_);
  and (_06646_, _06535_, word_in[31]);
  or (_26830_[7], _06646_, _06645_);
  and (_06647_, _06043_, _05753_);
  and (_06648_, _06647_, _05996_);
  and (_06649_, _06022_, _05784_);
  and (_06650_, _06649_, _05876_);
  not (_06651_, _06650_);
  or (_06652_, _06651_, _06538_);
  and (_06653_, _06028_, _05751_);
  and (_06654_, _06653_, _05767_);
  not (_06655_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  not (_06656_, _06031_);
  and (_06657_, _06369_, _06656_);
  and (_06658_, _06657_, _05667_);
  nor (_06659_, _06658_, _06655_);
  and (_06660_, _06658_, _06525_);
  or (_06661_, _06660_, _06659_);
  or (_06662_, _06661_, _06654_);
  not (_06663_, _06654_);
  or (_06664_, _06663_, word_in[8]);
  and (_06665_, _06664_, _06662_);
  or (_06666_, _06665_, _06650_);
  and (_06668_, _06666_, _06652_);
  or (_06669_, _06668_, _06648_);
  not (_06670_, _06648_);
  or (_06671_, _06670_, word_in[24]);
  and (_26831_[0], _06671_, _06669_);
  and (_06672_, _06650_, _06391_);
  and (_06673_, _06658_, _06548_);
  not (_06674_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_06675_, _06658_, _06674_);
  nor (_06676_, _06675_, _06673_);
  nor (_06677_, _06676_, _06654_);
  and (_06678_, _06654_, word_in[9]);
  or (_06679_, _06678_, _06677_);
  and (_06680_, _06679_, _06651_);
  or (_06682_, _06680_, _06672_);
  and (_06683_, _06682_, _06670_);
  and (_06684_, _06648_, word_in[25]);
  or (_26831_[1], _06684_, _06683_);
  and (_06685_, _06658_, _06412_);
  not (_06686_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_06687_, _06658_, _06686_);
  nor (_06688_, _06687_, _06685_);
  nor (_06689_, _06688_, _06654_);
  and (_06690_, _06654_, word_in[10]);
  or (_06691_, _06690_, _06689_);
  and (_06692_, _06691_, _06651_);
  and (_06693_, _06650_, _06572_);
  or (_06694_, _06693_, _06648_);
  or (_06695_, _06694_, _06692_);
  or (_06696_, _06670_, word_in[26]);
  and (_26831_[2], _06696_, _06695_);
  and (_06697_, _06650_, _06586_);
  and (_06698_, _06658_, _06427_);
  not (_06699_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_06700_, _06658_, _06699_);
  nor (_06702_, _06700_, _06698_);
  nor (_06703_, _06702_, _06654_);
  and (_06704_, _06654_, word_in[11]);
  or (_06705_, _06704_, _06703_);
  and (_06706_, _06705_, _06651_);
  or (_06708_, _06706_, _06697_);
  and (_06709_, _06708_, _06670_);
  and (_06710_, _06648_, word_in[27]);
  or (_26831_[3], _06710_, _06709_);
  not (_06711_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_06712_, _06658_, _06711_);
  and (_06713_, _06658_, _06450_);
  or (_06714_, _06713_, _06712_);
  or (_06715_, _06714_, _06654_);
  or (_06716_, _06663_, word_in[12]);
  and (_06717_, _06716_, _06715_);
  or (_06718_, _06717_, _06650_);
  or (_06719_, _06651_, _06591_);
  and (_06720_, _06719_, _06670_);
  and (_06721_, _06720_, _06718_);
  and (_06723_, _06648_, word_in[28]);
  or (_26831_[4], _06723_, _06721_);
  and (_06724_, _06650_, _06606_);
  and (_06725_, _06658_, _06469_);
  not (_06726_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_06727_, _06658_, _06726_);
  nor (_06728_, _06727_, _06725_);
  nor (_06729_, _06728_, _06654_);
  and (_06730_, _06654_, word_in[13]);
  or (_06731_, _06730_, _06729_);
  and (_06733_, _06731_, _06651_);
  or (_06734_, _06733_, _06724_);
  and (_06735_, _06734_, _06670_);
  and (_06736_, _06648_, word_in[29]);
  or (_26831_[5], _06736_, _06735_);
  and (_06737_, _06658_, _06623_);
  not (_06738_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_06739_, _06658_, _06738_);
  nor (_06740_, _06739_, _06737_);
  nor (_06741_, _06740_, _06654_);
  and (_06742_, _06654_, word_in[14]);
  or (_06743_, _06742_, _06741_);
  and (_06745_, _06743_, _06651_);
  and (_06746_, _06650_, _06620_);
  or (_06747_, _06746_, _06648_);
  or (_06748_, _06747_, _06745_);
  or (_06749_, _06670_, word_in[30]);
  and (_26831_[6], _06749_, _06748_);
  and (_06750_, _06658_, _06496_);
  nor (_06751_, _06658_, _05848_);
  nor (_06753_, _06751_, _06750_);
  nor (_06754_, _06753_, _06654_);
  and (_06755_, _06654_, word_in[15]);
  or (_06756_, _06755_, _06754_);
  and (_06757_, _06756_, _06651_);
  and (_06758_, _06650_, _06047_);
  or (_06759_, _06758_, _06648_);
  or (_06761_, _06759_, _06757_);
  or (_06762_, _06670_, word_in[31]);
  and (_26831_[7], _06762_, _06761_);
  and (_06763_, _24899_, _24006_);
  and (_06764_, _06763_, _24219_);
  not (_06765_, _06763_);
  and (_06766_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or (_01925_, _06766_, _06764_);
  and (_06767_, _06022_, _05751_);
  and (_06768_, _06767_, _05876_);
  not (_06769_, _06768_);
  and (_06770_, _06029_, _05767_);
  not (_06771_, _06032_);
  nor (_06773_, _06520_, _06771_);
  and (_06774_, _06773_, _06525_);
  not (_06775_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor (_06776_, _06773_, _06775_);
  nor (_06777_, _06776_, _06774_);
  nor (_06778_, _06777_, _06770_);
  and (_06779_, _06770_, word_in[8]);
  or (_06780_, _06779_, _06778_);
  and (_06781_, _06780_, _06769_);
  and (_06782_, _06044_, _05996_);
  and (_06783_, _06768_, _06538_);
  or (_06784_, _06783_, _06782_);
  or (_06785_, _06784_, _06781_);
  not (_06786_, _06782_);
  or (_06788_, _06786_, _06364_);
  and (_26832_[0], _06788_, _06785_);
  and (_06789_, _06773_, _06548_);
  not (_06790_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_06791_, _06773_, _06790_);
  nor (_06792_, _06791_, _06789_);
  nor (_06794_, _06792_, _06770_);
  and (_06795_, _06770_, word_in[9]);
  or (_06796_, _06795_, _06794_);
  and (_06797_, _06796_, _06769_);
  and (_06798_, _06768_, _06391_);
  or (_06799_, _06798_, _06782_);
  or (_06800_, _06799_, _06797_);
  and (_06801_, _06043_, word_in[25]);
  or (_06802_, _06786_, _06801_);
  and (_26832_[1], _06802_, _06800_);
  and (_06803_, _06773_, _06412_);
  not (_06804_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_06805_, _06773_, _06804_);
  nor (_06807_, _06805_, _06803_);
  nor (_06808_, _06807_, _06770_);
  and (_06809_, _06770_, word_in[10]);
  or (_06810_, _06809_, _06808_);
  and (_06811_, _06810_, _06769_);
  and (_06812_, _06768_, _06572_);
  or (_06813_, _06812_, _06782_);
  or (_06815_, _06813_, _06811_);
  or (_06816_, _06786_, _06407_);
  and (_26832_[2], _06816_, _06815_);
  not (_06818_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_06819_, _06773_, _06818_);
  and (_06820_, _06773_, _06427_);
  or (_06821_, _06820_, _06819_);
  or (_06822_, _06821_, _06770_);
  not (_06824_, _06770_);
  or (_06825_, _06824_, word_in[11]);
  and (_06826_, _06825_, _06822_);
  or (_06827_, _06826_, _06768_);
  or (_06828_, _06769_, _06586_);
  and (_06829_, _06828_, _06786_);
  and (_06830_, _06829_, _06827_);
  and (_06831_, _06782_, _06441_);
  or (_26832_[3], _06831_, _06830_);
  not (_06832_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_06833_, _06773_, _06832_);
  and (_06834_, _06773_, _06450_);
  or (_06835_, _06834_, _06833_);
  or (_06836_, _06835_, _06770_);
  or (_06837_, _06824_, word_in[12]);
  and (_06838_, _06837_, _06836_);
  or (_06839_, _06838_, _06768_);
  or (_06840_, _06769_, _06591_);
  and (_06841_, _06840_, _06786_);
  and (_06842_, _06841_, _06839_);
  and (_06843_, _06782_, _06446_);
  or (_26832_[4], _06843_, _06842_);
  and (_06844_, _06773_, _06469_);
  not (_06845_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_06846_, _06773_, _06845_);
  nor (_06847_, _06846_, _06844_);
  nor (_06848_, _06847_, _06770_);
  and (_06849_, _06770_, word_in[13]);
  or (_06850_, _06849_, _06848_);
  and (_06851_, _06850_, _06769_);
  and (_06852_, _06768_, _06606_);
  or (_06853_, _06852_, _06782_);
  or (_06854_, _06853_, _06851_);
  or (_06855_, _06786_, _06463_);
  and (_26832_[5], _06855_, _06854_);
  and (_06856_, _06773_, _06623_);
  not (_06857_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_06858_, _06773_, _06857_);
  nor (_06859_, _06858_, _06856_);
  nor (_06860_, _06859_, _06770_);
  and (_06861_, _06770_, word_in[14]);
  or (_06862_, _06861_, _06860_);
  and (_06863_, _06862_, _06769_);
  and (_06864_, _06768_, _06620_);
  or (_06865_, _06864_, _06782_);
  or (_06866_, _06865_, _06863_);
  and (_06867_, _06043_, word_in[30]);
  or (_06868_, _06786_, _06867_);
  and (_26832_[6], _06868_, _06866_);
  and (_06870_, _06773_, _06496_);
  nor (_06871_, _06773_, _05719_);
  nor (_06872_, _06871_, _06870_);
  nor (_06873_, _06872_, _06770_);
  and (_06874_, _06770_, word_in[15]);
  or (_06875_, _06874_, _06873_);
  and (_06876_, _06875_, _06769_);
  and (_06877_, _06768_, _06047_);
  or (_06878_, _06877_, _06782_);
  or (_06879_, _06878_, _06876_);
  or (_06880_, _06786_, _06052_);
  and (_26832_[7], _06880_, _06879_);
  and (_06882_, _06043_, _06074_);
  not (_06883_, _06882_);
  not (_06884_, _05921_);
  and (_06885_, _06023_, _06884_);
  and (_06887_, _06885_, _05906_);
  and (_06888_, _06887_, _06538_);
  not (_06889_, _06887_);
  and (_06890_, _06028_, _06073_);
  not (_06891_, _06890_);
  not (_06892_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_06893_, _06033_, _05760_);
  and (_06895_, _06893_, _06370_);
  nor (_06896_, _06895_, _06892_);
  and (_06898_, _06895_, word_in[0]);
  or (_06899_, _06898_, _06896_);
  and (_06900_, _06899_, _06891_);
  and (_06901_, _06890_, word_in[8]);
  or (_06902_, _06901_, _06900_);
  and (_06903_, _06902_, _06889_);
  or (_06904_, _06903_, _06888_);
  and (_06905_, _06904_, _06883_);
  and (_06906_, _06882_, word_in[24]);
  or (_26833_[0], _06906_, _06905_);
  and (_06907_, _06887_, _06391_);
  not (_06908_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_06909_, _06895_, _06908_);
  and (_06910_, _06895_, word_in[1]);
  or (_06911_, _06910_, _06909_);
  and (_06912_, _06911_, _06891_);
  and (_06913_, _06890_, word_in[9]);
  or (_06914_, _06913_, _06912_);
  and (_06915_, _06914_, _06889_);
  or (_06916_, _06915_, _06907_);
  and (_06917_, _06916_, _06883_);
  and (_06918_, _06882_, word_in[25]);
  or (_26833_[1], _06918_, _06917_);
  and (_06919_, _06887_, _06572_);
  not (_06920_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_06921_, _06895_, _06920_);
  and (_06922_, _06895_, word_in[2]);
  or (_06924_, _06922_, _06921_);
  and (_06925_, _06924_, _06891_);
  and (_06926_, _06890_, word_in[10]);
  or (_06927_, _06926_, _06925_);
  and (_06929_, _06927_, _06889_);
  or (_06930_, _06929_, _06919_);
  and (_06931_, _06930_, _06883_);
  and (_06932_, _06882_, word_in[26]);
  or (_26833_[2], _06932_, _06931_);
  and (_06933_, _06887_, _06586_);
  not (_06934_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_06935_, _06895_, _06934_);
  and (_06936_, _06895_, word_in[3]);
  or (_06937_, _06936_, _06935_);
  and (_06938_, _06937_, _06891_);
  and (_06939_, _06890_, word_in[11]);
  or (_06940_, _06939_, _06938_);
  and (_06941_, _06940_, _06889_);
  or (_06942_, _06941_, _06933_);
  and (_06943_, _06942_, _06883_);
  and (_06944_, _06882_, word_in[27]);
  or (_26833_[3], _06944_, _06943_);
  and (_06945_, _06887_, _06591_);
  not (_06946_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_06947_, _06895_, _06946_);
  and (_06949_, _06895_, word_in[4]);
  or (_06950_, _06949_, _06947_);
  and (_06951_, _06950_, _06891_);
  and (_06952_, _06890_, word_in[12]);
  or (_06953_, _06952_, _06951_);
  and (_06954_, _06953_, _06889_);
  or (_06956_, _06954_, _06945_);
  and (_06957_, _06956_, _06883_);
  and (_06958_, _06882_, word_in[28]);
  or (_26833_[4], _06958_, _06957_);
  and (_06959_, _06887_, _06606_);
  not (_06961_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_06962_, _06895_, _06961_);
  and (_06963_, _06895_, word_in[5]);
  or (_06965_, _06963_, _06962_);
  and (_06966_, _06965_, _06891_);
  and (_06968_, _06890_, word_in[13]);
  or (_06969_, _06968_, _06966_);
  and (_06970_, _06969_, _06889_);
  or (_06971_, _06970_, _06959_);
  and (_06972_, _06971_, _06883_);
  and (_06973_, _06882_, word_in[29]);
  or (_26833_[5], _06973_, _06972_);
  and (_06975_, _06887_, _06620_);
  not (_06976_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_06977_, _06895_, _06976_);
  and (_06979_, _06895_, word_in[6]);
  or (_06981_, _06979_, _06977_);
  and (_06982_, _06981_, _06891_);
  and (_06984_, _06890_, word_in[14]);
  or (_06985_, _06984_, _06982_);
  and (_06986_, _06985_, _06889_);
  or (_06987_, _06986_, _06975_);
  and (_06989_, _06987_, _06883_);
  and (_06991_, _06882_, word_in[30]);
  or (_26833_[6], _06991_, _06989_);
  and (_06993_, _06887_, _06047_);
  nor (_06995_, _06895_, _05855_);
  and (_06996_, _06895_, word_in[7]);
  or (_06998_, _06996_, _06995_);
  and (_07000_, _06998_, _06891_);
  and (_07001_, _06890_, word_in[15]);
  or (_07002_, _07001_, _07000_);
  and (_07004_, _07002_, _06889_);
  or (_07005_, _07004_, _06993_);
  and (_07006_, _07005_, _06883_);
  and (_07007_, _06882_, word_in[31]);
  or (_26833_[7], _07007_, _07006_);
  and (_07008_, _04920_, _24219_);
  and (_07009_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_02030_, _07009_, _07008_);
  and (_07011_, _06763_, _23887_);
  and (_07012_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_02042_, _07012_, _07011_);
  and (_07013_, _24095_, _24006_);
  and (_07014_, _07013_, _23548_);
  not (_07015_, _07013_);
  and (_07016_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_02052_, _07016_, _07014_);
  and (_07017_, _06043_, _06067_);
  not (_07018_, _07017_);
  and (_07019_, _06885_, _05753_);
  and (_07020_, _07019_, _06538_);
  not (_07021_, _07019_);
  and (_07022_, _06515_, _05797_);
  not (_07023_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_07025_, _06893_, _06521_);
  nor (_07026_, _07025_, _07023_);
  and (_07027_, _07025_, word_in[0]);
  nor (_07028_, _07027_, _07026_);
  nor (_07029_, _07028_, _07022_);
  and (_07030_, _07022_, word_in[8]);
  or (_07031_, _07030_, _07029_);
  and (_07032_, _07031_, _07021_);
  or (_07034_, _07032_, _07020_);
  and (_07035_, _07034_, _07018_);
  and (_07036_, _07017_, word_in[24]);
  or (_26834_[0], _07036_, _07035_);
  and (_07038_, _24349_, _24301_);
  and (_07040_, _07038_, _23996_);
  not (_07041_, _07038_);
  and (_07042_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_27227_, _07042_, _07040_);
  and (_07044_, _07019_, _06391_);
  and (_07045_, _07025_, word_in[1]);
  not (_07046_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_07048_, _07025_, _07046_);
  nor (_07050_, _07048_, _07045_);
  nor (_07052_, _07050_, _07022_);
  and (_07053_, _07022_, word_in[9]);
  or (_07055_, _07053_, _07052_);
  and (_07056_, _07055_, _07021_);
  or (_07057_, _07056_, _07044_);
  and (_07058_, _07057_, _07018_);
  and (_07060_, _07017_, word_in[25]);
  or (_26834_[1], _07060_, _07058_);
  and (_07062_, _07017_, word_in[26]);
  not (_07063_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_07064_, _07025_, _07063_);
  and (_07065_, _07025_, _06412_);
  or (_07066_, _07065_, _07064_);
  or (_07067_, _07066_, _07022_);
  not (_07068_, _07022_);
  or (_07069_, _07068_, word_in[10]);
  and (_07070_, _07069_, _07067_);
  or (_07071_, _07070_, _07019_);
  or (_07073_, _07021_, _06572_);
  and (_07074_, _07073_, _07018_);
  and (_07076_, _07074_, _07071_);
  or (_26834_[2], _07076_, _07062_);
  and (_07077_, _07017_, word_in[27]);
  not (_07078_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_07079_, _07025_, _07078_);
  and (_07080_, _07025_, _06427_);
  or (_07082_, _07080_, _07079_);
  or (_07084_, _07082_, _07022_);
  or (_07085_, _07068_, word_in[11]);
  and (_07086_, _07085_, _07084_);
  or (_07087_, _07086_, _07019_);
  or (_07088_, _07021_, _06586_);
  and (_07090_, _07088_, _07018_);
  and (_07091_, _07090_, _07087_);
  or (_26834_[3], _07091_, _07077_);
  and (_07093_, _07019_, _06591_);
  and (_07095_, _07025_, word_in[4]);
  not (_07096_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_07097_, _07025_, _07096_);
  nor (_07098_, _07097_, _07095_);
  nor (_07099_, _07098_, _07022_);
  and (_07101_, _07022_, word_in[12]);
  or (_07102_, _07101_, _07099_);
  and (_07104_, _07102_, _07021_);
  or (_07105_, _07104_, _07093_);
  and (_07106_, _07105_, _07018_);
  and (_07108_, _07017_, word_in[28]);
  or (_26834_[4], _07108_, _07106_);
  and (_07110_, _07017_, word_in[29]);
  and (_07111_, _07025_, word_in[5]);
  not (_07112_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_07114_, _07025_, _07112_);
  nor (_07116_, _07114_, _07111_);
  nor (_07118_, _07116_, _07022_);
  and (_07119_, _07022_, word_in[13]);
  or (_07120_, _07119_, _07118_);
  or (_07121_, _07120_, _07019_);
  or (_07122_, _07021_, _06606_);
  and (_07124_, _07122_, _07018_);
  and (_07126_, _07124_, _07121_);
  or (_26834_[5], _07126_, _07110_);
  not (_07127_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_07128_, _07025_, _07127_);
  and (_07129_, _07025_, word_in[6]);
  nor (_07131_, _07129_, _07128_);
  nor (_07132_, _07131_, _07022_);
  and (_07133_, _07022_, word_in[14]);
  or (_07134_, _07133_, _07132_);
  and (_07136_, _07134_, _07021_);
  and (_07137_, _07019_, _06620_);
  or (_07138_, _07137_, _07136_);
  and (_07139_, _07138_, _07018_);
  and (_07140_, _07017_, word_in[30]);
  or (_26834_[6], _07140_, _07139_);
  and (_07142_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and (_07143_, _06203_, _23887_);
  or (_02081_, _07143_, _07142_);
  and (_07144_, _07019_, _06047_);
  nor (_07146_, _07025_, _05732_);
  and (_07147_, _07025_, word_in[7]);
  nor (_07148_, _07147_, _07146_);
  nor (_07149_, _07148_, _07022_);
  and (_07150_, _07022_, word_in[15]);
  or (_07151_, _07150_, _07149_);
  and (_07152_, _07151_, _07021_);
  or (_07153_, _07152_, _07144_);
  and (_07154_, _07153_, _07018_);
  and (_07155_, _07017_, word_in[31]);
  or (_26834_[7], _07155_, _07154_);
  and (_07157_, _06129_, _24089_);
  and (_07158_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  or (_02099_, _07158_, _07157_);
  and (_07159_, _07013_, _23583_);
  and (_07160_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_02128_, _07160_, _07159_);
  and (_07161_, _06043_, _06073_);
  not (_07162_, _07161_);
  and (_07163_, _06885_, _05784_);
  and (_07165_, _07163_, _06538_);
  not (_07166_, _07163_);
  and (_07167_, _06653_, _05797_);
  and (_07168_, _06657_, _05760_);
  and (_07169_, _07168_, word_in[0]);
  not (_07170_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor (_07171_, _07168_, _07170_);
  nor (_07172_, _07171_, _07169_);
  nor (_07173_, _07172_, _07167_);
  and (_07174_, _07167_, word_in[8]);
  or (_07175_, _07174_, _07173_);
  and (_07176_, _07175_, _07166_);
  or (_07178_, _07176_, _07165_);
  and (_07179_, _07178_, _07162_);
  and (_07181_, _07161_, word_in[24]);
  or (_26835_[0], _07181_, _07179_);
  and (_07182_, _07163_, _06391_);
  not (_07183_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_07184_, _07168_, _07183_);
  and (_07186_, _07168_, word_in[1]);
  nor (_07187_, _07186_, _07184_);
  nor (_07189_, _07187_, _07167_);
  and (_07190_, _07167_, word_in[9]);
  or (_07191_, _07190_, _07189_);
  and (_07192_, _07191_, _07166_);
  or (_07193_, _07192_, _07182_);
  and (_07195_, _07193_, _07162_);
  and (_07196_, _07161_, word_in[25]);
  or (_26835_[1], _07196_, _07195_);
  and (_07198_, _06763_, _23548_);
  and (_07200_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_02151_, _07200_, _07198_);
  and (_07202_, _07163_, _06572_);
  not (_07203_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_07205_, _07168_, _07203_);
  and (_07206_, _07168_, word_in[2]);
  nor (_07207_, _07206_, _07205_);
  nor (_07208_, _07207_, _07167_);
  and (_07209_, _07167_, word_in[10]);
  or (_07210_, _07209_, _07208_);
  and (_07211_, _07210_, _07166_);
  or (_07212_, _07211_, _07202_);
  and (_07213_, _07212_, _07162_);
  and (_07215_, _07161_, word_in[26]);
  or (_26835_[2], _07215_, _07213_);
  and (_07217_, _07163_, _06586_);
  not (_07218_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_07219_, _07168_, _07218_);
  and (_07220_, _07168_, word_in[3]);
  nor (_07222_, _07220_, _07219_);
  nor (_07224_, _07222_, _07167_);
  and (_07225_, _07167_, word_in[11]);
  or (_07227_, _07225_, _07224_);
  and (_07228_, _07227_, _07166_);
  or (_07229_, _07228_, _07217_);
  and (_07230_, _07229_, _07162_);
  and (_07231_, _07161_, word_in[27]);
  or (_26835_[3], _07231_, _07230_);
  and (_07233_, _07163_, _06591_);
  not (_07234_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_07235_, _07168_, _07234_);
  and (_07236_, _07168_, word_in[4]);
  nor (_07237_, _07236_, _07235_);
  nor (_07238_, _07237_, _07167_);
  and (_07239_, _07167_, word_in[12]);
  or (_07240_, _07239_, _07238_);
  and (_07241_, _07240_, _07166_);
  or (_07242_, _07241_, _07233_);
  and (_07243_, _07242_, _07162_);
  and (_07244_, _07161_, word_in[28]);
  or (_26835_[4], _07244_, _07243_);
  and (_07246_, _07163_, _06606_);
  not (_07247_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_07248_, _07168_, _07247_);
  and (_07249_, _07168_, word_in[5]);
  nor (_07250_, _07249_, _07248_);
  nor (_07252_, _07250_, _07167_);
  and (_07253_, _07167_, word_in[13]);
  or (_07254_, _07253_, _07252_);
  and (_07255_, _07254_, _07166_);
  or (_07256_, _07255_, _07246_);
  and (_07257_, _07256_, _07162_);
  and (_07258_, _07161_, word_in[29]);
  or (_26835_[5], _07258_, _07257_);
  and (_07259_, _07163_, _06620_);
  not (_07260_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_07261_, _07168_, _07260_);
  and (_07262_, _07168_, word_in[6]);
  nor (_07263_, _07262_, _07261_);
  nor (_07264_, _07263_, _07167_);
  and (_07265_, _07167_, word_in[14]);
  or (_07267_, _07265_, _07264_);
  and (_07268_, _07267_, _07166_);
  or (_07269_, _07268_, _07259_);
  and (_07271_, _07269_, _07162_);
  and (_07272_, _07161_, word_in[30]);
  or (_26835_[6], _07272_, _07271_);
  and (_07273_, _07163_, _06047_);
  nor (_07274_, _07168_, _05862_);
  and (_07275_, _07168_, word_in[7]);
  nor (_07277_, _07275_, _07274_);
  nor (_07278_, _07277_, _07167_);
  and (_07279_, _07167_, word_in[15]);
  or (_07280_, _07279_, _07278_);
  and (_07281_, _07280_, _07166_);
  or (_07282_, _07281_, _07273_);
  and (_07283_, _07282_, _07162_);
  and (_07284_, _07161_, word_in[31]);
  or (_26835_[7], _07284_, _07283_);
  and (_07285_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and (_07286_, _06203_, _23548_);
  or (_02165_, _07286_, _07285_);
  and (_07287_, _06043_, _06080_);
  and (_07288_, _07287_, word_in[24]);
  and (_07289_, _06885_, _05751_);
  and (_07290_, _06029_, _05797_);
  and (_07291_, _06893_, _06032_);
  and (_07292_, _07291_, word_in[0]);
  not (_07294_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor (_07295_, _07291_, _07294_);
  nor (_07296_, _07295_, _07292_);
  nor (_07298_, _07296_, _07290_);
  and (_07299_, _07290_, word_in[8]);
  or (_07301_, _07299_, _07298_);
  or (_07302_, _07301_, _07289_);
  not (_07303_, _07287_);
  not (_07304_, _07289_);
  or (_07305_, _07304_, _06538_);
  and (_07307_, _07305_, _07303_);
  and (_07308_, _07307_, _07302_);
  or (_26836_[0], _07308_, _07288_);
  not (_07310_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_07311_, _07291_, _07310_);
  and (_07312_, _07291_, _06548_);
  or (_07313_, _07312_, _07311_);
  or (_07314_, _07313_, _07290_);
  not (_07315_, _07290_);
  or (_07316_, _07315_, word_in[9]);
  and (_07318_, _07316_, _07314_);
  or (_07319_, _07318_, _07289_);
  or (_07320_, _07304_, _06391_);
  and (_07321_, _07320_, _07303_);
  and (_07322_, _07321_, _07319_);
  and (_07323_, _07287_, word_in[25]);
  or (_26836_[1], _07323_, _07322_);
  and (_07325_, _07287_, word_in[26]);
  or (_07326_, _07304_, _06572_);
  and (_07327_, _07326_, _07303_);
  and (_07328_, _07291_, word_in[2]);
  not (_07329_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_07330_, _07291_, _07329_);
  nor (_07331_, _07330_, _07328_);
  nor (_07332_, _07331_, _07290_);
  and (_07333_, _07290_, word_in[10]);
  or (_07334_, _07333_, _07332_);
  or (_07335_, _07334_, _07289_);
  and (_07336_, _07335_, _07327_);
  or (_26836_[2], _07336_, _07325_);
  and (_07337_, _07287_, word_in[27]);
  not (_07339_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_07340_, _07291_, _07339_);
  and (_07342_, _07291_, _06427_);
  or (_07343_, _07342_, _07340_);
  or (_07345_, _07343_, _07290_);
  or (_07347_, _07315_, word_in[11]);
  and (_07348_, _07347_, _07345_);
  or (_07350_, _07348_, _07289_);
  or (_07351_, _07304_, _06586_);
  and (_07352_, _07351_, _07303_);
  and (_07354_, _07352_, _07350_);
  or (_26836_[3], _07354_, _07337_);
  and (_07356_, _07287_, word_in[28]);
  not (_07357_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_07358_, _07291_, _07357_);
  and (_07359_, _07291_, _06450_);
  or (_07361_, _07359_, _07358_);
  or (_07362_, _07361_, _07290_);
  or (_07363_, _07315_, word_in[12]);
  and (_07364_, _07363_, _07362_);
  or (_07365_, _07364_, _07289_);
  or (_07367_, _07304_, _06591_);
  and (_07368_, _07367_, _07303_);
  and (_07369_, _07368_, _07365_);
  or (_26836_[4], _07369_, _07356_);
  and (_07371_, _07287_, word_in[29]);
  or (_07372_, _07304_, _06606_);
  and (_07373_, _07372_, _07303_);
  and (_07374_, _07291_, word_in[5]);
  not (_07375_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_07376_, _07291_, _07375_);
  nor (_07377_, _07376_, _07374_);
  nor (_07378_, _07377_, _07290_);
  and (_07379_, _07290_, word_in[13]);
  or (_07380_, _07379_, _07378_);
  or (_07381_, _07380_, _07289_);
  and (_07382_, _07381_, _07373_);
  or (_26836_[5], _07382_, _07371_);
  and (_07383_, _07287_, word_in[30]);
  not (_07384_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_07385_, _07291_, _07384_);
  and (_07387_, _07291_, word_in[6]);
  nor (_07388_, _07387_, _07385_);
  nor (_07389_, _07388_, _07290_);
  and (_07390_, _07290_, word_in[14]);
  or (_07392_, _07390_, _07389_);
  and (_07393_, _07392_, _07304_);
  and (_07395_, _07289_, _06620_);
  or (_07396_, _07395_, _07393_);
  and (_07398_, _07396_, _07303_);
  or (_26836_[6], _07398_, _07383_);
  nor (_07400_, _07291_, _05726_);
  and (_07401_, _07291_, _06496_);
  or (_07402_, _07401_, _07400_);
  or (_07404_, _07402_, _07290_);
  or (_07405_, _07315_, word_in[15]);
  and (_07406_, _07405_, _07404_);
  or (_07408_, _07406_, _07289_);
  or (_07410_, _07304_, _06047_);
  and (_07411_, _07410_, _07303_);
  and (_07412_, _07411_, _07408_);
  and (_07413_, _07287_, word_in[31]);
  or (_26836_[7], _07413_, _07412_);
  and (_07415_, _07013_, _23887_);
  and (_07416_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_02261_, _07416_, _07415_);
  and (_07417_, _06043_, _05957_);
  and (_07419_, _07417_, _05751_);
  not (_07420_, _07419_);
  and (_07421_, _06022_, _06105_);
  and (_07422_, _07421_, word_in[16]);
  not (_07423_, _07421_);
  and (_07424_, _06028_, _05761_);
  not (_07426_, _07424_);
  not (_07428_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_07429_, _06033_, _05669_);
  and (_07430_, _07429_, _06370_);
  nor (_07431_, _07430_, _07428_);
  and (_07432_, _07430_, word_in[0]);
  or (_07434_, _07432_, _07431_);
  and (_07435_, _07434_, _07426_);
  and (_07436_, _07424_, word_in[8]);
  or (_07437_, _07436_, _07435_);
  and (_07438_, _07437_, _07423_);
  or (_07439_, _07438_, _07422_);
  and (_07440_, _07439_, _07420_);
  and (_07441_, _07419_, word_in[24]);
  or (_26837_[0], _07441_, _07440_);
  and (_07442_, _07421_, word_in[17]);
  not (_07443_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_07445_, _07430_, _07443_);
  and (_07446_, _07430_, word_in[1]);
  or (_07447_, _07446_, _07445_);
  and (_07448_, _07447_, _07426_);
  and (_07450_, _07424_, word_in[9]);
  or (_07451_, _07450_, _07448_);
  and (_07452_, _07451_, _07423_);
  or (_07453_, _07452_, _07442_);
  and (_07454_, _07453_, _07420_);
  and (_07455_, _07419_, word_in[25]);
  or (_26837_[1], _07455_, _07454_);
  and (_07457_, _07421_, word_in[18]);
  not (_07458_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_07459_, _07430_, _07458_);
  and (_07460_, _07430_, word_in[2]);
  or (_07461_, _07460_, _07459_);
  and (_07463_, _07461_, _07426_);
  and (_07464_, _07424_, word_in[10]);
  or (_07465_, _07464_, _07463_);
  and (_07466_, _07465_, _07423_);
  or (_07467_, _07466_, _07457_);
  and (_07468_, _07467_, _07420_);
  and (_07470_, _07419_, word_in[26]);
  or (_26837_[2], _07470_, _07468_);
  and (_07472_, _07421_, word_in[19]);
  not (_07473_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_07474_, _07430_, _07473_);
  and (_07475_, _07430_, word_in[3]);
  or (_07476_, _07475_, _07474_);
  and (_07477_, _07476_, _07426_);
  and (_07478_, _07424_, word_in[11]);
  or (_07480_, _07478_, _07477_);
  and (_07481_, _07480_, _07423_);
  or (_07482_, _07481_, _07472_);
  and (_07483_, _07482_, _07420_);
  and (_07484_, _07419_, word_in[27]);
  or (_26837_[3], _07484_, _07483_);
  and (_07485_, _07421_, word_in[20]);
  not (_07486_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_07487_, _07430_, _07486_);
  and (_07488_, _07430_, word_in[4]);
  or (_07489_, _07488_, _07487_);
  and (_07490_, _07489_, _07426_);
  and (_07491_, _07424_, word_in[12]);
  or (_07492_, _07491_, _07490_);
  and (_07493_, _07492_, _07423_);
  or (_07494_, _07493_, _07485_);
  and (_07495_, _07494_, _07420_);
  and (_07496_, _07419_, word_in[28]);
  or (_26837_[4], _07496_, _07495_);
  and (_07497_, _07421_, word_in[21]);
  not (_07498_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_07500_, _07430_, _07498_);
  and (_07502_, _07430_, word_in[5]);
  or (_07504_, _07502_, _07500_);
  and (_07505_, _07504_, _07426_);
  and (_07507_, _07424_, word_in[13]);
  or (_07508_, _07507_, _07505_);
  and (_07509_, _07508_, _07423_);
  or (_07510_, _07509_, _07497_);
  and (_07512_, _07510_, _07420_);
  and (_07514_, _07419_, word_in[29]);
  or (_26837_[5], _07514_, _07512_);
  and (_07516_, _07421_, word_in[22]);
  not (_07517_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_07518_, _07430_, _07517_);
  and (_07519_, _07430_, word_in[6]);
  or (_07520_, _07519_, _07518_);
  and (_07521_, _07520_, _07426_);
  and (_07522_, _07424_, word_in[14]);
  or (_07523_, _07522_, _07521_);
  and (_07524_, _07523_, _07423_);
  or (_07525_, _07524_, _07516_);
  and (_07526_, _07525_, _07420_);
  and (_07527_, _07419_, word_in[30]);
  or (_26837_[6], _07527_, _07526_);
  and (_07529_, _07421_, word_in[23]);
  nor (_07530_, _07430_, _05832_);
  and (_07531_, _07430_, word_in[7]);
  or (_07532_, _07531_, _07530_);
  and (_07533_, _07532_, _07426_);
  and (_07534_, _07424_, word_in[15]);
  or (_07536_, _07534_, _07533_);
  and (_07537_, _07536_, _07423_);
  or (_07538_, _07537_, _07529_);
  and (_07539_, _07538_, _07420_);
  and (_07541_, _07419_, word_in[31]);
  or (_26837_[7], _07541_, _07539_);
  and (_07543_, _04920_, _23887_);
  and (_07545_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_02327_, _07545_, _07543_);
  and (_07547_, _24497_, _24219_);
  and (_07548_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  or (_02342_, _07548_, _07547_);
  and (_07549_, _06043_, _06105_);
  and (_07551_, _06512_, _05885_);
  not (_07552_, _07551_);
  or (_07553_, _07552_, word_in[16]);
  and (_07555_, _06515_, _05763_);
  not (_07556_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_07557_, _07429_, _06521_);
  nor (_07559_, _07557_, _07556_);
  and (_07560_, _07557_, _06525_);
  or (_07561_, _07560_, _07559_);
  or (_07563_, _07561_, _07555_);
  not (_07564_, _07555_);
  or (_07566_, _07564_, word_in[8]);
  and (_07567_, _07566_, _07563_);
  or (_07568_, _07567_, _07551_);
  and (_07569_, _07568_, _07553_);
  or (_07570_, _07569_, _07549_);
  not (_07571_, _07549_);
  or (_07572_, _07571_, word_in[24]);
  and (_26838_[0], _07572_, _07570_);
  not (_07573_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_07574_, _07557_, _07573_);
  and (_07575_, _07557_, _06548_);
  or (_07576_, _07575_, _07574_);
  or (_07578_, _07576_, _07555_);
  or (_07579_, _07564_, word_in[9]);
  and (_07581_, _07579_, _07578_);
  or (_07582_, _07581_, _07551_);
  or (_07583_, _07552_, word_in[17]);
  and (_07584_, _07583_, _07571_);
  and (_07585_, _07584_, _07582_);
  and (_07587_, _07549_, word_in[25]);
  or (_26838_[1], _07587_, _07585_);
  and (_07589_, _07551_, word_in[18]);
  not (_07590_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_07591_, _07557_, _07590_);
  and (_07592_, _07557_, word_in[2]);
  nor (_07593_, _07592_, _07591_);
  nor (_07594_, _07593_, _07555_);
  and (_07595_, _07555_, word_in[10]);
  or (_07596_, _07595_, _07594_);
  and (_07597_, _07596_, _07552_);
  or (_07598_, _07597_, _07589_);
  and (_07599_, _07598_, _07571_);
  and (_07600_, _07549_, word_in[26]);
  or (_26838_[2], _07600_, _07599_);
  and (_07601_, _07551_, word_in[19]);
  not (_07602_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_07604_, _07557_, _07602_);
  and (_07605_, _07557_, word_in[3]);
  nor (_07606_, _07605_, _07604_);
  nor (_07608_, _07606_, _07555_);
  and (_07609_, _07555_, word_in[11]);
  or (_07610_, _07609_, _07608_);
  and (_07611_, _07610_, _07552_);
  or (_07612_, _07611_, _07601_);
  and (_07613_, _07612_, _07571_);
  and (_07615_, _07549_, word_in[27]);
  or (_26838_[3], _07615_, _07613_);
  not (_07616_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_07617_, _07557_, _07616_);
  and (_07618_, _07557_, _06450_);
  or (_07619_, _07618_, _07617_);
  or (_07620_, _07619_, _07555_);
  or (_07621_, _07564_, word_in[12]);
  and (_07622_, _07621_, _07620_);
  or (_07623_, _07622_, _07551_);
  or (_07625_, _07552_, _06591_);
  and (_07627_, _07625_, _07571_);
  and (_07628_, _07627_, _07623_);
  and (_07629_, _07549_, word_in[28]);
  or (_26838_[4], _07629_, _07628_);
  or (_07630_, _07552_, word_in[21]);
  not (_07631_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_07632_, _07557_, _07631_);
  and (_07633_, _07557_, _06469_);
  or (_07634_, _07633_, _07632_);
  or (_07635_, _07634_, _07555_);
  or (_07636_, _07564_, word_in[13]);
  and (_07637_, _07636_, _07635_);
  or (_07638_, _07637_, _07551_);
  and (_07640_, _07638_, _07630_);
  and (_07641_, _07640_, _07571_);
  and (_07642_, _07549_, word_in[29]);
  or (_26838_[5], _07642_, _07641_);
  and (_07643_, _07551_, word_in[22]);
  and (_07644_, _07557_, word_in[6]);
  not (_07647_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_07649_, _07557_, _07647_);
  nor (_07650_, _07649_, _07644_);
  nor (_07651_, _07650_, _07555_);
  and (_07652_, _07555_, word_in[14]);
  or (_07653_, _07652_, _07651_);
  and (_07654_, _07653_, _07552_);
  or (_07655_, _07654_, _07643_);
  and (_07656_, _07655_, _07571_);
  and (_07657_, _07549_, word_in[30]);
  or (_26838_[6], _07657_, _07656_);
  nor (_07658_, _07557_, _05709_);
  and (_07659_, _07557_, _06496_);
  or (_07660_, _07659_, _07658_);
  or (_07661_, _07660_, _07555_);
  or (_07662_, _07564_, word_in[15]);
  and (_07663_, _07662_, _07661_);
  or (_07664_, _07663_, _07551_);
  or (_07665_, _07552_, _06047_);
  and (_07666_, _07665_, _07571_);
  and (_07667_, _07666_, _07664_);
  and (_07668_, _07549_, word_in[31]);
  or (_26838_[7], _07668_, _07667_);
  nor (_26841_[2], _26684_, rst);
  and (_07669_, _06647_, _05957_);
  and (_07670_, _06649_, _05885_);
  not (_07671_, _07670_);
  or (_07672_, _07671_, _06538_);
  and (_07673_, _06653_, _05763_);
  not (_07674_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_07675_, _06657_, _05669_);
  nor (_07676_, _07675_, _07674_);
  and (_07677_, _07675_, word_in[0]);
  or (_07678_, _07677_, _07676_);
  or (_07679_, _07678_, _07673_);
  not (_07680_, _07673_);
  or (_07681_, _07680_, word_in[8]);
  and (_07682_, _07681_, _07679_);
  or (_07683_, _07682_, _07670_);
  and (_07684_, _07683_, _07672_);
  or (_07685_, _07684_, _07669_);
  not (_07686_, _07669_);
  or (_07687_, _07686_, word_in[24]);
  and (_26824_[0], _07687_, _07685_);
  not (_07688_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_07689_, _07675_, _07688_);
  and (_07690_, _07675_, word_in[1]);
  or (_07691_, _07690_, _07689_);
  or (_07692_, _07691_, _07673_);
  or (_07693_, _07680_, word_in[9]);
  and (_07694_, _07693_, _07692_);
  or (_07695_, _07694_, _07670_);
  or (_07696_, _07671_, _06391_);
  and (_07697_, _07696_, _07686_);
  and (_07698_, _07697_, _07695_);
  and (_07699_, _07669_, word_in[25]);
  or (_26824_[1], _07699_, _07698_);
  not (_07700_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_07701_, _07675_, _07700_);
  and (_07702_, _07675_, word_in[2]);
  or (_07704_, _07702_, _07701_);
  or (_07705_, _07704_, _07673_);
  or (_07706_, _07680_, word_in[10]);
  and (_07707_, _07706_, _07705_);
  or (_07708_, _07707_, _07670_);
  or (_07709_, _07671_, _06572_);
  and (_07710_, _07709_, _07686_);
  and (_07711_, _07710_, _07708_);
  and (_07712_, _07669_, word_in[26]);
  or (_26824_[2], _07712_, _07711_);
  or (_07713_, _07671_, _06586_);
  not (_07714_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_07715_, _07675_, _07714_);
  and (_07716_, _07675_, word_in[3]);
  or (_07717_, _07716_, _07715_);
  or (_07718_, _07717_, _07673_);
  or (_07719_, _07680_, word_in[11]);
  and (_07720_, _07719_, _07718_);
  or (_07721_, _07720_, _07670_);
  and (_07722_, _07721_, _07713_);
  or (_07724_, _07722_, _07669_);
  or (_07725_, _07686_, word_in[27]);
  and (_26824_[3], _07725_, _07724_);
  not (_07726_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_07727_, _07675_, _07726_);
  and (_07728_, _07675_, word_in[4]);
  or (_07729_, _07728_, _07727_);
  or (_07730_, _07729_, _07673_);
  or (_07731_, _07680_, word_in[12]);
  and (_07732_, _07731_, _07730_);
  or (_07733_, _07732_, _07670_);
  or (_07734_, _07671_, _06591_);
  and (_07735_, _07734_, _07686_);
  and (_07736_, _07735_, _07733_);
  and (_07737_, _07669_, word_in[28]);
  or (_26824_[4], _07737_, _07736_);
  not (_07738_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_07739_, _07675_, _07738_);
  and (_07740_, _07675_, word_in[5]);
  or (_07741_, _07740_, _07739_);
  or (_07743_, _07741_, _07673_);
  or (_07744_, _07680_, word_in[13]);
  and (_07745_, _07744_, _07743_);
  or (_07746_, _07745_, _07670_);
  or (_07747_, _07671_, _06606_);
  and (_07748_, _07747_, _07686_);
  and (_07749_, _07748_, _07746_);
  and (_07750_, _07669_, word_in[29]);
  or (_26824_[5], _07750_, _07749_);
  or (_07751_, _07671_, _06620_);
  not (_07752_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_07753_, _07675_, _07752_);
  and (_07754_, _07675_, word_in[6]);
  or (_07755_, _07754_, _07753_);
  or (_07756_, _07755_, _07673_);
  or (_07757_, _07680_, word_in[14]);
  and (_07758_, _07757_, _07756_);
  or (_07759_, _07758_, _07670_);
  and (_07760_, _07759_, _07751_);
  or (_07761_, _07760_, _07669_);
  or (_07763_, _07686_, word_in[30]);
  and (_26824_[6], _07763_, _07761_);
  nor (_07764_, _07675_, _05827_);
  and (_07765_, _07675_, word_in[7]);
  or (_07766_, _07765_, _07764_);
  or (_07767_, _07766_, _07673_);
  or (_07768_, _07680_, word_in[15]);
  and (_07769_, _07768_, _07767_);
  or (_07770_, _07769_, _07670_);
  or (_07771_, _07671_, _06047_);
  and (_07772_, _07771_, _07686_);
  and (_07773_, _07772_, _07770_);
  and (_07774_, _07669_, word_in[31]);
  or (_26824_[7], _07774_, _07773_);
  and (_07775_, _25414_, _23887_);
  and (_07776_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_02454_, _07776_, _07775_);
  and (_07777_, _25414_, _24219_);
  and (_07778_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or (_02457_, _07778_, _07777_);
  and (_07779_, _25413_, _24140_);
  and (_07780_, _07779_, _23996_);
  not (_07781_, _07779_);
  and (_07782_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  or (_27158_, _07782_, _07780_);
  and (_07783_, _07779_, _23583_);
  and (_07784_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  or (_02464_, _07784_, _07783_);
  and (_07785_, _07779_, _23548_);
  and (_07786_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  or (_02466_, _07786_, _07785_);
  and (_07787_, _02368_, _24089_);
  and (_07788_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  or (_27151_, _07788_, _07787_);
  and (_07789_, _02368_, _23887_);
  and (_07790_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  or (_02477_, _07790_, _07789_);
  and (_07791_, _02413_, _24051_);
  and (_07792_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_02482_, _07792_, _07791_);
  and (_07793_, _06767_, _05885_);
  and (_07794_, _06029_, _05763_);
  not (_07795_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_07796_, _07429_, _06032_);
  nor (_07797_, _07796_, _07795_);
  and (_07798_, _07796_, _06525_);
  or (_07799_, _07798_, _07797_);
  or (_07800_, _07799_, _07794_);
  not (_07801_, word_in[8]);
  nand (_07802_, _07794_, _07801_);
  and (_07803_, _07802_, _07800_);
  or (_07804_, _07803_, _07793_);
  and (_07805_, _06044_, _05957_);
  not (_07806_, _07805_);
  not (_07807_, _07793_);
  or (_07808_, _07807_, word_in[16]);
  and (_07809_, _07808_, _07806_);
  and (_07810_, _07809_, _07804_);
  and (_07811_, _07805_, _06364_);
  or (_26825_[0], _07811_, _07810_);
  and (_07813_, _02413_, _23583_);
  and (_07814_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_02487_, _07814_, _07813_);
  and (_07815_, _07796_, word_in[1]);
  not (_07816_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_07817_, _07796_, _07816_);
  nor (_07818_, _07817_, _07815_);
  nor (_07819_, _07818_, _07794_);
  and (_07820_, _07794_, word_in[9]);
  or (_07821_, _07820_, _07819_);
  and (_07822_, _07821_, _07807_);
  and (_07823_, _07793_, word_in[17]);
  or (_07824_, _07823_, _07805_);
  or (_07825_, _07824_, _07822_);
  or (_07826_, _07806_, _06801_);
  and (_26825_[1], _07826_, _07825_);
  and (_07827_, _07796_, word_in[2]);
  not (_07828_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_07829_, _07796_, _07828_);
  nor (_07830_, _07829_, _07827_);
  nor (_07831_, _07830_, _07794_);
  and (_07832_, _07794_, word_in[10]);
  or (_07833_, _07832_, _07831_);
  and (_07834_, _07833_, _07807_);
  and (_07835_, _07793_, word_in[18]);
  or (_07836_, _07835_, _07805_);
  or (_07837_, _07836_, _07834_);
  or (_07838_, _07806_, _06407_);
  and (_26825_[2], _07838_, _07837_);
  and (_07839_, _07796_, word_in[3]);
  not (_07840_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_07841_, _07796_, _07840_);
  nor (_07842_, _07841_, _07839_);
  nor (_07843_, _07842_, _07794_);
  and (_07844_, _07794_, word_in[11]);
  or (_07845_, _07844_, _07843_);
  and (_07846_, _07845_, _07807_);
  and (_07847_, _07793_, word_in[19]);
  or (_07848_, _07847_, _07846_);
  and (_07849_, _07848_, _07806_);
  and (_07850_, _07805_, word_in[27]);
  or (_26825_[3], _07850_, _07849_);
  and (_07851_, _02455_, _24051_);
  and (_07852_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_02493_, _07852_, _07851_);
  and (_07853_, _07796_, word_in[4]);
  not (_07854_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_07855_, _07796_, _07854_);
  nor (_07856_, _07855_, _07853_);
  nor (_07857_, _07856_, _07794_);
  and (_07858_, _07794_, word_in[12]);
  or (_07859_, _07858_, _07857_);
  and (_07860_, _07859_, _07807_);
  and (_07861_, _07793_, _06591_);
  or (_07862_, _07861_, _07860_);
  and (_07863_, _07862_, _07806_);
  and (_07864_, _07805_, word_in[28]);
  or (_26825_[4], _07864_, _07863_);
  and (_07865_, _02455_, _23583_);
  and (_07866_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_02496_, _07866_, _07865_);
  and (_07867_, _07796_, word_in[5]);
  not (_07869_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_07871_, _07796_, _07869_);
  nor (_07872_, _07871_, _07867_);
  nor (_07873_, _07872_, _07794_);
  and (_07874_, _07794_, word_in[13]);
  or (_07876_, _07874_, _07873_);
  and (_07878_, _07876_, _07807_);
  and (_07880_, _07793_, word_in[21]);
  or (_07882_, _07880_, _07805_);
  or (_07883_, _07882_, _07878_);
  or (_07885_, _07806_, _06463_);
  and (_26825_[5], _07885_, _07883_);
  and (_07886_, _07796_, word_in[6]);
  not (_07887_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_07888_, _07796_, _07887_);
  nor (_07890_, _07888_, _07886_);
  nor (_07892_, _07890_, _07794_);
  and (_07893_, _07794_, word_in[14]);
  or (_07895_, _07893_, _07892_);
  and (_07897_, _07895_, _07807_);
  and (_07899_, _07793_, word_in[22]);
  or (_07900_, _07899_, _07805_);
  or (_07901_, _07900_, _07897_);
  or (_07903_, _07806_, _06867_);
  and (_26825_[6], _07903_, _07901_);
  and (_07906_, _07796_, word_in[7]);
  nor (_07907_, _07796_, _05697_);
  nor (_07909_, _07907_, _07906_);
  nor (_07911_, _07909_, _07794_);
  and (_07913_, _07794_, word_in[15]);
  or (_07915_, _07913_, _07911_);
  and (_07916_, _07915_, _07807_);
  and (_07918_, _07793_, _06047_);
  or (_07919_, _07918_, _07916_);
  and (_07920_, _07919_, _07806_);
  and (_07921_, _07805_, word_in[31]);
  or (_26825_[7], _07921_, _07920_);
  and (_07922_, _02517_, _24134_);
  and (_07924_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  or (_02506_, _07924_, _07922_);
  and (_07925_, _02517_, _24089_);
  and (_07926_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  or (_02510_, _07926_, _07925_);
  and (_07927_, _02890_, _23583_);
  and (_07928_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  or (_02529_, _07928_, _07927_);
  and (_07929_, _04865_, _23996_);
  and (_07930_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or (_02533_, _07930_, _07929_);
  and (_07931_, _04812_, _24089_);
  and (_07932_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_02538_, _07932_, _07931_);
  and (_07933_, _05431_, _23887_);
  and (_07934_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  or (_27129_, _07934_, _07933_);
  and (_07935_, _05431_, _24219_);
  and (_07936_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  or (_02547_, _07936_, _07935_);
  and (_07937_, _05456_, _23996_);
  and (_07938_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_27128_, _07938_, _07937_);
  and (_07939_, _03360_, _23996_);
  and (_07940_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_02554_, _07940_, _07939_);
  and (_07941_, _05456_, _23583_);
  and (_07942_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_27125_, _07942_, _07941_);
  and (_07943_, _05456_, _23548_);
  and (_07945_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_02559_, _07945_, _07943_);
  and (_07946_, _06024_, _05906_);
  not (_07947_, _07946_);
  and (_07948_, _06028_, _06221_);
  not (_07949_, _07948_);
  not (_07950_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_07951_, _06370_, _06034_);
  nor (_07953_, _07951_, _07950_);
  and (_07954_, _07951_, word_in[0]);
  or (_07955_, _07954_, _07953_);
  and (_07956_, _07955_, _07949_);
  and (_07957_, _07948_, word_in[8]);
  or (_07958_, _07957_, _07956_);
  and (_07960_, _07958_, _07947_);
  and (_07962_, _06043_, _06008_);
  and (_07963_, _07962_, _05751_);
  and (_07964_, _07946_, _06538_);
  or (_07966_, _07964_, _07963_);
  or (_07967_, _07966_, _07960_);
  not (_07969_, _07963_);
  or (_07970_, _07969_, _06364_);
  and (_26826_[0], _07970_, _07967_);
  and (_07971_, _05491_, _24051_);
  and (_07973_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  or (_02567_, _07973_, _07971_);
  not (_07974_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_07976_, _07951_, _07974_);
  and (_07977_, _07951_, word_in[1]);
  or (_07978_, _07977_, _07976_);
  or (_07979_, _07978_, _07948_);
  or (_07980_, _07949_, word_in[9]);
  and (_07982_, _07980_, _07979_);
  or (_07984_, _07982_, _07946_);
  or (_07985_, _07947_, _06391_);
  and (_07986_, _07985_, _07984_);
  or (_07987_, _07986_, _07963_);
  or (_07989_, _07969_, _06801_);
  and (_26826_[1], _07989_, _07987_);
  and (_07991_, _07946_, _06572_);
  not (_07992_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_07994_, _07951_, _07992_);
  and (_07996_, _07951_, word_in[2]);
  or (_07998_, _07996_, _07994_);
  and (_07999_, _07998_, _07949_);
  and (_08000_, _07948_, word_in[10]);
  or (_08001_, _08000_, _07999_);
  and (_08003_, _08001_, _07947_);
  or (_08004_, _08003_, _07991_);
  and (_08006_, _08004_, _07969_);
  and (_08007_, _07963_, _06407_);
  or (_26826_[2], _08007_, _08006_);
  not (_08008_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_08009_, _07951_, _08008_);
  and (_08010_, _07951_, word_in[3]);
  or (_08011_, _08010_, _08009_);
  or (_08013_, _08011_, _07948_);
  or (_08014_, _07949_, word_in[11]);
  and (_08015_, _08014_, _08013_);
  and (_08016_, _08015_, _07947_);
  and (_08018_, _07946_, _06586_);
  or (_08019_, _08018_, _07963_);
  or (_08021_, _08019_, _08016_);
  or (_08022_, _07969_, _06441_);
  and (_26826_[3], _08022_, _08021_);
  and (_08024_, _05491_, _24219_);
  and (_08025_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  or (_02575_, _08025_, _08024_);
  not (_08026_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_08027_, _07951_, _08026_);
  and (_08028_, _07951_, word_in[4]);
  or (_08029_, _08028_, _08027_);
  and (_08030_, _08029_, _07949_);
  and (_08031_, _07948_, word_in[12]);
  or (_08032_, _08031_, _08030_);
  and (_08033_, _08032_, _07947_);
  and (_08034_, _07946_, _06591_);
  or (_08035_, _08034_, _07963_);
  or (_08036_, _08035_, _08033_);
  or (_08037_, _07969_, _06446_);
  and (_26826_[4], _08037_, _08036_);
  and (_08038_, _24409_, _24134_);
  and (_08039_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  or (_02579_, _08039_, _08038_);
  not (_08040_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_08041_, _07951_, _08040_);
  and (_08042_, _07951_, word_in[5]);
  or (_08043_, _08042_, _08041_);
  or (_08044_, _08043_, _07948_);
  or (_08045_, _07949_, word_in[13]);
  and (_08046_, _08045_, _08044_);
  and (_08047_, _08046_, _07947_);
  and (_08048_, _07946_, _06606_);
  or (_08049_, _08048_, _07963_);
  or (_08050_, _08049_, _08047_);
  or (_08051_, _07969_, _06463_);
  and (_26826_[5], _08051_, _08050_);
  not (_08052_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_08053_, _07951_, _08052_);
  and (_08054_, _07951_, word_in[6]);
  or (_08055_, _08054_, _08053_);
  or (_08056_, _08055_, _07948_);
  or (_08057_, _07949_, word_in[14]);
  and (_08058_, _08057_, _08056_);
  and (_08059_, _08058_, _07947_);
  and (_08060_, _07946_, _06620_);
  or (_08061_, _08060_, _07963_);
  or (_08062_, _08061_, _08059_);
  or (_08063_, _07969_, _06867_);
  and (_26826_[6], _08063_, _08062_);
  nor (_08064_, _07951_, _05818_);
  and (_08065_, _07951_, word_in[7]);
  or (_08066_, _08065_, _08064_);
  and (_08067_, _08066_, _07949_);
  and (_08068_, _07948_, word_in[15]);
  or (_08069_, _08068_, _08067_);
  and (_08070_, _08069_, _07947_);
  and (_08071_, _07946_, _06047_);
  or (_08072_, _08071_, _07963_);
  or (_08073_, _08072_, _08070_);
  or (_08074_, _07969_, _06052_);
  and (_26826_[7], _08074_, _08073_);
  not (_08075_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_08076_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait , _08075_);
  and (_26885_, _08076_, _22731_);
  and (_08077_, _24409_, _23548_);
  and (_08078_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  or (_27119_, _08078_, _08077_);
  and (_08079_, _05485_, _24089_);
  and (_08080_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_27135_, _08080_, _08079_);
  and (_08081_, _05485_, _24219_);
  and (_08082_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_27133_, _08082_, _08081_);
  and (_08083_, _05431_, _23996_);
  and (_08084_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  or (_27132_, _08084_, _08083_);
  and (_08085_, _05485_, _23887_);
  and (_08086_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_27134_, _08086_, _08085_);
  and (_08088_, _25414_, _24089_);
  and (_08089_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_27160_, _08089_, _08088_);
  and (_08090_, _07779_, _24051_);
  and (_08091_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  or (_27157_, _08091_, _08090_);
  and (_08092_, _02368_, _24134_);
  and (_08093_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  or (_27153_, _08093_, _08092_);
  and (_08094_, _02413_, _23996_);
  and (_08095_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_27150_, _08095_, _08094_);
  and (_08096_, _02455_, _23996_);
  and (_08097_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_27146_, _08097_, _08096_);
  and (_08098_, _06024_, _05753_);
  not (_08099_, _08098_);
  and (_08100_, _06515_, _05800_);
  and (_08101_, _06521_, _06034_);
  and (_08102_, _08101_, word_in[0]);
  not (_08104_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_08105_, _08101_, _08104_);
  nor (_08106_, _08105_, _08102_);
  nor (_08107_, _08106_, _08100_);
  and (_08108_, _08100_, word_in[8]);
  or (_08109_, _08108_, _08107_);
  and (_08110_, _08109_, _08099_);
  and (_08111_, _07962_, _05906_);
  and (_08112_, _08098_, _06538_);
  or (_08113_, _08112_, _08111_);
  or (_08114_, _08113_, _08110_);
  not (_08115_, _08111_);
  or (_08116_, _08115_, _06364_);
  and (_26827_[0], _08116_, _08114_);
  not (_08117_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_08118_, _08101_, _08117_);
  and (_08119_, _08101_, _06548_);
  or (_08120_, _08119_, _08118_);
  or (_08121_, _08120_, _08100_);
  not (_08122_, _08100_);
  or (_08124_, _08122_, word_in[9]);
  and (_08125_, _08124_, _08121_);
  or (_08126_, _08125_, _08098_);
  or (_08127_, _08099_, _06391_);
  and (_08128_, _08127_, _08115_);
  and (_08129_, _08128_, _08126_);
  and (_08130_, _08111_, _06801_);
  or (_26827_[1], _08130_, _08129_);
  and (_08131_, _02517_, _24219_);
  and (_08132_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  or (_27142_, _08132_, _08131_);
  and (_08133_, _08101_, word_in[2]);
  not (_08134_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_08135_, _08101_, _08134_);
  nor (_08136_, _08135_, _08133_);
  nor (_08137_, _08136_, _08100_);
  and (_08138_, _08100_, word_in[10]);
  or (_08139_, _08138_, _08137_);
  and (_08140_, _08139_, _08099_);
  and (_08141_, _08098_, _06572_);
  or (_08143_, _08141_, _08111_);
  or (_08144_, _08143_, _08140_);
  or (_08145_, _08115_, _06407_);
  and (_26827_[2], _08145_, _08144_);
  and (_08146_, _02890_, _24051_);
  and (_08147_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  or (_27141_, _08147_, _08146_);
  not (_08148_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_08149_, _08101_, _08148_);
  and (_08150_, _08101_, _06427_);
  or (_08151_, _08150_, _08149_);
  or (_08152_, _08151_, _08100_);
  or (_08153_, _08122_, word_in[11]);
  and (_08154_, _08153_, _08152_);
  or (_08155_, _08154_, _08098_);
  or (_08156_, _08099_, _06586_);
  and (_08157_, _08156_, _08115_);
  and (_08158_, _08157_, _08155_);
  and (_08159_, _08111_, _06441_);
  or (_26827_[3], _08159_, _08158_);
  and (_08160_, _02890_, _23548_);
  and (_08161_, _02892_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  or (_27140_, _08161_, _08160_);
  not (_08162_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_08163_, _08101_, _08162_);
  and (_08164_, _08101_, _06450_);
  or (_08165_, _08164_, _08163_);
  or (_08166_, _08165_, _08100_);
  or (_08167_, _08122_, word_in[12]);
  and (_08168_, _08167_, _08166_);
  or (_08170_, _08168_, _08098_);
  or (_08171_, _08099_, _06591_);
  and (_08172_, _08171_, _08115_);
  and (_08173_, _08172_, _08170_);
  and (_08174_, _08111_, _06446_);
  or (_26827_[4], _08174_, _08173_);
  and (_08175_, _04812_, _24134_);
  and (_08176_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_27139_, _08176_, _08175_);
  and (_08177_, _08098_, _06606_);
  and (_08178_, _08101_, word_in[5]);
  not (_08179_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_08180_, _08101_, _08179_);
  nor (_08181_, _08180_, _08178_);
  nor (_08182_, _08181_, _08100_);
  and (_08183_, _08100_, word_in[13]);
  or (_08184_, _08183_, _08182_);
  and (_08185_, _08184_, _08099_);
  or (_08186_, _08185_, _08177_);
  and (_08187_, _08186_, _08115_);
  and (_08188_, _08111_, _06463_);
  or (_26827_[5], _08188_, _08187_);
  and (_08189_, _05431_, _24089_);
  and (_08190_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  or (_27130_, _08190_, _08189_);
  and (_08191_, _08101_, word_in[6]);
  not (_08192_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_08193_, _08101_, _08192_);
  nor (_08194_, _08193_, _08191_);
  nor (_08195_, _08194_, _08100_);
  and (_08196_, _08100_, word_in[14]);
  or (_08197_, _08196_, _08195_);
  and (_08198_, _08197_, _08099_);
  and (_08199_, _08098_, _06620_);
  or (_08200_, _08199_, _08111_);
  or (_08201_, _08200_, _08198_);
  or (_08202_, _08115_, _06867_);
  and (_26827_[6], _08202_, _08201_);
  nor (_08203_, _08101_, _05704_);
  and (_08204_, _08101_, _06496_);
  or (_08205_, _08204_, _08203_);
  or (_08206_, _08205_, _08100_);
  or (_08207_, _08122_, word_in[15]);
  and (_08208_, _08207_, _08206_);
  or (_08209_, _08208_, _08098_);
  or (_08210_, _08099_, _06047_);
  and (_08211_, _08210_, _08115_);
  and (_08212_, _08211_, _08209_);
  and (_08213_, _08111_, _06052_);
  or (_26827_[7], _08213_, _08212_);
  and (_08214_, _05456_, _24051_);
  and (_08215_, _05458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_27127_, _08215_, _08214_);
  nand (_08216_, _01816_, _24126_);
  and (_08217_, _02210_, _02320_);
  and (_08218_, _08217_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not (_08219_, _08218_);
  nor (_08220_, _08219_, _01814_);
  not (_08221_, _08220_);
  nor (_08222_, _08221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_08223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_08224_, _08223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_08225_, _08224_, _02210_);
  and (_08226_, _08225_, _02196_);
  nand (_08227_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_08228_, _08227_, _01814_);
  and (_08229_, _08221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_08230_, _08229_, _08228_);
  or (_08231_, _08230_, _08222_);
  or (_08232_, _08231_, _01816_);
  and (_08234_, _08232_, _22731_);
  and (_02667_, _08234_, _08216_);
  and (_08235_, _05491_, _23887_);
  and (_08236_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  or (_27123_, _08236_, _08235_);
  and (_08239_, _24350_, _23887_);
  and (_08241_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_27058_, _08241_, _08239_);
  and (_08243_, _24409_, _23583_);
  and (_08244_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  or (_27120_, _08244_, _08243_);
  and (_08245_, _04812_, _23548_);
  and (_08246_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_27137_, _08246_, _08245_);
  and (_08248_, _05485_, _24134_);
  and (_08250_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_27136_, _08250_, _08248_);
  and (_08251_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_08252_, _04897_, _23887_);
  or (_27008_, _08252_, _08251_);
  and (_08254_, _02455_, _24219_);
  and (_08255_, _02458_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_27144_, _08255_, _08254_);
  and (_08257_, _06024_, _05784_);
  not (_08258_, _08257_);
  and (_08260_, _06653_, _05800_);
  and (_08262_, _06657_, _05962_);
  and (_08263_, _08262_, word_in[0]);
  not (_08264_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor (_08265_, _08262_, _08264_);
  nor (_08267_, _08265_, _08263_);
  nor (_08269_, _08267_, _08260_);
  and (_08271_, _08260_, word_in[8]);
  or (_08273_, _08271_, _08269_);
  and (_08274_, _08273_, _08258_);
  and (_08276_, _06647_, _06008_);
  and (_08277_, _08257_, _06538_);
  or (_08279_, _08277_, _08276_);
  or (_08281_, _08279_, _08274_);
  not (_08282_, _08276_);
  or (_08283_, _08282_, _06364_);
  and (_26828_[0], _08283_, _08281_);
  and (_08285_, _05491_, _24134_);
  and (_08286_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  or (_27124_, _08286_, _08285_);
  not (_08287_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_08289_, _08262_, _08287_);
  and (_08291_, _08262_, word_in[1]);
  nor (_08292_, _08291_, _08289_);
  nor (_08293_, _08292_, _08260_);
  and (_08295_, _08260_, word_in[9]);
  or (_08296_, _08295_, _08293_);
  and (_08297_, _08296_, _08258_);
  and (_08298_, _08257_, _06391_);
  or (_08299_, _08298_, _08276_);
  or (_08300_, _08299_, _08297_);
  or (_08301_, _08282_, _06801_);
  and (_26828_[1], _08301_, _08300_);
  and (_08302_, _24409_, _23996_);
  and (_08303_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  or (_27121_, _08303_, _08302_);
  not (_08304_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_08305_, _08262_, _08304_);
  and (_08306_, _08262_, word_in[2]);
  nor (_08307_, _08306_, _08305_);
  nor (_08308_, _08307_, _08260_);
  and (_08309_, _08260_, word_in[10]);
  or (_08310_, _08309_, _08308_);
  and (_08311_, _08310_, _08258_);
  and (_08312_, _08257_, _06572_);
  or (_08313_, _08312_, _08276_);
  or (_08314_, _08313_, _08311_);
  or (_08315_, _08282_, _06407_);
  and (_26828_[2], _08315_, _08314_);
  not (_08316_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_08317_, _08262_, _08316_);
  and (_08318_, _08262_, word_in[3]);
  nor (_08319_, _08318_, _08317_);
  nor (_08320_, _08319_, _08260_);
  and (_08321_, _08260_, word_in[11]);
  or (_08322_, _08321_, _08320_);
  and (_08323_, _08322_, _08258_);
  and (_08324_, _08257_, _06586_);
  or (_08325_, _08324_, _08276_);
  or (_08326_, _08325_, _08323_);
  or (_08327_, _08282_, _06441_);
  and (_26828_[3], _08327_, _08326_);
  nand (_08328_, _25608_, _23542_);
  and (_08329_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_08330_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_08332_, _08330_, _08329_);
  or (_08333_, _08332_, _25608_);
  and (_08334_, _08333_, _25617_);
  and (_08335_, _08334_, _08328_);
  and (_08336_, _25603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_08337_, _08336_, _08335_);
  and (_02719_, _08337_, _22731_);
  not (_08338_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_08339_, _08262_, _08338_);
  and (_08340_, _08262_, word_in[4]);
  nor (_08341_, _08340_, _08339_);
  nor (_08342_, _08341_, _08260_);
  and (_08343_, _08260_, word_in[12]);
  or (_08344_, _08343_, _08342_);
  and (_08345_, _08344_, _08258_);
  and (_08346_, _08257_, _06591_);
  or (_08347_, _08346_, _08276_);
  or (_08348_, _08347_, _08345_);
  or (_08349_, _08282_, _06446_);
  and (_26828_[4], _08349_, _08348_);
  and (_08350_, _25414_, _24051_);
  and (_08351_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_02721_, _08351_, _08350_);
  not (_08352_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_08353_, _08262_, _08352_);
  and (_08354_, _08262_, word_in[5]);
  nor (_08355_, _08354_, _08353_);
  nor (_08356_, _08355_, _08260_);
  and (_08357_, _08260_, word_in[13]);
  or (_08358_, _08357_, _08356_);
  and (_08359_, _08358_, _08258_);
  and (_08360_, _08257_, _06606_);
  or (_08361_, _08360_, _08276_);
  or (_08362_, _08361_, _08359_);
  or (_08363_, _08282_, _06463_);
  and (_26828_[5], _08363_, _08362_);
  and (_08364_, _02368_, _23996_);
  and (_08365_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  or (_02725_, _08365_, _08364_);
  not (_08366_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_08367_, _08262_, _08366_);
  and (_08368_, _08262_, word_in[6]);
  nor (_08370_, _08368_, _08367_);
  nor (_08371_, _08370_, _08260_);
  and (_08372_, _08260_, word_in[14]);
  or (_08373_, _08372_, _08371_);
  and (_08374_, _08373_, _08258_);
  and (_08375_, _08257_, _06620_);
  or (_08376_, _08375_, _08276_);
  or (_08377_, _08376_, _08374_);
  or (_08379_, _08282_, _06867_);
  and (_26828_[6], _08379_, _08377_);
  nor (_08380_, _08262_, _05811_);
  and (_08382_, _08262_, word_in[7]);
  nor (_08383_, _08382_, _08380_);
  nor (_08384_, _08383_, _08260_);
  and (_08385_, _08260_, word_in[15]);
  or (_08386_, _08385_, _08384_);
  and (_08387_, _08386_, _08258_);
  and (_08388_, _08257_, _06047_);
  or (_08389_, _08388_, _08276_);
  or (_08390_, _08389_, _08387_);
  or (_08391_, _08282_, _06052_);
  and (_26828_[7], _08391_, _08390_);
  and (_08392_, _02517_, _23548_);
  and (_08394_, _02519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  or (_02736_, _08394_, _08392_);
  and (_08395_, _05431_, _24051_);
  and (_08396_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  or (_02741_, _08396_, _08395_);
  and (_08398_, _04812_, _23887_);
  and (_08399_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_02747_, _08399_, _08398_);
  not (_08401_, _25608_);
  nor (_08402_, _08401_, _24126_);
  and (_08403_, _24533_, _24181_);
  and (_08404_, _08403_, _25488_);
  and (_08405_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_08406_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_08407_, _08406_, _08405_);
  nor (_08409_, _08407_, _25608_);
  or (_08411_, _08409_, _08404_);
  or (_08412_, _08411_, _08402_);
  not (_08413_, _08404_);
  or (_08414_, _08413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_08415_, _08414_, _22731_);
  and (_02751_, _08415_, _08412_);
  and (_08416_, _02413_, _24219_);
  and (_08417_, _02415_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_27147_, _08417_, _08416_);
  nand (_08418_, _25603_, _24082_);
  or (_08419_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  not (_08420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nand (_08421_, _25609_, _08420_);
  and (_08422_, _08421_, _08419_);
  or (_08423_, _08422_, _25603_);
  and (_08424_, _08423_, _22731_);
  and (_02763_, _08424_, _08418_);
  or (_08425_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or (_08426_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_08427_, _08426_, _08425_);
  or (_08428_, _08427_, _25603_);
  nand (_08429_, _25603_, _24210_);
  and (_08430_, _08429_, _22731_);
  and (_02766_, _08430_, _08428_);
  and (_08431_, _03013_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  and (_08432_, _03011_, _23548_);
  or (_02770_, _08432_, _08431_);
  and (_08433_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and (_08434_, _06203_, _24134_);
  or (_02773_, _08434_, _08433_);
  and (_08435_, _24159_, _24006_);
  and (_08436_, _08435_, _23583_);
  not (_08437_, _08435_);
  and (_08438_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  or (_02781_, _08438_, _08436_);
  and (_08439_, _25499_, _23577_);
  and (_08440_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_08441_, _08440_, _25523_);
  nand (_08442_, _25509_, _25507_);
  nor (_08443_, _08442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_08444_, _08442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_08445_, _08444_, _25531_);
  or (_08446_, _08445_, _08443_);
  or (_08447_, _08446_, _08441_);
  not (_08448_, _25531_);
  or (_08449_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_08450_, _08449_, _25502_);
  and (_08451_, _08450_, _08447_);
  and (_08452_, _25501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_08453_, _08452_, _08451_);
  or (_08454_, _08453_, _08439_);
  and (_02788_, _08454_, _22731_);
  and (_08455_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_08456_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_08457_, _08456_, _25523_);
  and (_08458_, _25519_, _25507_);
  nor (_08459_, _08458_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_08460_, _08459_, _25543_);
  or (_08461_, _08460_, _25531_);
  or (_08462_, _08461_, _08457_);
  or (_08463_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_08464_, _08463_, _25502_);
  and (_08465_, _08464_, _08462_);
  or (_08466_, _08465_, _08455_);
  and (_08467_, _25556_, _25488_);
  and (_08468_, _08467_, _24179_);
  and (_08469_, _08468_, _02689_);
  or (_08470_, _08469_, _08466_);
  and (_02791_, _08470_, _22731_);
  and (_08471_, _06035_, word_in[0]);
  not (_08472_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_08473_, _06035_, _08472_);
  nor (_08474_, _08473_, _08471_);
  nor (_08475_, _08474_, _06030_);
  and (_08476_, _06030_, word_in[8]);
  or (_08477_, _08476_, _08475_);
  and (_08478_, _08477_, _06027_);
  and (_08479_, _06538_, _06026_);
  or (_08480_, _08479_, _06046_);
  or (_08481_, _08480_, _08478_);
  or (_08482_, _06364_, _06051_);
  and (_26829_[0], _08482_, _08481_);
  and (_08483_, _06035_, word_in[1]);
  not (_08484_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_08485_, _06035_, _08484_);
  nor (_08486_, _08485_, _08483_);
  nor (_08487_, _08486_, _06030_);
  and (_08488_, _06030_, word_in[9]);
  or (_08489_, _08488_, _08487_);
  and (_08491_, _08489_, _06027_);
  and (_08492_, _06391_, _06026_);
  or (_08493_, _08492_, _06046_);
  or (_08494_, _08493_, _08491_);
  or (_08495_, _06801_, _06051_);
  and (_26829_[1], _08495_, _08494_);
  and (_08496_, _06763_, _23996_);
  and (_08497_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_02797_, _08497_, _08496_);
  not (_08498_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_08499_, _06035_, _08498_);
  and (_08500_, _06412_, _06035_);
  or (_08501_, _08500_, _08499_);
  or (_08502_, _08501_, _06030_);
  not (_08503_, _06030_);
  or (_08504_, _08503_, word_in[10]);
  and (_08505_, _08504_, _08502_);
  or (_08506_, _08505_, _06026_);
  or (_08507_, _06572_, _06027_);
  and (_08508_, _08507_, _08506_);
  or (_08509_, _08508_, _06046_);
  or (_08510_, _06407_, _06051_);
  and (_26829_[2], _08510_, _08509_);
  or (_08511_, _08503_, word_in[11]);
  not (_08512_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_08513_, _06035_, _08512_);
  and (_08514_, _06427_, _06035_);
  or (_08515_, _08514_, _08513_);
  or (_08516_, _08515_, _06030_);
  and (_08517_, _08516_, _06027_);
  and (_08518_, _08517_, _08511_);
  and (_08519_, _06586_, _06026_);
  or (_08520_, _08519_, _06046_);
  or (_08521_, _08520_, _08518_);
  or (_08522_, _06441_, _06051_);
  and (_26829_[3], _08522_, _08521_);
  and (_08523_, _24474_, _24006_);
  and (_08524_, _08523_, _23548_);
  not (_08525_, _08523_);
  and (_08526_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  or (_27081_, _08526_, _08524_);
  and (_08527_, _06035_, word_in[4]);
  not (_08528_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_08529_, _06035_, _08528_);
  nor (_08530_, _08529_, _08527_);
  nor (_08531_, _08530_, _06030_);
  and (_08532_, _06030_, word_in[12]);
  or (_08533_, _08532_, _08531_);
  and (_08534_, _08533_, _06027_);
  and (_08535_, _06591_, _06026_);
  or (_08536_, _08535_, _06046_);
  or (_08537_, _08536_, _08534_);
  or (_08538_, _06446_, _06051_);
  and (_26829_[4], _08538_, _08537_);
  and (_08539_, _25479_, _24177_);
  nand (_08540_, _08539_, _23504_);
  not (_08541_, _25489_);
  or (_08542_, _08539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_08543_, _08542_, _08541_);
  and (_08544_, _08543_, _08540_);
  nor (_08545_, _08541_, _23542_);
  or (_08546_, _08545_, _08544_);
  and (_02805_, _08546_, _22731_);
  not (_08547_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_08548_, _06035_, _08547_);
  and (_08549_, _06469_, _06035_);
  or (_08550_, _08549_, _08548_);
  or (_08551_, _08550_, _06030_);
  or (_08552_, _08503_, word_in[13]);
  and (_08553_, _08552_, _08551_);
  or (_08554_, _08553_, _06026_);
  or (_08555_, _06606_, _06027_);
  and (_08556_, _08555_, _08554_);
  or (_08557_, _08556_, _06046_);
  or (_08558_, _06463_, _06051_);
  and (_26829_[5], _08558_, _08557_);
  and (_08559_, _24223_, _24006_);
  and (_08560_, _08559_, _24134_);
  not (_08561_, _08559_);
  and (_08562_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  or (_02808_, _08562_, _08560_);
  or (_08563_, _08503_, word_in[14]);
  not (_08564_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_08565_, _06035_, _08564_);
  and (_08566_, _06623_, _06035_);
  or (_08567_, _08566_, _08565_);
  or (_08568_, _08567_, _06030_);
  and (_08569_, _08568_, _06027_);
  and (_08570_, _08569_, _08563_);
  and (_08571_, _06620_, _06026_);
  or (_08573_, _08571_, _06046_);
  or (_08574_, _08573_, _08570_);
  or (_08575_, _06867_, _06051_);
  and (_26829_[6], _08575_, _08574_);
  and (_08576_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_08577_, _06339_, _24134_);
  or (_02822_, _08577_, _08576_);
  and (_08578_, _24319_, _24006_);
  and (_08579_, _08578_, _23996_);
  not (_08580_, _08578_);
  and (_08581_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  or (_02828_, _08581_, _08579_);
  and (_08582_, _25479_, _24607_);
  nand (_08583_, _08582_, _23504_);
  or (_08584_, _08582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_08585_, _08584_, _08541_);
  and (_08586_, _08585_, _08583_);
  nor (_08587_, _08541_, _24043_);
  or (_08588_, _08587_, _08586_);
  and (_02843_, _08588_, _22731_);
  and (_08589_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_08590_, _06339_, _23996_);
  or (_02850_, _08590_, _08589_);
  and (_08591_, _02039_, _24899_);
  not (_08592_, _08591_);
  and (_08593_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  and (_08594_, _08591_, _23548_);
  or (_02853_, _08594_, _08593_);
  and (_08595_, _24442_, _23548_);
  and (_08596_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  or (_02864_, _08596_, _08595_);
  and (_08598_, _05460_, _23583_);
  and (_08599_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_27073_, _08599_, _08598_);
  and (_08600_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  and (_08601_, _08591_, _23887_);
  or (_02878_, _08601_, _08600_);
  and (_08603_, _05689_, word_in[0]);
  nand (_08604_, _05613_, _07556_);
  or (_08605_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_08607_, _08605_, _08604_);
  and (_08608_, _08607_, _05649_);
  nand (_08609_, _05613_, _08104_);
  or (_08610_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_08611_, _08610_, _08609_);
  and (_08612_, _08611_, _05629_);
  nand (_08613_, _05613_, _07795_);
  or (_08614_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_08615_, _08614_, _08613_);
  and (_08616_, _08615_, _05632_);
  or (_08617_, _08616_, _08612_);
  or (_08618_, _08617_, _08608_);
  nand (_08619_, _05613_, _08472_);
  or (_08620_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_08621_, _08620_, _08619_);
  and (_08622_, _08621_, _05639_);
  or (_08623_, _08622_, _05724_);
  or (_08624_, _08623_, _08618_);
  nand (_08625_, _05613_, _06518_);
  or (_08626_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_08627_, _08626_, _08625_);
  and (_08628_, _08627_, _05649_);
  nand (_08630_, _05613_, _06775_);
  or (_08631_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_08632_, _08631_, _08630_);
  and (_08633_, _08632_, _05632_);
  nand (_08635_, _05613_, _07023_);
  or (_08636_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_08637_, _08636_, _08635_);
  and (_08638_, _08637_, _05629_);
  or (_08639_, _08638_, _08633_);
  or (_08640_, _08639_, _08628_);
  nand (_08641_, _05613_, _07294_);
  or (_08642_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_08643_, _08642_, _08641_);
  and (_08644_, _08643_, _05639_);
  or (_08645_, _08644_, _05617_);
  or (_08646_, _08645_, _08640_);
  and (_08647_, _08646_, _08624_);
  and (_08648_, _08647_, _05688_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _08648_, _08603_);
  and (_08649_, _05689_, word_in[1]);
  nand (_08651_, _05613_, _07573_);
  or (_08652_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_08653_, _08652_, _08651_);
  and (_08654_, _08653_, _05649_);
  nand (_08656_, _05613_, _08117_);
  or (_08657_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_08658_, _08657_, _08656_);
  and (_08659_, _08658_, _05629_);
  nand (_08660_, _05613_, _07816_);
  or (_08661_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_08663_, _08661_, _08660_);
  and (_08664_, _08663_, _05632_);
  or (_08665_, _08664_, _08659_);
  or (_08666_, _08665_, _08654_);
  nand (_08668_, _05613_, _08484_);
  or (_08669_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_08670_, _08669_, _08668_);
  and (_08671_, _08670_, _05639_);
  or (_08672_, _08671_, _05724_);
  or (_08673_, _08672_, _08666_);
  nand (_08674_, _05613_, _06545_);
  or (_08675_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_08676_, _08675_, _08674_);
  and (_08677_, _08676_, _05649_);
  nand (_08678_, _05613_, _06790_);
  or (_08679_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_08680_, _08679_, _08678_);
  and (_08681_, _08680_, _05632_);
  nand (_08682_, _05613_, _07046_);
  or (_08683_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_08684_, _08683_, _08682_);
  and (_08685_, _08684_, _05629_);
  or (_08686_, _08685_, _08681_);
  or (_08687_, _08686_, _08677_);
  nand (_08688_, _05613_, _07310_);
  or (_08689_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_08690_, _08689_, _08688_);
  and (_08691_, _08690_, _05639_);
  or (_08692_, _08691_, _05617_);
  or (_08693_, _08692_, _08687_);
  and (_08695_, _08693_, _08673_);
  and (_08696_, _08695_, _05688_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _08696_, _08649_);
  and (_08697_, _05689_, word_in[2]);
  nand (_08698_, _05613_, _07590_);
  or (_08699_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_08700_, _08699_, _08698_);
  and (_08702_, _08700_, _05649_);
  nand (_08703_, _05613_, _07828_);
  or (_08704_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_08705_, _08704_, _08703_);
  and (_08706_, _08705_, _05632_);
  nand (_08707_, _05613_, _08134_);
  or (_08708_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_08709_, _08708_, _08707_);
  and (_08710_, _08709_, _05629_);
  or (_08712_, _08710_, _08706_);
  or (_08713_, _08712_, _08702_);
  nand (_08714_, _05613_, _08498_);
  or (_08715_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_08716_, _08715_, _08714_);
  and (_08717_, _08716_, _05639_);
  or (_08718_, _08717_, _05724_);
  or (_08719_, _08718_, _08713_);
  nand (_08720_, _05613_, _06562_);
  or (_08721_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_08722_, _08721_, _08720_);
  and (_08723_, _08722_, _05649_);
  nand (_08725_, _05613_, _06804_);
  or (_08726_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_08727_, _08726_, _08725_);
  and (_08729_, _08727_, _05632_);
  nand (_08730_, _05613_, _07063_);
  or (_08731_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_08732_, _08731_, _08730_);
  and (_08733_, _08732_, _05629_);
  or (_08734_, _08733_, _08729_);
  or (_08735_, _08734_, _08723_);
  nand (_08736_, _05613_, _07329_);
  or (_08737_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_08739_, _08737_, _08736_);
  and (_08740_, _08739_, _05639_);
  or (_08741_, _08740_, _05617_);
  or (_08742_, _08741_, _08735_);
  and (_08743_, _08742_, _08719_);
  and (_08744_, _08743_, _05688_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _08744_, _08697_);
  and (_08745_, _05689_, word_in[3]);
  nand (_08747_, _05613_, _07840_);
  or (_08748_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_08749_, _08748_, _08747_);
  and (_08750_, _08749_, _05632_);
  nand (_08751_, _05613_, _08148_);
  or (_08752_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_08753_, _08752_, _08751_);
  and (_08754_, _08753_, _05629_);
  nand (_08755_, _05613_, _07602_);
  or (_08756_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_08757_, _08756_, _08755_);
  and (_08758_, _08757_, _05649_);
  or (_08759_, _08758_, _08754_);
  or (_08760_, _08759_, _08750_);
  nand (_08761_, _05613_, _08512_);
  or (_08762_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_08763_, _08762_, _08761_);
  and (_08764_, _08763_, _05639_);
  or (_08765_, _08764_, _05724_);
  or (_08766_, _08765_, _08760_);
  nand (_08768_, _05613_, _06818_);
  or (_08769_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_08770_, _08769_, _08768_);
  and (_08771_, _08770_, _05632_);
  nand (_08772_, _05613_, _06578_);
  or (_08773_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_08774_, _08773_, _08772_);
  and (_08775_, _08774_, _05649_);
  nand (_08776_, _05613_, _07078_);
  or (_08777_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_08778_, _08777_, _08776_);
  and (_08779_, _08778_, _05629_);
  or (_08781_, _08779_, _08775_);
  or (_08783_, _08781_, _08771_);
  nand (_08784_, _05613_, _07339_);
  or (_08785_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_08786_, _08785_, _08784_);
  and (_08787_, _08786_, _05639_);
  or (_08788_, _08787_, _05617_);
  or (_08789_, _08788_, _08783_);
  and (_08790_, _08789_, _08766_);
  and (_08791_, _08790_, _05688_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _08791_, _08745_);
  and (_08792_, _05689_, word_in[4]);
  nand (_08793_, _05613_, _07854_);
  or (_08794_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_08795_, _08794_, _08793_);
  and (_08796_, _08795_, _05632_);
  nand (_08797_, _05613_, _08162_);
  or (_08798_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_08800_, _08798_, _08797_);
  and (_08801_, _08800_, _05629_);
  nand (_08803_, _05613_, _07616_);
  or (_08804_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_08805_, _08804_, _08803_);
  and (_08806_, _08805_, _05649_);
  or (_08807_, _08806_, _08801_);
  or (_08808_, _08807_, _08796_);
  nand (_08810_, _05613_, _08528_);
  or (_08811_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_08813_, _08811_, _08810_);
  and (_08815_, _08813_, _05639_);
  or (_08816_, _08815_, _05724_);
  or (_08818_, _08816_, _08808_);
  nand (_08819_, _05613_, _06832_);
  or (_08820_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_08821_, _08820_, _08819_);
  and (_08822_, _08821_, _05632_);
  nand (_08823_, _05613_, _06594_);
  or (_08824_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_08826_, _08824_, _08823_);
  and (_08827_, _08826_, _05649_);
  nand (_08828_, _05613_, _07096_);
  or (_08829_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_08830_, _08829_, _08828_);
  and (_08831_, _08830_, _05629_);
  or (_08832_, _08831_, _08827_);
  or (_08833_, _08832_, _08822_);
  nand (_08834_, _05613_, _07357_);
  or (_08835_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_08836_, _08835_, _08834_);
  and (_08837_, _08836_, _05639_);
  or (_08838_, _08837_, _05617_);
  or (_08839_, _08838_, _08833_);
  and (_08840_, _08839_, _08818_);
  and (_08841_, _08840_, _05688_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _08841_, _08792_);
  and (_08842_, _05689_, word_in[5]);
  nand (_08843_, _05613_, _07631_);
  or (_08844_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_08846_, _08844_, _08843_);
  and (_08848_, _08846_, _05649_);
  nand (_08849_, _05613_, _07869_);
  or (_08850_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_08852_, _08850_, _08849_);
  and (_08853_, _08852_, _05632_);
  nand (_08854_, _05613_, _08179_);
  or (_08856_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_08857_, _08856_, _08854_);
  and (_08858_, _08857_, _05629_);
  or (_08859_, _08858_, _08853_);
  or (_08860_, _08859_, _08848_);
  nand (_08861_, _05613_, _08547_);
  or (_08863_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_08864_, _08863_, _08861_);
  and (_08866_, _08864_, _05639_);
  or (_08867_, _08866_, _05724_);
  or (_08868_, _08867_, _08860_);
  nand (_08869_, _05613_, _06609_);
  or (_08870_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_08871_, _08870_, _08869_);
  and (_08872_, _08871_, _05649_);
  nand (_08874_, _05613_, _06845_);
  or (_08875_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_08876_, _08875_, _08874_);
  and (_08877_, _08876_, _05632_);
  nand (_08878_, _05613_, _07112_);
  or (_08879_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_08880_, _08879_, _08878_);
  and (_08881_, _08880_, _05629_);
  or (_08882_, _08881_, _08877_);
  or (_08883_, _08882_, _08872_);
  nand (_08884_, _05613_, _07375_);
  or (_08885_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_08886_, _08885_, _08884_);
  and (_08888_, _08886_, _05639_);
  or (_08889_, _08888_, _05617_);
  or (_08890_, _08889_, _08883_);
  and (_08891_, _08890_, _08868_);
  and (_08893_, _08891_, _05688_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _08893_, _08842_);
  and (_08894_, _05689_, word_in[6]);
  nand (_08895_, _05613_, _07647_);
  or (_08897_, _05613_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_08898_, _08897_, _08895_);
  and (_08899_, _08898_, _05649_);
  nand (_08900_, _05613_, _08192_);
  or (_08901_, _05613_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_08902_, _08901_, _08900_);
  and (_08904_, _08902_, _05629_);
  nand (_08906_, _05613_, _07887_);
  or (_08908_, _05613_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_08909_, _08908_, _08906_);
  and (_08910_, _08909_, _05632_);
  or (_08911_, _08910_, _08904_);
  or (_08913_, _08911_, _08899_);
  nand (_08914_, _05613_, _08564_);
  or (_08915_, _05613_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_08916_, _08915_, _08914_);
  and (_08917_, _08916_, _05639_);
  or (_08918_, _08917_, _05724_);
  or (_08919_, _08918_, _08913_);
  nand (_08920_, _05613_, _06625_);
  or (_08921_, _05613_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_08922_, _08921_, _08920_);
  and (_08924_, _08922_, _05649_);
  nand (_08926_, _05613_, _06857_);
  or (_08927_, _05613_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_08928_, _08927_, _08926_);
  and (_08929_, _08928_, _05632_);
  nand (_08930_, _05613_, _07127_);
  or (_08931_, _05613_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_08933_, _08931_, _08930_);
  and (_08934_, _08933_, _05629_);
  or (_08935_, _08934_, _08929_);
  or (_08936_, _08935_, _08924_);
  nand (_08937_, _05613_, _07384_);
  or (_08938_, _05613_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_08939_, _08938_, _08937_);
  and (_08940_, _08939_, _05639_);
  or (_08941_, _08940_, _05617_);
  or (_08942_, _08941_, _08936_);
  and (_08943_, _08942_, _08919_);
  and (_08944_, _08943_, _05688_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _08944_, _08894_);
  and (_08945_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  and (_08946_, _08591_, _24051_);
  or (_27018_, _08946_, _08945_);
  and (_08948_, _05810_, word_in[8]);
  nand (_08950_, _05613_, _07674_);
  or (_08951_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_08952_, _08951_, _08950_);
  and (_08953_, _08952_, _05787_);
  nand (_08954_, _05613_, _07428_);
  or (_08955_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_08956_, _08955_, _08954_);
  and (_08957_, _08956_, _05785_);
  or (_08958_, _08957_, _08953_);
  and (_08959_, _08958_, _05763_);
  nand (_08960_, _05613_, _06655_);
  or (_08961_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_08962_, _08961_, _08960_);
  and (_08963_, _08962_, _05787_);
  nand (_08964_, _05613_, _06375_);
  or (_08965_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_08966_, _08965_, _08964_);
  and (_08967_, _08966_, _05785_);
  or (_08968_, _08967_, _08963_);
  and (_08969_, _08968_, _05767_);
  nand (_08970_, _05613_, _07170_);
  or (_08972_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_08973_, _08972_, _08970_);
  and (_08974_, _08973_, _05787_);
  nand (_08975_, _05613_, _06892_);
  or (_08976_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_08977_, _08976_, _08975_);
  and (_08978_, _08977_, _05785_);
  or (_08979_, _08978_, _08974_);
  and (_08980_, _08979_, _05797_);
  or (_08981_, _08980_, _08969_);
  nand (_08982_, _05613_, _08264_);
  or (_08983_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_08984_, _08983_, _08982_);
  and (_08985_, _08984_, _05787_);
  nand (_08987_, _05613_, _07950_);
  or (_08988_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_08990_, _08988_, _08987_);
  and (_08991_, _08990_, _05785_);
  or (_08993_, _08991_, _08985_);
  and (_08994_, _08993_, _05800_);
  or (_08996_, _08994_, _08981_);
  nor (_08997_, _08996_, _08959_);
  nor (_08998_, _08997_, _05810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _08998_, _08948_);
  and (_09000_, _05810_, word_in[9]);
  nand (_09001_, _05613_, _07688_);
  or (_09003_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_09005_, _09003_, _09001_);
  and (_09006_, _09005_, _05787_);
  nand (_09007_, _05613_, _07443_);
  or (_09010_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_09011_, _09010_, _09007_);
  and (_09012_, _09011_, _05785_);
  or (_09013_, _09012_, _09006_);
  and (_09015_, _09013_, _05763_);
  nand (_09016_, _05613_, _06674_);
  or (_09018_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_09019_, _09018_, _09016_);
  and (_09020_, _09019_, _05787_);
  nand (_09021_, _05613_, _06393_);
  or (_09022_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_09023_, _09022_, _09021_);
  and (_09024_, _09023_, _05785_);
  or (_09025_, _09024_, _09020_);
  and (_09026_, _09025_, _05767_);
  nand (_09027_, _05613_, _07183_);
  or (_09028_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_09029_, _09028_, _09027_);
  and (_09030_, _09029_, _05787_);
  nand (_09031_, _05613_, _06908_);
  or (_09033_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_09035_, _09033_, _09031_);
  and (_09036_, _09035_, _05785_);
  or (_09037_, _09036_, _09030_);
  and (_09039_, _09037_, _05797_);
  or (_09040_, _09039_, _09026_);
  nand (_09041_, _05613_, _08287_);
  or (_09043_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_09044_, _09043_, _09041_);
  and (_09045_, _09044_, _05787_);
  nand (_09046_, _05613_, _07974_);
  or (_09047_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_09049_, _09047_, _09046_);
  and (_09050_, _09049_, _05785_);
  or (_09051_, _09050_, _09045_);
  and (_09052_, _09051_, _05800_);
  or (_09053_, _09052_, _09040_);
  nor (_09054_, _09053_, _09015_);
  nor (_09055_, _09054_, _05810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _09055_, _09000_);
  and (_09058_, _05810_, word_in[10]);
  nand (_09060_, _05613_, _07700_);
  or (_09062_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_09064_, _09062_, _09060_);
  and (_09065_, _09064_, _05787_);
  nand (_09066_, _05613_, _07458_);
  or (_09067_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_09068_, _09067_, _09066_);
  and (_09070_, _09068_, _05785_);
  or (_09071_, _09070_, _09065_);
  and (_09072_, _09071_, _05763_);
  nand (_09073_, _05613_, _06686_);
  or (_09074_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_09075_, _09074_, _09073_);
  and (_09076_, _09075_, _05787_);
  nand (_09077_, _05613_, _06410_);
  or (_09078_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_09080_, _09078_, _09077_);
  and (_09081_, _09080_, _05785_);
  or (_09082_, _09081_, _09076_);
  and (_09083_, _09082_, _05767_);
  nand (_09084_, _05613_, _07203_);
  or (_09085_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_09086_, _09085_, _09084_);
  and (_09087_, _09086_, _05787_);
  nand (_09088_, _05613_, _06920_);
  or (_09089_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_09090_, _09089_, _09088_);
  and (_09091_, _09090_, _05785_);
  or (_09092_, _09091_, _09087_);
  and (_09094_, _09092_, _05797_);
  or (_09095_, _09094_, _09083_);
  nand (_09097_, _05613_, _08304_);
  or (_09098_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_09099_, _09098_, _09097_);
  and (_09100_, _09099_, _05787_);
  nand (_09101_, _05613_, _07992_);
  or (_09102_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_09104_, _09102_, _09101_);
  and (_09105_, _09104_, _05785_);
  or (_09106_, _09105_, _09100_);
  and (_09107_, _09106_, _05800_);
  or (_09109_, _09107_, _09095_);
  nor (_09110_, _09109_, _09072_);
  nor (_09111_, _09110_, _05810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _09111_, _09058_);
  and (_09114_, _05810_, word_in[11]);
  nand (_09115_, _05613_, _07714_);
  or (_09116_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_09117_, _09116_, _09115_);
  and (_09120_, _09117_, _05787_);
  nand (_09121_, _05613_, _07473_);
  or (_09123_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_09124_, _09123_, _09121_);
  and (_09125_, _09124_, _05785_);
  or (_09126_, _09125_, _09120_);
  and (_09127_, _09126_, _05763_);
  nand (_09128_, _05613_, _06699_);
  or (_09129_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_09131_, _09129_, _09128_);
  and (_09132_, _09131_, _05787_);
  nand (_09134_, _05613_, _06425_);
  or (_09135_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_09137_, _09135_, _09134_);
  and (_09138_, _09137_, _05785_);
  or (_09140_, _09138_, _09132_);
  and (_09142_, _09140_, _05767_);
  nand (_09143_, _05613_, _07218_);
  or (_09144_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_09146_, _09144_, _09143_);
  and (_09149_, _09146_, _05787_);
  nand (_09150_, _05613_, _06934_);
  or (_09151_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_09153_, _09151_, _09150_);
  and (_09154_, _09153_, _05785_);
  or (_09155_, _09154_, _09149_);
  and (_09156_, _09155_, _05797_);
  or (_09158_, _09156_, _09142_);
  nand (_09160_, _05613_, _08316_);
  or (_09161_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_09162_, _09161_, _09160_);
  and (_09163_, _09162_, _05787_);
  nand (_09164_, _05613_, _08008_);
  or (_09165_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_09166_, _09165_, _09164_);
  and (_09167_, _09166_, _05785_);
  or (_09168_, _09167_, _09163_);
  and (_09169_, _09168_, _05800_);
  or (_09170_, _09169_, _09158_);
  nor (_09171_, _09170_, _09127_);
  nor (_09172_, _09171_, _05810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _09172_, _09114_);
  and (_09173_, _05810_, word_in[12]);
  nand (_09174_, _05613_, _07726_);
  or (_09175_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_09176_, _09175_, _09174_);
  and (_09178_, _09176_, _05787_);
  nand (_09179_, _05613_, _07486_);
  or (_09181_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_09182_, _09181_, _09179_);
  and (_09184_, _09182_, _05785_);
  or (_09185_, _09184_, _09178_);
  and (_09186_, _09185_, _05763_);
  nand (_09187_, _05613_, _08338_);
  or (_09189_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_09190_, _09189_, _09187_);
  and (_09192_, _09190_, _05787_);
  nand (_09193_, _05613_, _08026_);
  or (_09194_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_09195_, _09194_, _09193_);
  and (_09197_, _09195_, _05785_);
  or (_09199_, _09197_, _09192_);
  and (_09200_, _09199_, _05800_);
  nand (_09202_, _05613_, _07234_);
  or (_09203_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_09204_, _09203_, _09202_);
  and (_09205_, _09204_, _05787_);
  nand (_09206_, _05613_, _06946_);
  or (_09208_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_09210_, _09208_, _09206_);
  and (_09212_, _09210_, _05785_);
  or (_09213_, _09212_, _09205_);
  and (_09215_, _09213_, _05797_);
  nand (_09217_, _05613_, _06711_);
  or (_09219_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_09221_, _09219_, _09217_);
  and (_09222_, _09221_, _05787_);
  nand (_09223_, _05613_, _06448_);
  or (_09225_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_09227_, _09225_, _09223_);
  and (_09229_, _09227_, _05785_);
  or (_09231_, _09229_, _09222_);
  and (_09233_, _09231_, _05767_);
  or (_09234_, _09233_, _09215_);
  or (_09235_, _09234_, _09200_);
  nor (_09236_, _09235_, _09186_);
  nor (_09237_, _09236_, _05810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _09237_, _09173_);
  and (_09238_, _05810_, word_in[13]);
  nand (_09239_, _05613_, _07738_);
  or (_09240_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_09241_, _09240_, _09239_);
  and (_09242_, _09241_, _05787_);
  nand (_09243_, _05613_, _07498_);
  or (_09244_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_09245_, _09244_, _09243_);
  and (_09246_, _09245_, _05785_);
  or (_09247_, _09246_, _09242_);
  and (_09248_, _09247_, _05763_);
  nand (_09249_, _05613_, _08352_);
  or (_09250_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_09251_, _09250_, _09249_);
  and (_09252_, _09251_, _05787_);
  nand (_09253_, _05613_, _08040_);
  or (_09254_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_09255_, _09254_, _09253_);
  and (_09257_, _09255_, _05785_);
  or (_09258_, _09257_, _09252_);
  and (_09259_, _09258_, _05800_);
  nand (_09260_, _05613_, _07247_);
  or (_09261_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_09262_, _09261_, _09260_);
  and (_09263_, _09262_, _05787_);
  nand (_09264_, _05613_, _06961_);
  or (_09265_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_09266_, _09265_, _09264_);
  and (_09267_, _09266_, _05785_);
  or (_09269_, _09267_, _09263_);
  and (_09271_, _09269_, _05797_);
  nand (_09272_, _05613_, _06726_);
  or (_09273_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_09274_, _09273_, _09272_);
  and (_09275_, _09274_, _05787_);
  nand (_09277_, _05613_, _06466_);
  or (_09278_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_09279_, _09278_, _09277_);
  and (_09280_, _09279_, _05785_);
  or (_09281_, _09280_, _09275_);
  and (_09282_, _09281_, _05767_);
  or (_09283_, _09282_, _09271_);
  or (_09284_, _09283_, _09259_);
  nor (_09285_, _09284_, _09248_);
  nor (_09286_, _09285_, _05810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _09286_, _09238_);
  and (_09288_, _05810_, word_in[14]);
  nand (_09289_, _05613_, _07752_);
  or (_09290_, _05613_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_09291_, _09290_, _09289_);
  and (_09292_, _09291_, _05787_);
  nand (_09293_, _05613_, _07517_);
  or (_09294_, _05613_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_09295_, _09294_, _09293_);
  and (_09296_, _09295_, _05785_);
  or (_09297_, _09296_, _09292_);
  and (_09298_, _09297_, _05763_);
  nand (_09299_, _05613_, _08366_);
  or (_09300_, _05613_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_09301_, _09300_, _09299_);
  and (_09302_, _09301_, _05787_);
  nand (_09303_, _05613_, _08052_);
  or (_09304_, _05613_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_09305_, _09304_, _09303_);
  and (_09306_, _09305_, _05785_);
  or (_09307_, _09306_, _09302_);
  and (_09308_, _09307_, _05800_);
  nand (_09309_, _05613_, _07260_);
  or (_09310_, _05613_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_09311_, _09310_, _09309_);
  and (_09312_, _09311_, _05787_);
  nand (_09313_, _05613_, _06976_);
  or (_09314_, _05613_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_09315_, _09314_, _09313_);
  and (_09316_, _09315_, _05785_);
  or (_09318_, _09316_, _09312_);
  and (_09319_, _09318_, _05797_);
  nand (_09320_, _05613_, _06738_);
  or (_09321_, _05613_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_09322_, _09321_, _09320_);
  and (_09323_, _09322_, _05787_);
  nand (_09324_, _05613_, _06481_);
  or (_09325_, _05613_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_09326_, _09325_, _09324_);
  and (_09327_, _09326_, _05785_);
  or (_09329_, _09327_, _09323_);
  and (_09330_, _09329_, _05767_);
  or (_09332_, _09330_, _09319_);
  or (_09333_, _09332_, _09308_);
  nor (_09334_, _09333_, _09298_);
  nor (_09335_, _09334_, _05810_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _09335_, _09288_);
  and (_09336_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  and (_09337_, _08591_, _23996_);
  or (_02933_, _09337_, _09336_);
  and (_09338_, _05918_, word_in[16]);
  and (_09339_, _08627_, _05639_);
  and (_09340_, _08643_, _05629_);
  or (_09341_, _09340_, _09339_);
  and (_09342_, _08637_, _05632_);
  and (_09343_, _08632_, _05649_);
  or (_09344_, _09343_, _09342_);
  or (_09345_, _09344_, _09341_);
  or (_09346_, _09345_, _05921_);
  and (_09348_, _08611_, _05632_);
  and (_09349_, _08607_, _05639_);
  or (_09350_, _09349_, _09348_);
  and (_09351_, _08621_, _05629_);
  and (_09352_, _08615_, _05649_);
  or (_09353_, _09352_, _09351_);
  nor (_09354_, _09353_, _09350_);
  nand (_09355_, _09354_, _05921_);
  nand (_09356_, _09355_, _09346_);
  nor (_09358_, _09356_, _05918_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _09358_, _09338_);
  and (_09359_, _05918_, word_in[17]);
  and (_09360_, _08684_, _05632_);
  and (_09361_, _08676_, _05639_);
  or (_09362_, _09361_, _09360_);
  and (_09363_, _08690_, _05629_);
  and (_09364_, _08680_, _05649_);
  or (_09365_, _09364_, _09363_);
  or (_09366_, _09365_, _09362_);
  or (_09368_, _09366_, _05921_);
  and (_09369_, _08653_, _05639_);
  and (_09370_, _08670_, _05629_);
  or (_09371_, _09370_, _09369_);
  and (_09372_, _08658_, _05632_);
  and (_09373_, _08663_, _05649_);
  or (_09374_, _09373_, _09372_);
  nor (_09375_, _09374_, _09371_);
  nand (_09376_, _09375_, _05921_);
  nand (_09377_, _09376_, _09368_);
  nor (_09378_, _09377_, _05918_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _09378_, _09359_);
  and (_09379_, _05918_, word_in[18]);
  and (_09380_, _08722_, _05639_);
  and (_09381_, _08739_, _05629_);
  or (_09382_, _09381_, _09380_);
  and (_09383_, _08732_, _05632_);
  and (_09384_, _08727_, _05649_);
  or (_09385_, _09384_, _09383_);
  or (_09386_, _09385_, _09382_);
  or (_09387_, _09386_, _05921_);
  and (_09388_, _08700_, _05639_);
  and (_09389_, _08716_, _05629_);
  or (_09390_, _09389_, _09388_);
  and (_09392_, _08709_, _05632_);
  and (_09393_, _08705_, _05649_);
  or (_09394_, _09393_, _09392_);
  nor (_09395_, _09394_, _09390_);
  nand (_09396_, _09395_, _05921_);
  nand (_09397_, _09396_, _09387_);
  nor (_09398_, _09397_, _05918_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _09398_, _09379_);
  and (_09399_, _05918_, word_in[19]);
  and (_09400_, _08778_, _05632_);
  and (_09401_, _08774_, _05639_);
  or (_09403_, _09401_, _09400_);
  and (_09404_, _08786_, _05629_);
  and (_09405_, _08770_, _05649_);
  or (_09406_, _09405_, _09404_);
  or (_09407_, _09406_, _09403_);
  or (_09408_, _09407_, _05921_);
  and (_09409_, _08757_, _05639_);
  and (_09410_, _08763_, _05629_);
  or (_09411_, _09410_, _09409_);
  and (_09413_, _08753_, _05632_);
  and (_09414_, _08749_, _05649_);
  or (_09415_, _09414_, _09413_);
  nor (_09417_, _09415_, _09411_);
  nand (_09418_, _09417_, _05921_);
  nand (_09419_, _09418_, _09408_);
  nor (_09420_, _09419_, _05918_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _09420_, _09399_);
  and (_09421_, _05918_, word_in[20]);
  and (_09422_, _08826_, _05639_);
  and (_09423_, _08836_, _05629_);
  or (_09424_, _09423_, _09422_);
  and (_09425_, _08830_, _05632_);
  and (_09426_, _08821_, _05649_);
  or (_09428_, _09426_, _09425_);
  or (_09429_, _09428_, _09424_);
  or (_09430_, _09429_, _05921_);
  and (_09431_, _08805_, _05639_);
  and (_09432_, _08813_, _05629_);
  or (_09433_, _09432_, _09431_);
  and (_09434_, _08800_, _05632_);
  and (_09435_, _08795_, _05649_);
  or (_09436_, _09435_, _09434_);
  nor (_09437_, _09436_, _09433_);
  nand (_09438_, _09437_, _05921_);
  nand (_09439_, _09438_, _09430_);
  nor (_09440_, _09439_, _05918_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _09440_, _09421_);
  and (_09441_, _05918_, word_in[21]);
  and (_09442_, _08871_, _05639_);
  and (_09443_, _08886_, _05629_);
  or (_09444_, _09443_, _09442_);
  and (_09445_, _08880_, _05632_);
  and (_09446_, _08876_, _05649_);
  or (_09447_, _09446_, _09445_);
  or (_09449_, _09447_, _09444_);
  or (_09450_, _09449_, _05921_);
  and (_09451_, _08857_, _05632_);
  and (_09452_, _08846_, _05639_);
  or (_09453_, _09452_, _09451_);
  and (_09454_, _08864_, _05629_);
  and (_09455_, _08852_, _05649_);
  or (_09456_, _09455_, _09454_);
  nor (_09457_, _09456_, _09453_);
  nand (_09458_, _09457_, _05921_);
  nand (_09459_, _09458_, _09450_);
  nor (_09460_, _09459_, _05918_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _09460_, _09441_);
  and (_09461_, _05918_, word_in[22]);
  and (_09463_, _08933_, _05632_);
  and (_09464_, _08922_, _05639_);
  or (_09465_, _09464_, _09463_);
  and (_09466_, _08939_, _05629_);
  and (_09467_, _08928_, _05649_);
  or (_09468_, _09467_, _09466_);
  or (_09469_, _09468_, _09465_);
  or (_09470_, _09469_, _05921_);
  and (_09471_, _08902_, _05632_);
  and (_09472_, _08898_, _05639_);
  or (_09473_, _09472_, _09471_);
  and (_09474_, _08916_, _05629_);
  and (_09475_, _08909_, _05649_);
  or (_09476_, _09475_, _09474_);
  nor (_09477_, _09476_, _09473_);
  nand (_09478_, _09477_, _05921_);
  nand (_09480_, _09478_, _09470_);
  nor (_09481_, _09480_, _05918_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _09481_, _09461_);
  and (_09482_, _05991_, word_in[24]);
  and (_09483_, _08956_, _05787_);
  and (_09484_, _08952_, _05785_);
  or (_09485_, _09484_, _09483_);
  and (_09486_, _09485_, _05957_);
  and (_09487_, _08966_, _05787_);
  and (_09488_, _08962_, _05785_);
  or (_09489_, _09488_, _09487_);
  and (_09490_, _09489_, _05996_);
  and (_09491_, _08977_, _05787_);
  and (_09492_, _08973_, _05785_);
  or (_09493_, _09492_, _09491_);
  and (_09494_, _09493_, _06003_);
  and (_09495_, _08990_, _05787_);
  and (_09496_, _08984_, _05785_);
  or (_09497_, _09496_, _09495_);
  and (_09498_, _09497_, _06008_);
  or (_09500_, _09498_, _09494_);
  or (_09501_, _09500_, _09490_);
  nor (_09502_, _09501_, _09486_);
  nor (_09503_, _09502_, _05991_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _09503_, _09482_);
  and (_09504_, _05991_, word_in[25]);
  and (_09505_, _09011_, _05787_);
  and (_09506_, _09005_, _05785_);
  or (_09507_, _09506_, _09505_);
  and (_09508_, _09507_, _05957_);
  and (_09509_, _09023_, _05787_);
  and (_09510_, _09019_, _05785_);
  or (_09511_, _09510_, _09509_);
  and (_09512_, _09511_, _05996_);
  and (_09514_, _09035_, _05787_);
  and (_09515_, _09029_, _05785_);
  or (_09516_, _09515_, _09514_);
  and (_09517_, _09516_, _06003_);
  and (_09518_, _09049_, _05787_);
  and (_09519_, _09044_, _05785_);
  or (_09520_, _09519_, _09518_);
  and (_09521_, _09520_, _06008_);
  or (_09522_, _09521_, _09517_);
  or (_09523_, _09522_, _09512_);
  nor (_09524_, _09523_, _09508_);
  nor (_09525_, _09524_, _05991_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _09525_, _09504_);
  and (_09526_, _05991_, word_in[26]);
  and (_09527_, _09068_, _05787_);
  and (_09528_, _09064_, _05785_);
  or (_09529_, _09528_, _09527_);
  and (_09530_, _09529_, _05957_);
  and (_09531_, _09080_, _05787_);
  and (_09532_, _09075_, _05785_);
  or (_09533_, _09532_, _09531_);
  and (_09534_, _09533_, _05996_);
  and (_09535_, _09090_, _05787_);
  and (_09536_, _09086_, _05785_);
  or (_09537_, _09536_, _09535_);
  and (_09538_, _09537_, _06003_);
  and (_09540_, _09104_, _05787_);
  and (_09541_, _09099_, _05785_);
  or (_09542_, _09541_, _09540_);
  and (_09543_, _09542_, _06008_);
  or (_09545_, _09543_, _09538_);
  or (_09546_, _09545_, _09534_);
  nor (_09547_, _09546_, _09530_);
  nor (_09548_, _09547_, _05991_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _09548_, _09526_);
  and (_09549_, _05991_, word_in[27]);
  and (_09550_, _09137_, _05787_);
  and (_09551_, _09131_, _05785_);
  or (_09552_, _09551_, _09550_);
  and (_09553_, _09552_, _05996_);
  and (_09554_, _09124_, _05787_);
  and (_09555_, _09117_, _05785_);
  or (_09556_, _09555_, _09554_);
  and (_09557_, _09556_, _05957_);
  and (_09558_, _09153_, _05787_);
  and (_09559_, _09146_, _05785_);
  or (_09561_, _09559_, _09558_);
  and (_09562_, _09561_, _06003_);
  and (_09563_, _09166_, _05787_);
  and (_09564_, _09162_, _05785_);
  or (_09565_, _09564_, _09563_);
  and (_09566_, _09565_, _06008_);
  or (_09567_, _09566_, _09562_);
  or (_09568_, _09567_, _09557_);
  nor (_09569_, _09568_, _09553_);
  nor (_09570_, _09569_, _05991_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _09570_, _09549_);
  and (_09571_, _05991_, word_in[28]);
  and (_09572_, _09227_, _05787_);
  and (_09573_, _09221_, _05785_);
  or (_09574_, _09573_, _09572_);
  and (_09575_, _09574_, _05996_);
  and (_09576_, _09182_, _05787_);
  and (_09577_, _09176_, _05785_);
  or (_09578_, _09577_, _09576_);
  and (_09579_, _09578_, _05957_);
  and (_09581_, _09210_, _05787_);
  and (_09582_, _09204_, _05785_);
  or (_09583_, _09582_, _09581_);
  and (_09584_, _09583_, _06003_);
  and (_09585_, _09195_, _05787_);
  and (_09586_, _09190_, _05785_);
  or (_09587_, _09586_, _09585_);
  and (_09588_, _09587_, _06008_);
  or (_09589_, _09588_, _09584_);
  or (_09590_, _09589_, _09579_);
  nor (_09591_, _09590_, _09575_);
  nor (_09592_, _09591_, _05991_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _09592_, _09571_);
  and (_09593_, _05991_, word_in[29]);
  and (_09594_, _09245_, _05787_);
  and (_09595_, _09241_, _05785_);
  or (_09596_, _09595_, _09594_);
  and (_09597_, _09596_, _05957_);
  and (_09598_, _09279_, _05787_);
  and (_09599_, _09274_, _05785_);
  or (_09601_, _09599_, _09598_);
  and (_09602_, _09601_, _05996_);
  and (_09603_, _09266_, _05787_);
  and (_09604_, _09262_, _05785_);
  or (_09605_, _09604_, _09603_);
  and (_09606_, _09605_, _06003_);
  and (_09607_, _09255_, _05787_);
  and (_09608_, _09251_, _05785_);
  or (_09609_, _09608_, _09607_);
  and (_09610_, _09609_, _06008_);
  or (_09611_, _09610_, _09606_);
  or (_09612_, _09611_, _09602_);
  nor (_09614_, _09612_, _09597_);
  nor (_09615_, _09614_, _05991_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _09615_, _09593_);
  and (_09616_, _05991_, word_in[30]);
  and (_09617_, _09295_, _05787_);
  and (_09618_, _09291_, _05785_);
  or (_09619_, _09618_, _09617_);
  and (_09620_, _09619_, _05957_);
  and (_09622_, _09326_, _05787_);
  and (_09623_, _09322_, _05785_);
  or (_09624_, _09623_, _09622_);
  and (_09625_, _09624_, _05996_);
  and (_09626_, _09315_, _05787_);
  and (_09627_, _09311_, _05785_);
  or (_09628_, _09627_, _09626_);
  and (_09629_, _09628_, _06003_);
  and (_09631_, _09305_, _05787_);
  and (_09632_, _09301_, _05785_);
  or (_09633_, _09632_, _09631_);
  and (_09634_, _09633_, _06008_);
  or (_09635_, _09634_, _09629_);
  or (_09636_, _09635_, _09625_);
  nor (_09637_, _09636_, _09620_);
  nor (_09638_, _09637_, _05991_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _09638_, _09616_);
  and (_09639_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_09640_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_09641_, _22740_, _09640_);
  or (_09642_, _09641_, _09639_);
  and (_26862_[1], _09642_, _22731_);
  and (_09643_, _24350_, _24134_);
  and (_09644_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_27062_, _09644_, _09643_);
  and (_09645_, _02039_, _23941_);
  not (_09646_, _09645_);
  and (_09647_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  and (_09648_, _09645_, _24219_);
  or (_03000_, _09648_, _09647_);
  and (_09651_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  and (_09652_, _09645_, _23887_);
  or (_03012_, _09652_, _09651_);
  and (_09653_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  and (_09654_, _09645_, _24089_);
  or (_03027_, _09654_, _09653_);
  and (_09655_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  and (_09656_, _09645_, _24134_);
  or (_03047_, _09656_, _09655_);
  and (_09657_, _24415_, _24089_);
  and (_09658_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  or (_03051_, _09658_, _09657_);
  and (_09659_, _24485_, _24134_);
  and (_09660_, _24487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  or (_03053_, _09660_, _09659_);
  and (_09661_, _25206_, _23583_);
  and (_09663_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_03056_, _09663_, _09661_);
  and (_09665_, _25442_, _23996_);
  and (_09667_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_27035_, _09667_, _09665_);
  and (_09668_, _25648_, _24134_);
  and (_09669_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  or (_27032_, _09669_, _09668_);
  and (_09670_, _24365_, _24236_);
  and (_09671_, _09670_, _23996_);
  not (_09672_, _09670_);
  and (_09673_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  or (_03063_, _09673_, _09671_);
  and (_09674_, _25648_, _23887_);
  and (_09675_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  or (_03064_, _09675_, _09674_);
  and (_09676_, _02039_, _24349_);
  not (_09677_, _09676_);
  and (_09678_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_09679_, _09676_, _23548_);
  or (_03069_, _09679_, _09678_);
  and (_09680_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_09681_, _09676_, _24089_);
  or (_03076_, _09681_, _09680_);
  and (_09682_, _24442_, _24134_);
  and (_09683_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  or (_03079_, _09683_, _09682_);
  and (_09684_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  and (_09685_, _02338_, _24219_);
  or (_03092_, _09685_, _09684_);
  and (_09687_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  and (_09689_, _02836_, _24051_);
  or (_03095_, _09689_, _09687_);
  and (_09690_, _02990_, _23583_);
  and (_09692_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  or (_03099_, _09692_, _09690_);
  and (_09693_, _02990_, _24219_);
  and (_09694_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  or (_27053_, _09694_, _09693_);
  and (_09695_, _03186_, _24089_);
  and (_09696_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  or (_03103_, _09696_, _09695_);
  and (_09697_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_09698_, _09676_, _24051_);
  or (_27022_, _09698_, _09697_);
  and (_09699_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_09700_, _09676_, _23996_);
  or (_03112_, _09700_, _09699_);
  and (_09701_, _02065_, _23583_);
  and (_09702_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  or (_03116_, _09702_, _09701_);
  and (_09703_, _24051_, _24008_);
  and (_09704_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or (_03117_, _09704_, _09703_);
  and (_09705_, _02039_, _24236_);
  not (_09706_, _09705_);
  and (_09707_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_09708_, _09705_, _24219_);
  or (_03123_, _09708_, _09707_);
  and (_09709_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_09710_, _09705_, _23583_);
  or (_03125_, _09710_, _09709_);
  and (_09711_, _24889_, _24051_);
  and (_09712_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_03130_, _09712_, _09711_);
  and (_09713_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_09714_, _09705_, _24089_);
  or (_03154_, _09714_, _09713_);
  and (_09715_, _04920_, _23583_);
  and (_09716_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_03156_, _09716_, _09715_);
  and (_09717_, _24159_, _23945_);
  and (_09718_, _09717_, _24089_);
  not (_09719_, _09717_);
  and (_09720_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_03160_, _09720_, _09718_);
  and (_09722_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_09723_, _09705_, _24134_);
  or (_03163_, _09723_, _09722_);
  and (_09724_, _24237_, _23583_);
  and (_09725_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_27063_, _09725_, _09724_);
  and (_09726_, _24330_, _24134_);
  and (_09727_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_03177_, _09727_, _09726_);
  and (_09728_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_09729_, _09705_, _23996_);
  or (_03179_, _09729_, _09728_);
  and (_09730_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_09731_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_09732_, _22740_, _09731_);
  or (_09733_, _09732_, _09730_);
  and (_26862_[0], _09733_, _22731_);
  and (_09734_, _02478_, _24219_);
  and (_09736_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or (_03196_, _09736_, _09734_);
  and (_09737_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  and (_09738_, _04853_, _24134_);
  or (_03206_, _09738_, _09737_);
  and (_09739_, _25442_, _23887_);
  and (_09740_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_03216_, _09740_, _09739_);
  and (_09742_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  and (_09744_, _04853_, _24051_);
  or (_03223_, _09744_, _09742_);
  and (_09746_, _02990_, _23996_);
  and (_09747_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  or (_03240_, _09747_, _09746_);
  and (_09749_, _23890_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_09750_, _23845_, _26578_);
  and (_09751_, _23909_, _23800_);
  or (_09752_, _03899_, _09751_);
  or (_09753_, _09752_, _09750_);
  not (_09754_, _26736_);
  or (_09756_, _24253_, _23913_);
  or (_09757_, _09756_, _09754_);
  or (_09758_, _09757_, _09753_);
  or (_09759_, _23916_, _23839_);
  or (_09760_, _26739_, _23901_);
  or (_09761_, _09760_, _09759_);
  and (_09762_, _23841_, _23708_);
  and (_09763_, _24247_, _23896_);
  or (_09764_, _09763_, _24248_);
  or (_09765_, _09764_, _09762_);
  or (_09767_, _09765_, _23906_);
  or (_09769_, _09767_, _09761_);
  or (_09771_, _09769_, _23934_);
  or (_09772_, _09771_, _09758_);
  and (_09773_, _09772_, _23855_);
  or (_26850_[0], _09773_, _09749_);
  and (_09774_, _24496_, _24319_);
  and (_09775_, _09774_, _24051_);
  not (_09777_, _09774_);
  and (_09778_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  or (_03262_, _09778_, _09775_);
  and (_09779_, _23944_, _22977_);
  and (_09780_, _09779_, _24159_);
  and (_09781_, _09780_, _23996_);
  not (_09782_, _09780_);
  and (_09783_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or (_27006_, _09783_, _09781_);
  and (_09784_, _07013_, _24219_);
  and (_09785_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or (_03268_, _09785_, _09784_);
  and (_09787_, _09780_, _24134_);
  and (_09789_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or (_27005_, _09789_, _09787_);
  not (_09790_, _05520_);
  not (_09791_, _05535_);
  and (_09792_, _05548_, _05547_);
  and (_09793_, _05513_, _05511_);
  and (_09794_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  and (_09795_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  or (_09796_, _09795_, _09794_);
  and (_09797_, _09796_, _09792_);
  and (_09798_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  and (_09799_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  or (_09801_, _09799_, _09798_);
  and (_09802_, _09801_, _05549_);
  or (_09803_, _09802_, _09797_);
  or (_09804_, _09803_, _09791_);
  not (_09805_, _05542_);
  and (_09806_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  and (_09808_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_09811_, _09808_, _09806_);
  and (_09812_, _09811_, _09792_);
  and (_09813_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  and (_09814_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_09815_, _09814_, _09813_);
  and (_09816_, _09815_, _05549_);
  or (_09817_, _09816_, _09812_);
  or (_09818_, _09817_, _05535_);
  and (_09819_, _09818_, _09805_);
  and (_09820_, _09819_, _09804_);
  or (_09821_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_09822_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  and (_09823_, _09822_, _09821_);
  and (_09824_, _09823_, _09792_);
  or (_09825_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_09827_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  and (_09828_, _09827_, _09825_);
  and (_09829_, _09828_, _05549_);
  or (_09830_, _09829_, _09824_);
  or (_09831_, _09830_, _09791_);
  or (_09832_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  or (_09833_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  and (_09834_, _09833_, _09832_);
  and (_09836_, _09834_, _09792_);
  or (_09838_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_09839_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  and (_09840_, _09839_, _09838_);
  and (_09841_, _09840_, _05549_);
  or (_09842_, _09841_, _09836_);
  or (_09843_, _09842_, _05535_);
  and (_09845_, _09843_, _05542_);
  and (_09847_, _09845_, _09831_);
  or (_09848_, _09847_, _09820_);
  and (_09849_, _09848_, _05518_);
  not (_09850_, _05518_);
  and (_09851_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  and (_09852_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_09853_, _09852_, _09851_);
  and (_09855_, _09853_, _09792_);
  and (_09856_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  and (_09857_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  or (_09858_, _09857_, _09856_);
  and (_09859_, _09858_, _05549_);
  or (_09860_, _09859_, _09855_);
  or (_09861_, _09860_, _09791_);
  and (_09862_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  and (_09863_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  or (_09865_, _09863_, _09862_);
  and (_09866_, _09865_, _09792_);
  and (_09867_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  and (_09869_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  or (_09870_, _09869_, _09867_);
  and (_09871_, _09870_, _05549_);
  or (_09872_, _09871_, _09866_);
  or (_09873_, _09872_, _05535_);
  and (_09874_, _09873_, _09805_);
  and (_09876_, _09874_, _09861_);
  or (_09877_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  or (_09878_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  and (_09879_, _09878_, _05549_);
  and (_09880_, _09879_, _09877_);
  or (_09882_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  or (_09883_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  and (_09885_, _09883_, _09792_);
  and (_09887_, _09885_, _09882_);
  or (_09888_, _09887_, _09880_);
  or (_09889_, _09888_, _09791_);
  or (_09890_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_09892_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  and (_09893_, _09892_, _05549_);
  and (_09895_, _09893_, _09890_);
  or (_09897_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_09898_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  and (_09899_, _09898_, _09792_);
  and (_09900_, _09899_, _09897_);
  or (_09901_, _09900_, _09895_);
  or (_09902_, _09901_, _05535_);
  and (_09903_, _09902_, _05542_);
  and (_09904_, _09903_, _09889_);
  or (_09905_, _09904_, _09876_);
  and (_09906_, _09905_, _09850_);
  or (_09907_, _09906_, _09849_);
  and (_09909_, _09907_, _09790_);
  and (_09910_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_09912_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_09913_, _09912_, _09910_);
  and (_09915_, _09913_, _09792_);
  and (_09917_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_09919_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_09921_, _09919_, _09917_);
  and (_09923_, _09921_, _05549_);
  or (_09924_, _09923_, _09915_);
  and (_09925_, _09924_, _05535_);
  and (_09926_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_09927_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_09928_, _09927_, _09926_);
  and (_09930_, _09928_, _09792_);
  and (_09931_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_09932_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_09933_, _09932_, _09931_);
  and (_09934_, _09933_, _05549_);
  or (_09935_, _09934_, _09930_);
  and (_09936_, _09935_, _09791_);
  or (_09937_, _09936_, _09925_);
  and (_09938_, _09937_, _09805_);
  or (_09940_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_09941_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_09942_, _09941_, _05549_);
  and (_09943_, _09942_, _09940_);
  or (_09944_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_09945_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_09946_, _09945_, _09792_);
  and (_09947_, _09946_, _09944_);
  or (_09948_, _09947_, _09943_);
  and (_09949_, _09948_, _05535_);
  or (_09951_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_09952_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_09954_, _09952_, _05549_);
  and (_09956_, _09954_, _09951_);
  or (_09957_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_09958_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_09960_, _09958_, _09792_);
  and (_09962_, _09960_, _09957_);
  or (_09963_, _09962_, _09956_);
  and (_09964_, _09963_, _09791_);
  or (_09965_, _09964_, _09949_);
  and (_09967_, _09965_, _05542_);
  or (_09968_, _09967_, _09938_);
  and (_09969_, _09968_, _09850_);
  and (_09971_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  and (_09973_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_09975_, _09973_, _09971_);
  and (_09976_, _09975_, _09792_);
  and (_09978_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  and (_09979_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  or (_09981_, _09979_, _09978_);
  and (_09982_, _09981_, _05549_);
  or (_09983_, _09982_, _09976_);
  and (_09984_, _09983_, _05535_);
  and (_09985_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  and (_09987_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  or (_09988_, _09987_, _09985_);
  and (_09989_, _09988_, _09792_);
  and (_09990_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  and (_09991_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  or (_09992_, _09991_, _09990_);
  and (_09993_, _09992_, _05549_);
  or (_09994_, _09993_, _09989_);
  and (_09995_, _09994_, _09791_);
  or (_09997_, _09995_, _09984_);
  and (_09998_, _09997_, _09805_);
  or (_09999_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_10000_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  and (_10002_, _10000_, _09999_);
  and (_10004_, _10002_, _09792_);
  or (_10005_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_10007_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  and (_10009_, _10007_, _10005_);
  and (_10010_, _10009_, _05549_);
  or (_10011_, _10010_, _10004_);
  and (_10013_, _10011_, _05535_);
  or (_10014_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_10015_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  and (_10016_, _10015_, _10014_);
  and (_10017_, _10016_, _09792_);
  or (_10019_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_10020_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  and (_10021_, _10020_, _10019_);
  and (_10022_, _10021_, _05549_);
  or (_10023_, _10022_, _10017_);
  and (_10024_, _10023_, _09791_);
  or (_10025_, _10024_, _10013_);
  and (_10026_, _10025_, _05542_);
  or (_10027_, _10026_, _09998_);
  and (_10028_, _10027_, _05518_);
  or (_10029_, _10028_, _09969_);
  and (_10030_, _10029_, _05520_);
  or (_10031_, _10030_, _09909_);
  or (_10032_, _10031_, _05526_);
  not (_10033_, _05526_);
  and (_10034_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  and (_10035_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_10036_, _10035_, _10034_);
  and (_10037_, _10036_, _09792_);
  and (_10038_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  and (_10039_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  or (_10041_, _10039_, _10038_);
  and (_10042_, _10041_, _05549_);
  or (_10044_, _10042_, _10037_);
  or (_10046_, _10044_, _09791_);
  and (_10047_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  and (_10049_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_10051_, _10049_, _10047_);
  and (_10052_, _10051_, _09792_);
  and (_10053_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  and (_10054_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_10056_, _10054_, _10053_);
  and (_10057_, _10056_, _05549_);
  or (_10058_, _10057_, _10052_);
  or (_10060_, _10058_, _05535_);
  and (_10062_, _10060_, _09805_);
  and (_10063_, _10062_, _10046_);
  or (_10064_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_10065_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  and (_10066_, _10065_, _05549_);
  and (_10067_, _10066_, _10064_);
  or (_10068_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_10069_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  and (_10071_, _10069_, _09792_);
  and (_10072_, _10071_, _10068_);
  or (_10073_, _10072_, _10067_);
  or (_10074_, _10073_, _09791_);
  or (_10075_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_10076_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  and (_10077_, _10076_, _05549_);
  and (_10078_, _10077_, _10075_);
  or (_10079_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_10080_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  and (_10081_, _10080_, _09792_);
  and (_10082_, _10081_, _10079_);
  or (_10083_, _10082_, _10078_);
  or (_10084_, _10083_, _05535_);
  and (_10085_, _10084_, _05542_);
  and (_10086_, _10085_, _10074_);
  or (_10087_, _10086_, _10063_);
  and (_10088_, _10087_, _09850_);
  and (_10089_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  and (_10091_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_10092_, _10091_, _10089_);
  and (_10094_, _10092_, _09792_);
  and (_10095_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  and (_10096_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_10098_, _10096_, _10095_);
  and (_10099_, _10098_, _05549_);
  or (_10100_, _10099_, _10094_);
  or (_10101_, _10100_, _09791_);
  and (_10103_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  and (_10104_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_10105_, _10104_, _10103_);
  and (_10106_, _10105_, _09792_);
  and (_10108_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  and (_10109_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_10110_, _10109_, _10108_);
  and (_10112_, _10110_, _05549_);
  or (_10114_, _10112_, _10106_);
  or (_10116_, _10114_, _05535_);
  and (_10117_, _10116_, _09805_);
  and (_10119_, _10117_, _10101_);
  or (_10121_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_10122_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  and (_10123_, _10122_, _10121_);
  and (_10124_, _10123_, _09792_);
  or (_10125_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_10127_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  and (_10128_, _10127_, _10125_);
  and (_10129_, _10128_, _05549_);
  or (_10131_, _10129_, _10124_);
  or (_10133_, _10131_, _09791_);
  or (_10134_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_10135_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  and (_10137_, _10135_, _10134_);
  and (_10138_, _10137_, _09792_);
  or (_10139_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_10141_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  and (_10142_, _10141_, _10139_);
  and (_10143_, _10142_, _05549_);
  or (_10145_, _10143_, _10138_);
  or (_10146_, _10145_, _05535_);
  and (_10148_, _10146_, _05542_);
  and (_10149_, _10148_, _10133_);
  or (_10150_, _10149_, _10119_);
  and (_10152_, _10150_, _05518_);
  or (_10153_, _10152_, _10088_);
  and (_10155_, _10153_, _09790_);
  or (_10156_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_10157_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  and (_10158_, _10157_, _10156_);
  and (_10159_, _10158_, _09792_);
  or (_10160_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_10162_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  and (_10163_, _10162_, _10160_);
  and (_10164_, _10163_, _05549_);
  or (_10165_, _10164_, _10159_);
  and (_10167_, _10165_, _09791_);
  or (_10168_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_10169_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  and (_10171_, _10169_, _10168_);
  and (_10172_, _10171_, _09792_);
  or (_10174_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_10176_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  and (_10178_, _10176_, _10174_);
  and (_10180_, _10178_, _05549_);
  or (_10182_, _10180_, _10172_);
  and (_10183_, _10182_, _05535_);
  or (_10184_, _10183_, _10167_);
  and (_10185_, _10184_, _05542_);
  and (_10187_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  and (_10188_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  or (_10189_, _10188_, _10187_);
  and (_10191_, _10189_, _09792_);
  and (_10192_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  and (_10193_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  or (_10195_, _10193_, _10192_);
  and (_10197_, _10195_, _05549_);
  or (_10199_, _10197_, _10191_);
  and (_10200_, _10199_, _09791_);
  and (_10202_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  and (_10203_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  or (_10204_, _10203_, _10202_);
  and (_10205_, _10204_, _09792_);
  and (_10206_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  and (_10207_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_10208_, _10207_, _10206_);
  and (_10209_, _10208_, _05549_);
  or (_10210_, _10209_, _10205_);
  and (_10211_, _10210_, _05535_);
  or (_10212_, _10211_, _10200_);
  and (_10213_, _10212_, _09805_);
  or (_10215_, _10213_, _10185_);
  and (_10216_, _10215_, _05518_);
  or (_10217_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_10218_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  and (_10219_, _10218_, _05549_);
  and (_10221_, _10219_, _10217_);
  or (_10222_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or (_10223_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  and (_10224_, _10223_, _09792_);
  and (_10225_, _10224_, _10222_);
  or (_10226_, _10225_, _10221_);
  and (_10227_, _10226_, _09791_);
  or (_10228_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  or (_10229_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  and (_10230_, _10229_, _05549_);
  and (_10231_, _10230_, _10228_);
  or (_10232_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  or (_10233_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  and (_10234_, _10233_, _09792_);
  and (_10235_, _10234_, _10232_);
  or (_10236_, _10235_, _10231_);
  and (_10237_, _10236_, _05535_);
  or (_10238_, _10237_, _10227_);
  and (_10239_, _10238_, _05542_);
  and (_10240_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  and (_10241_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_10243_, _10241_, _10240_);
  and (_10245_, _10243_, _09792_);
  and (_10246_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  and (_10247_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  or (_10248_, _10247_, _10246_);
  and (_10249_, _10248_, _05549_);
  or (_10251_, _10249_, _10245_);
  and (_10252_, _10251_, _09791_);
  and (_10253_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  and (_10254_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_10255_, _10254_, _10253_);
  and (_10256_, _10255_, _09792_);
  and (_10257_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  and (_10258_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or (_10259_, _10258_, _10257_);
  and (_10261_, _10259_, _05549_);
  or (_10262_, _10261_, _10256_);
  and (_10263_, _10262_, _05535_);
  or (_10264_, _10263_, _10252_);
  and (_10265_, _10264_, _09805_);
  or (_10267_, _10265_, _10239_);
  and (_10268_, _10267_, _09850_);
  or (_10269_, _10268_, _10216_);
  and (_10270_, _10269_, _05520_);
  or (_10271_, _10270_, _10155_);
  or (_10272_, _10271_, _10033_);
  and (_10273_, _10272_, _10032_);
  or (_10274_, _10273_, _00143_);
  and (_10275_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_10276_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  or (_10277_, _10276_, _10275_);
  and (_10278_, _10277_, _05549_);
  and (_10279_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  and (_10280_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  or (_10281_, _10280_, _10279_);
  and (_10282_, _10281_, _09792_);
  or (_10283_, _10282_, _10278_);
  or (_10284_, _10283_, _09791_);
  and (_10285_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  and (_10286_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  or (_10287_, _10286_, _10285_);
  and (_10288_, _10287_, _05549_);
  and (_10289_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_10290_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  or (_10291_, _10290_, _10289_);
  and (_10292_, _10291_, _09792_);
  or (_10294_, _10292_, _10288_);
  or (_10295_, _10294_, _05535_);
  and (_10296_, _10295_, _09805_);
  and (_10297_, _10296_, _10284_);
  or (_10298_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  or (_10299_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  and (_10300_, _10299_, _09792_);
  and (_10301_, _10300_, _10298_);
  or (_10302_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  or (_10303_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_10305_, _10303_, _05549_);
  and (_10306_, _10305_, _10302_);
  or (_10307_, _10306_, _10301_);
  or (_10308_, _10307_, _09791_);
  or (_10309_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  or (_10310_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  and (_10311_, _10310_, _09792_);
  and (_10312_, _10311_, _10309_);
  or (_10313_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  or (_10314_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_10315_, _10314_, _05549_);
  and (_10316_, _10315_, _10313_);
  or (_10317_, _10316_, _10312_);
  or (_10318_, _10317_, _05535_);
  and (_10319_, _10318_, _05542_);
  and (_10320_, _10319_, _10308_);
  or (_10321_, _10320_, _10297_);
  and (_10322_, _10321_, _09850_);
  and (_10323_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  and (_10325_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  or (_10326_, _10325_, _09792_);
  or (_10327_, _10326_, _10323_);
  and (_10328_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  and (_10329_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  or (_10330_, _10329_, _05549_);
  or (_10331_, _10330_, _10328_);
  and (_10332_, _10331_, _10327_);
  or (_10333_, _10332_, _09791_);
  and (_10334_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  and (_10335_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  or (_10336_, _10335_, _09792_);
  or (_10338_, _10336_, _10334_);
  and (_10339_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  and (_10340_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  or (_10341_, _10340_, _05549_);
  or (_10342_, _10341_, _10339_);
  and (_10343_, _10342_, _10338_);
  or (_10344_, _10343_, _05535_);
  and (_10345_, _10344_, _09805_);
  and (_10346_, _10345_, _10333_);
  or (_10348_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  or (_10349_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  and (_10350_, _10349_, _10348_);
  or (_10351_, _10350_, _05549_);
  or (_10352_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  or (_10353_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  and (_10354_, _10353_, _10352_);
  or (_10355_, _10354_, _09792_);
  and (_10356_, _10355_, _10351_);
  or (_10357_, _10356_, _09791_);
  or (_10359_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  or (_10360_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  and (_10361_, _10360_, _10359_);
  or (_10362_, _10361_, _05549_);
  or (_10363_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_10364_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  and (_10365_, _10364_, _10363_);
  or (_10367_, _10365_, _09792_);
  and (_10368_, _10367_, _10362_);
  or (_10369_, _10368_, _05535_);
  and (_10370_, _10369_, _05542_);
  and (_10371_, _10370_, _10357_);
  or (_10372_, _10371_, _10346_);
  and (_10373_, _10372_, _05518_);
  or (_10374_, _10373_, _10322_);
  and (_10376_, _10374_, _09790_);
  and (_10377_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  and (_10378_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  or (_10380_, _10378_, _10377_);
  and (_10381_, _10380_, _09792_);
  and (_10383_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  and (_10384_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  or (_10385_, _10384_, _10383_);
  and (_10386_, _10385_, _05549_);
  or (_10387_, _10386_, _10381_);
  and (_10388_, _10387_, _05535_);
  and (_10389_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  and (_10390_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  or (_10391_, _10390_, _10389_);
  and (_10392_, _10391_, _09792_);
  and (_10393_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  and (_10394_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  or (_10395_, _10394_, _10393_);
  and (_10396_, _10395_, _05549_);
  or (_10397_, _10396_, _10392_);
  and (_10398_, _10397_, _09791_);
  or (_10399_, _10398_, _10388_);
  and (_10400_, _10399_, _09805_);
  or (_10401_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  or (_10402_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  and (_10403_, _10402_, _10401_);
  and (_10404_, _10403_, _09792_);
  or (_10405_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  or (_10406_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  and (_10407_, _10406_, _10405_);
  and (_10408_, _10407_, _05549_);
  or (_10409_, _10408_, _10404_);
  and (_10410_, _10409_, _05535_);
  or (_10411_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  or (_10412_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  and (_10413_, _10412_, _10411_);
  and (_10414_, _10413_, _09792_);
  or (_10415_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  or (_10416_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  and (_10417_, _10416_, _10415_);
  and (_10418_, _10417_, _05549_);
  or (_10419_, _10418_, _10414_);
  and (_10421_, _10419_, _09791_);
  or (_10422_, _10421_, _10410_);
  and (_10423_, _10422_, _05542_);
  or (_10424_, _10423_, _10400_);
  and (_10425_, _10424_, _09850_);
  and (_10426_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  and (_10427_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or (_10429_, _10427_, _10426_);
  and (_10430_, _10429_, _09792_);
  and (_10432_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  and (_10433_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or (_10435_, _10433_, _10432_);
  and (_10436_, _10435_, _05549_);
  or (_10437_, _10436_, _10430_);
  and (_10438_, _10437_, _05535_);
  and (_10439_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  and (_10440_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or (_10441_, _10440_, _10439_);
  and (_10443_, _10441_, _09792_);
  and (_10444_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  and (_10445_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or (_10447_, _10445_, _10444_);
  and (_10448_, _10447_, _05549_);
  or (_10449_, _10448_, _10443_);
  and (_10450_, _10449_, _09791_);
  or (_10451_, _10450_, _10438_);
  and (_10452_, _10451_, _09805_);
  or (_10453_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or (_10455_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  and (_10456_, _10455_, _10453_);
  and (_10457_, _10456_, _09792_);
  or (_10458_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or (_10459_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  and (_10462_, _10459_, _10458_);
  and (_10463_, _10462_, _05549_);
  or (_10464_, _10463_, _10457_);
  and (_10465_, _10464_, _05535_);
  or (_10466_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or (_10467_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  and (_10468_, _10467_, _10466_);
  and (_10469_, _10468_, _09792_);
  or (_10470_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  or (_10471_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  and (_10472_, _10471_, _10470_);
  and (_10473_, _10472_, _05549_);
  or (_10474_, _10473_, _10469_);
  and (_10475_, _10474_, _09791_);
  or (_10476_, _10475_, _10465_);
  and (_10477_, _10476_, _05542_);
  or (_10478_, _10477_, _10452_);
  and (_10479_, _10478_, _05518_);
  or (_10480_, _10479_, _10425_);
  and (_10481_, _10480_, _05520_);
  or (_10483_, _10481_, _10376_);
  or (_10484_, _10483_, _05526_);
  and (_10485_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  and (_10486_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_10487_, _10486_, _10485_);
  and (_10488_, _10487_, _09792_);
  and (_10489_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  and (_10490_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  or (_10491_, _10490_, _10489_);
  and (_10492_, _10491_, _05549_);
  or (_10493_, _10492_, _10488_);
  or (_10494_, _10493_, _09791_);
  and (_10495_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  and (_10496_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  or (_10497_, _10496_, _10495_);
  and (_10498_, _10497_, _09792_);
  and (_10499_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  and (_10500_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  or (_10501_, _10500_, _10499_);
  and (_10502_, _10501_, _05549_);
  or (_10503_, _10502_, _10498_);
  or (_10504_, _10503_, _05535_);
  and (_10505_, _10504_, _09805_);
  and (_10507_, _10505_, _10494_);
  or (_10509_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  or (_10510_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  and (_10511_, _10510_, _05549_);
  and (_10512_, _10511_, _10509_);
  or (_10514_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  or (_10515_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  and (_10517_, _10515_, _09792_);
  and (_10518_, _10517_, _10514_);
  or (_10519_, _10518_, _10512_);
  or (_10520_, _10519_, _09791_);
  or (_10521_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  or (_10522_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  and (_10524_, _10522_, _05549_);
  and (_10525_, _10524_, _10521_);
  or (_10526_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  or (_10527_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  and (_10529_, _10527_, _09792_);
  and (_10530_, _10529_, _10526_);
  or (_10531_, _10530_, _10525_);
  or (_10532_, _10531_, _05535_);
  and (_10533_, _10532_, _05542_);
  and (_10535_, _10533_, _10520_);
  or (_10536_, _10535_, _10507_);
  and (_10537_, _10536_, _09850_);
  and (_10538_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  and (_10540_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_10542_, _10540_, _10538_);
  and (_10543_, _10542_, _09792_);
  and (_10544_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  and (_10545_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or (_10546_, _10545_, _10544_);
  and (_10547_, _10546_, _05549_);
  or (_10548_, _10547_, _10543_);
  or (_10549_, _10548_, _09791_);
  and (_10550_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  and (_10552_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or (_10553_, _10552_, _10550_);
  and (_10554_, _10553_, _09792_);
  and (_10555_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  and (_10556_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  or (_10557_, _10556_, _10555_);
  and (_10558_, _10557_, _05549_);
  or (_10559_, _10558_, _10554_);
  or (_10561_, _10559_, _05535_);
  and (_10563_, _10561_, _09805_);
  and (_10564_, _10563_, _10549_);
  or (_10566_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or (_10567_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  and (_10568_, _10567_, _10566_);
  and (_10570_, _10568_, _09792_);
  or (_10571_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_10573_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  and (_10575_, _10573_, _10571_);
  and (_10576_, _10575_, _05549_);
  or (_10578_, _10576_, _10570_);
  or (_10579_, _10578_, _09791_);
  or (_10580_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  or (_10581_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  and (_10582_, _10581_, _10580_);
  and (_10584_, _10582_, _09792_);
  or (_10585_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_10586_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  and (_10587_, _10586_, _10585_);
  and (_10588_, _10587_, _05549_);
  or (_10590_, _10588_, _10584_);
  or (_10591_, _10590_, _05535_);
  and (_10593_, _10591_, _05542_);
  and (_10594_, _10593_, _10579_);
  or (_10595_, _10594_, _10564_);
  and (_10596_, _10595_, _05518_);
  or (_10597_, _10596_, _10537_);
  and (_10598_, _10597_, _09790_);
  or (_10600_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  or (_10602_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and (_10603_, _10602_, _10600_);
  and (_10604_, _10603_, _09792_);
  or (_10605_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  or (_10606_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_10608_, _10606_, _10605_);
  and (_10610_, _10608_, _05549_);
  or (_10611_, _10610_, _10604_);
  and (_10612_, _10611_, _09791_);
  or (_10614_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  or (_10615_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and (_10616_, _10615_, _10614_);
  and (_10617_, _10616_, _09792_);
  or (_10619_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  or (_10621_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_10623_, _10621_, _10619_);
  and (_10625_, _10623_, _05549_);
  or (_10626_, _10625_, _10617_);
  and (_10627_, _10626_, _05535_);
  or (_10628_, _10627_, _10612_);
  and (_10629_, _10628_, _05542_);
  and (_10631_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  and (_10632_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  or (_10633_, _10632_, _10631_);
  and (_10634_, _10633_, _09792_);
  and (_10635_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  and (_10636_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  or (_10637_, _10636_, _10635_);
  and (_10638_, _10637_, _05549_);
  or (_10640_, _10638_, _10634_);
  and (_10641_, _10640_, _09791_);
  and (_10642_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  and (_10643_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  or (_10644_, _10643_, _10642_);
  and (_10646_, _10644_, _09792_);
  and (_10647_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  and (_10649_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  or (_10651_, _10649_, _10647_);
  and (_10652_, _10651_, _05549_);
  or (_10654_, _10652_, _10646_);
  and (_10655_, _10654_, _05535_);
  or (_10657_, _10655_, _10641_);
  and (_10659_, _10657_, _09805_);
  or (_10660_, _10659_, _10629_);
  and (_10661_, _10660_, _05518_);
  or (_10662_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_10663_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  and (_10664_, _10663_, _05549_);
  and (_10665_, _10664_, _10662_);
  or (_10666_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or (_10667_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  and (_10669_, _10667_, _09792_);
  and (_10670_, _10669_, _10666_);
  or (_10672_, _10670_, _10665_);
  and (_10673_, _10672_, _09791_);
  or (_10674_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  or (_10676_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  and (_10677_, _10676_, _05549_);
  and (_10678_, _10677_, _10674_);
  or (_10679_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or (_10680_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  and (_10682_, _10680_, _09792_);
  and (_10683_, _10682_, _10679_);
  or (_10684_, _10683_, _10678_);
  and (_10685_, _10684_, _05535_);
  or (_10687_, _10685_, _10673_);
  and (_10689_, _10687_, _05542_);
  and (_10691_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  and (_10693_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_10695_, _10693_, _10691_);
  and (_10697_, _10695_, _09792_);
  and (_10698_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  and (_10699_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_10700_, _10699_, _10698_);
  and (_10701_, _10700_, _05549_);
  or (_10702_, _10701_, _10697_);
  and (_10704_, _10702_, _09791_);
  and (_10706_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  and (_10707_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_10708_, _10707_, _10706_);
  and (_10709_, _10708_, _09792_);
  and (_10710_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  and (_10712_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or (_10714_, _10712_, _10710_);
  and (_10715_, _10714_, _05549_);
  or (_10717_, _10715_, _10709_);
  and (_10718_, _10717_, _05535_);
  or (_10719_, _10718_, _10704_);
  and (_10721_, _10719_, _09805_);
  or (_10722_, _10721_, _10689_);
  and (_10724_, _10722_, _09850_);
  or (_10725_, _10724_, _10661_);
  and (_10726_, _10725_, _05520_);
  or (_10728_, _10726_, _10598_);
  or (_10729_, _10728_, _10033_);
  and (_10730_, _10729_, _10484_);
  or (_10731_, _10730_, _04413_);
  and (_10732_, _10731_, _10274_);
  or (_10733_, _10732_, _05563_);
  not (_10735_, _05563_);
  or (_10737_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_10738_, _10737_, _22731_);
  and (_27313_[6], _10738_, _10733_);
  and (_10740_, _09774_, _24089_);
  and (_10741_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  or (_03297_, _10741_, _10740_);
  and (_10742_, _03026_, _23548_);
  and (_10743_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_03300_, _10743_, _10742_);
  and (_10744_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  and (_10745_, _04853_, _23548_);
  or (_03321_, _10745_, _10744_);
  and (_10746_, _24408_, _24372_);
  and (_10748_, _10746_, _24219_);
  not (_10749_, _10746_);
  and (_10750_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  or (_03336_, _10750_, _10748_);
  and (_10751_, _24408_, _24146_);
  and (_10752_, _10751_, _23996_);
  not (_10754_, _10751_);
  and (_10755_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  or (_03339_, _10755_, _10752_);
  and (_10756_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  and (_10757_, _04853_, _24219_);
  or (_03342_, _10757_, _10756_);
  and (_10758_, _10751_, _24089_);
  and (_10759_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  or (_03345_, _10759_, _10758_);
  and (_10760_, _10751_, _24219_);
  and (_10761_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  or (_03352_, _10761_, _10760_);
  and (_10762_, _24408_, _24140_);
  and (_10763_, _10762_, _24134_);
  not (_10765_, _10762_);
  and (_10766_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  or (_27113_, _10766_, _10763_);
  and (_10767_, _10762_, _23548_);
  and (_10768_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_27111_, _10768_, _10767_);
  and (_10769_, _02512_, _24159_);
  not (_10770_, _10769_);
  and (_10771_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  and (_10772_, _10769_, _24219_);
  or (_03389_, _10772_, _10771_);
  and (_10773_, _02512_, _24297_);
  not (_10774_, _10773_);
  and (_10775_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and (_10776_, _10773_, _23996_);
  or (_03399_, _10776_, _10775_);
  and (_10777_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_10778_, _10773_, _23583_);
  or (_03401_, _10778_, _10777_);
  and (_10779_, _09780_, _23548_);
  and (_10781_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or (_03415_, _10781_, _10779_);
  and (_10782_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_10783_, _04897_, _23583_);
  or (_03418_, _10783_, _10782_);
  and (_10784_, _09780_, _24219_);
  and (_10785_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or (_03422_, _10785_, _10784_);
  and (_10786_, _05465_, _24134_);
  and (_10787_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  or (_03426_, _10787_, _10786_);
  and (_10788_, _02512_, _24016_);
  not (_10789_, _10788_);
  and (_10790_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and (_10791_, _10788_, _23583_);
  or (_03427_, _10791_, _10790_);
  and (_10792_, _02512_, _24236_);
  not (_10793_, _10792_);
  and (_10794_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  and (_10795_, _10792_, _23996_);
  or (_27105_, _10795_, _10794_);
  and (_10797_, _09779_, _24297_);
  and (_10798_, _10797_, _23996_);
  not (_10799_, _10797_);
  and (_10800_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  or (_03440_, _10800_, _10798_);
  and (_10801_, _24451_, _23887_);
  and (_10802_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_03443_, _10802_, _10801_);
  and (_10803_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  and (_10804_, _10792_, _24089_);
  or (_27104_, _10804_, _10803_);
  and (_10805_, _02512_, _23941_);
  not (_10806_, _10805_);
  and (_10807_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_10808_, _10805_, _23996_);
  or (_03456_, _10808_, _10807_);
  and (_10809_, _02512_, _24899_);
  not (_10811_, _10809_);
  and (_10813_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and (_10815_, _10809_, _23996_);
  or (_03467_, _10815_, _10813_);
  and (_10816_, _09780_, _24089_);
  and (_10817_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or (_03472_, _10817_, _10816_);
  and (_10819_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_10821_, _10809_, _23887_);
  or (_03475_, _10821_, _10819_);
  and (_10822_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and (_10823_, _10809_, _24219_);
  or (_03477_, _10823_, _10822_);
  and (_10824_, _09780_, _23583_);
  and (_10825_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or (_03480_, _10825_, _10824_);
  and (_10827_, _02512_, _24474_);
  not (_10829_, _10827_);
  and (_10830_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  and (_10832_, _10827_, _23996_);
  or (_03483_, _10832_, _10830_);
  and (_10834_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  and (_10835_, _10827_, _23548_);
  or (_03486_, _10835_, _10834_);
  and (_10836_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  and (_10837_, _10792_, _23548_);
  or (_27101_, _10837_, _10836_);
  and (_10839_, _02512_, _24349_);
  not (_10840_, _10839_);
  and (_10841_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  and (_10843_, _10839_, _24134_);
  or (_03498_, _10843_, _10841_);
  and (_10845_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  and (_10846_, _10839_, _23583_);
  or (_03507_, _10846_, _10845_);
  and (_10847_, _10746_, _23887_);
  and (_10848_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  or (_03509_, _10848_, _10847_);
  and (_10849_, _09774_, _23583_);
  and (_10850_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or (_03511_, _10850_, _10849_);
  and (_10851_, _10762_, _23583_);
  and (_10852_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_03519_, _10852_, _10851_);
  and (_10854_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  and (_10855_, _10769_, _24051_);
  or (_03529_, _10855_, _10854_);
  and (_10856_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  and (_10858_, _10769_, _23887_);
  or (_03533_, _10858_, _10856_);
  and (_10859_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_10860_, _10773_, _24219_);
  or (_27108_, _10860_, _10859_);
  and (_10861_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and (_10862_, _10788_, _24051_);
  or (_03539_, _10862_, _10861_);
  and (_10863_, _10797_, _23583_);
  and (_10865_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  or (_27002_, _10865_, _10863_);
  and (_10867_, _24140_, _22982_);
  and (_10868_, _10867_, _24089_);
  not (_10869_, _10867_);
  and (_10871_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  or (_03548_, _10871_, _10868_);
  and (_10872_, _10797_, _23887_);
  and (_10873_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  or (_03553_, _10873_, _10872_);
  and (_10874_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and (_10875_, _10805_, _23887_);
  or (_03560_, _10875_, _10874_);
  and (_10876_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  and (_10877_, _10827_, _23583_);
  or (_03573_, _10877_, _10876_);
  and (_10878_, _24302_, _23583_);
  and (_10879_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  or (_03576_, _10879_, _10878_);
  and (_10880_, _09670_, _23583_);
  and (_10882_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  or (_03584_, _10882_, _10880_);
  and (_10884_, _10762_, _23996_);
  and (_10885_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_03598_, _10885_, _10884_);
  and (_10887_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and (_10888_, _10773_, _24089_);
  or (_03605_, _10888_, _10887_);
  and (_10889_, _06763_, _24134_);
  and (_10890_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  or (_03609_, _10890_, _10889_);
  and (_10892_, _10797_, _24134_);
  and (_10894_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  or (_27004_, _10894_, _10892_);
  and (_10895_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and (_10896_, _10809_, _24089_);
  or (_03627_, _10896_, _10895_);
  and (_10898_, _10797_, _24051_);
  and (_10900_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  or (_27003_, _10900_, _10898_);
  and (_10902_, _10797_, _24089_);
  and (_10903_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  or (_03631_, _10903_, _10902_);
  and (_10904_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and (_10905_, _06203_, _24051_);
  or (_03648_, _10905_, _10904_);
  and (_10906_, _09779_, _24016_);
  and (_10907_, _10906_, _24089_);
  not (_10908_, _10906_);
  and (_10909_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  or (_03659_, _10909_, _10907_);
  and (_10911_, _03026_, _24219_);
  and (_10912_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_03664_, _10912_, _10911_);
  and (_10913_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  and (_10914_, _10839_, _23887_);
  or (_03671_, _10914_, _10913_);
  and (_10916_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  and (_10917_, _10839_, _24219_);
  or (_03673_, _10917_, _10916_);
  and (_10919_, _03186_, _23548_);
  and (_10920_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  or (_03675_, _10920_, _10919_);
  and (_10922_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  and (_10924_, _10839_, _23548_);
  or (_27098_, _10924_, _10922_);
  and (_10926_, _03186_, _23887_);
  and (_10927_, _03188_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  or (_27050_, _10927_, _10926_);
  and (_10929_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  and (_10930_, _10839_, _24089_);
  or (_03695_, _10930_, _10929_);
  and (_10931_, _10906_, _24134_);
  and (_10932_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  or (_03697_, _10932_, _10931_);
  and (_10935_, _03026_, _24089_);
  and (_10937_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_03701_, _10937_, _10935_);
  and (_10939_, _03026_, _23887_);
  and (_10940_, _03029_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_03704_, _10940_, _10939_);
  and (_10943_, _10906_, _24051_);
  and (_10945_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  or (_03716_, _10945_, _10943_);
  and (_10947_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  and (_10949_, _10839_, _24051_);
  or (_03718_, _10949_, _10947_);
  and (_26841_[1], _26769_, _22731_);
  and (_10952_, _10840_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  and (_10954_, _10839_, _23996_);
  or (_03726_, _10954_, _10952_);
  and (_10956_, _02990_, _23887_);
  and (_10957_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  or (_27054_, _10957_, _10956_);
  or (_10959_, _02351_, _04800_);
  and (_10961_, _10959_, _22737_);
  and (_10962_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_10963_, _10962_, _02360_);
  or (_10965_, _10963_, _02010_);
  or (_10966_, _10965_, _10961_);
  and (_26849_[2], _10966_, _22731_);
  and (_10969_, _02990_, _24134_);
  and (_10971_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  or (_03741_, _10971_, _10969_);
  and (_10972_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  and (_10973_, _10792_, _24219_);
  or (_03749_, _10973_, _10972_);
  and (_10975_, _02990_, _24051_);
  and (_10977_, _02992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  or (_03753_, _10977_, _10975_);
  and (_10979_, _23890_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and (_10981_, _23892_, _23779_);
  or (_10983_, _09762_, _23923_);
  or (_10985_, _10983_, _10981_);
  or (_10986_, _23839_, _23793_);
  or (_10988_, _10986_, _26739_);
  or (_10989_, _10988_, _10985_);
  or (_10990_, _10989_, _09753_);
  and (_10991_, _10990_, _23855_);
  or (_26850_[1], _10991_, _10979_);
  and (_10992_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  and (_10994_, _10827_, _24219_);
  or (_03761_, _10994_, _10992_);
  and (_10996_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and (_10997_, _06203_, _24089_);
  or (_03766_, _10997_, _10996_);
  and (_10998_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  and (_11000_, _10827_, _23887_);
  or (_03768_, _11000_, _10998_);
  and (_11002_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  and (_11003_, _10827_, _24089_);
  or (_03780_, _11003_, _11002_);
  and (_11004_, _02339_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  and (_11006_, _02338_, _24051_);
  or (_27027_, _11006_, _11004_);
  and (_11007_, _09717_, _24219_);
  and (_11008_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_27070_, _11008_, _11007_);
  and (_11009_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  and (_11010_, _10827_, _24051_);
  or (_03800_, _11010_, _11009_);
  and (_11012_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_11013_, _02040_, _24219_);
  or (_03804_, _11013_, _11012_);
  and (_11015_, _02041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  and (_11016_, _02040_, _24134_);
  or (_03812_, _11016_, _11015_);
  and (_11018_, _10829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  and (_11019_, _10827_, _24134_);
  or (_03817_, _11019_, _11018_);
  and (_11020_, _10797_, _24219_);
  and (_11022_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  or (_03820_, _11022_, _11020_);
  and (_11025_, _25648_, _24219_);
  and (_11026_, _25650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  or (_03827_, _11026_, _11025_);
  and (_11028_, _10906_, _23996_);
  and (_11029_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  or (_03836_, _11029_, _11028_);
  and (_11031_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and (_11032_, _10809_, _23548_);
  or (_03848_, _11032_, _11031_);
  and (_11033_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and (_11034_, _06203_, _23583_);
  or (_27088_, _11034_, _11033_);
  and (_11037_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and (_11038_, _10809_, _23583_);
  or (_03854_, _11038_, _11037_);
  and (_11040_, _25442_, _23548_);
  and (_11041_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_03856_, _11041_, _11040_);
  and (_11044_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and (_11045_, _10809_, _24051_);
  or (_03864_, _11045_, _11044_);
  and (_11046_, _09779_, _24236_);
  and (_11047_, _11046_, _24134_);
  not (_11049_, _11046_);
  and (_11051_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  or (_03867_, _11051_, _11047_);
  and (_11052_, _11046_, _23996_);
  and (_11053_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or (_03900_, _11053_, _11052_);
  and (_11054_, _25442_, _24051_);
  and (_11055_, _25444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_03907_, _11055_, _11054_);
  and (_11057_, _10811_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  and (_11058_, _10809_, _24134_);
  or (_03918_, _11058_, _11057_);
  and (_11059_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_11060_, _10805_, _24219_);
  or (_03921_, _11060_, _11059_);
  and (_11061_, _25206_, _23996_);
  and (_11062_, _25208_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_03924_, _11062_, _11061_);
  and (_11063_, _09717_, _23548_);
  and (_11064_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_03932_, _11064_, _11063_);
  and (_11065_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and (_11066_, _10805_, _23548_);
  or (_03948_, _11066_, _11065_);
  and (_11067_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_11069_, _10805_, _23583_);
  or (_27097_, _11069_, _11067_);
  and (_11070_, _10867_, _24051_);
  and (_11072_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  or (_27262_, _11072_, _11070_);
  and (_11073_, _24415_, _23548_);
  and (_11075_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  or (_03961_, _11075_, _11073_);
  and (_11078_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_11079_, _10805_, _24089_);
  or (_03969_, _11079_, _11078_);
  and (_11080_, _24381_, _23548_);
  and (_11082_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_03971_, _11082_, _11080_);
  and (_11083_, _10906_, _23887_);
  and (_11084_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  or (_03974_, _11084_, _11083_);
  and (_11086_, _24415_, _23996_);
  and (_11087_, _24417_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  or (_03986_, _11087_, _11086_);
  and (_11089_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and (_11090_, _10805_, _24051_);
  or (_03989_, _11090_, _11089_);
  or (_11092_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_03992_, _11092_, _03428_);
  and (_11093_, _24381_, _23996_);
  and (_11094_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_03994_, _11094_, _11093_);
  and (_11095_, _10906_, _23548_);
  and (_11096_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  or (_27001_, _11096_, _11095_);
  and (_11097_, _24381_, _24089_);
  and (_11098_, _24383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_03999_, _11098_, _11097_);
  not (_11099_, _02294_);
  or (_11100_, _11099_, _23577_);
  and (_11101_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_11102_, _02257_, _02248_);
  nor (_11104_, _11102_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_11105_, _11104_, _06159_);
  and (_11107_, _11105_, _06158_);
  and (_11108_, _02623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_11110_, _11108_, _11107_);
  nor (_11112_, _11110_, _02616_);
  or (_11114_, _11112_, _11101_);
  or (_11116_, _11114_, _02294_);
  and (_11118_, _11116_, _22731_);
  and (_04002_, _11118_, _11100_);
  and (_11119_, _24330_, _24051_);
  and (_11120_, _24332_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_04005_, _11120_, _11119_);
  and (_11122_, _10806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  and (_11123_, _10805_, _24134_);
  or (_04007_, _11123_, _11122_);
  nor (_11125_, _24210_, rst);
  or (_11127_, _11125_, _02295_);
  and (_11129_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_11130_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_11131_, _11130_, _02283_);
  and (_11132_, _11131_, _02263_);
  and (_11134_, _02248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_11136_, _02248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_11137_, _11136_, _11134_);
  and (_11138_, _11137_, _06158_);
  nor (_11139_, _11138_, _11132_);
  nor (_11140_, _11139_, _02616_);
  or (_11141_, _11140_, _02294_);
  or (_11143_, _11141_, _11129_);
  and (_04010_, _11143_, _11127_);
  and (_11145_, _10906_, _24219_);
  and (_11147_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  or (_04013_, _11147_, _11145_);
  not (_11148_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_11149_, _02620_, _02237_);
  and (_11150_, _06162_, _02271_);
  nor (_11151_, _11150_, _11149_);
  and (_11152_, _11151_, _11148_);
  nor (_11153_, _11151_, _11148_);
  nor (_11154_, _11153_, _11152_);
  or (_11155_, _11154_, _02616_);
  nand (_11157_, _02616_, _24210_);
  and (_11158_, _11157_, _11155_);
  and (_11159_, _11158_, _02295_);
  and (_11160_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or (_04015_, _11160_, _11159_);
  and (_11163_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  and (_11164_, _10792_, _23887_);
  or (_27102_, _11164_, _11163_);
  and (_11165_, _24350_, _24219_);
  and (_11166_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_04026_, _11166_, _11165_);
  or (_11168_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_26894_, _11168_, _03087_);
  and (_11169_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  and (_11171_, _10792_, _23583_);
  or (_27103_, _11171_, _11169_);
  and (_11174_, _24134_, _23946_);
  and (_11175_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  or (_04037_, _11175_, _11174_);
  and (_11177_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  and (_11179_, _10792_, _24051_);
  or (_04040_, _11179_, _11177_);
  or (_11181_, _02300_, _23577_);
  nand (_11182_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_11183_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_11184_, _02206_, _02205_);
  and (_11185_, _11184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nand (_11186_, _11185_, _11183_);
  and (_11187_, _11186_, _11182_);
  nor (_11189_, _11187_, _01814_);
  and (_11191_, _02207_, _11184_);
  nand (_11193_, _11191_, _02193_);
  and (_11194_, _11193_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_11195_, _11194_, _11189_);
  or (_11196_, _11195_, _01816_);
  and (_11198_, _11196_, _22731_);
  and (_04044_, _11198_, _11181_);
  or (_11201_, _02193_, _23880_);
  and (_11203_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_11205_, _11203_, _08224_);
  and (_11206_, _11205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_11207_, _11206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_11208_, _11206_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_11209_, _11208_, _02197_);
  and (_11210_, _11209_, _11207_);
  and (_11211_, _02210_, _01820_);
  or (_11212_, _11211_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_11214_, _11211_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_11216_, _11214_, _02320_);
  and (_11217_, _11216_, _11212_);
  and (_11218_, _01821_, _01818_);
  nand (_11219_, _11218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_11221_, _01820_, _01818_);
  and (_11223_, _11221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_11225_, _11223_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_11226_, _11225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_11227_, _11226_, _11219_);
  or (_11229_, _11227_, _11217_);
  or (_11230_, _11229_, _11210_);
  or (_11231_, _11230_, _01814_);
  and (_11233_, _11231_, _11201_);
  or (_11235_, _11233_, _01816_);
  or (_11236_, _02300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_11238_, _11236_, _22731_);
  and (_04046_, _11238_, _11235_);
  and (_11239_, _24237_, _23887_);
  and (_11241_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_04050_, _11241_, _11239_);
  and (_11243_, _11046_, _24219_);
  and (_11244_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or (_04055_, _11244_, _11243_);
  and (_11245_, _10793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  and (_11246_, _10792_, _24134_);
  or (_04068_, _11246_, _11245_);
  and (_11247_, _24237_, _24219_);
  and (_11248_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_04072_, _11248_, _11247_);
  and (_11250_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and (_11251_, _10788_, _24219_);
  or (_27106_, _11251_, _11250_);
  or (_11252_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_04075_, _11252_, _03414_);
  or (_11253_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_11254_, _11253_, _22731_);
  not (_11256_, _24189_);
  or (_11257_, _11256_, _23880_);
  and (_04077_, _11257_, _11254_);
  and (_11259_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and (_11260_, _10788_, _23548_);
  or (_04087_, _11260_, _11259_);
  and (_11261_, _24017_, _23996_);
  and (_11263_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  or (_04089_, _11263_, _11261_);
  and (_11264_, _09779_, _24349_);
  and (_11265_, _11264_, _23996_);
  not (_11266_, _11264_);
  and (_11267_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or (_04092_, _11267_, _11265_);
  and (_11269_, _24089_, _24017_);
  and (_11270_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  or (_04097_, _11270_, _11269_);
  or (_11271_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_04101_, _11271_, _03419_);
  and (_11272_, _05465_, _24051_);
  and (_11273_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  or (_04107_, _11273_, _11272_);
  and (_11274_, _11264_, _24134_);
  and (_11275_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  or (_04109_, _11275_, _11274_);
  and (_11276_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and (_11277_, _10788_, _23887_);
  or (_04112_, _11277_, _11276_);
  and (_11278_, _05465_, _23583_);
  and (_11279_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  or (_27068_, _11279_, _11278_);
  and (_11280_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_11281_, _10788_, _24089_);
  or (_04116_, _11281_, _11280_);
  and (_11282_, _09717_, _23583_);
  and (_11284_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_27071_, _11284_, _11282_);
  and (_11286_, _04865_, _23887_);
  and (_11288_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or (_04126_, _11288_, _11286_);
  and (_11290_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  and (_11291_, _10788_, _24134_);
  or (_27107_, _11291_, _11290_);
  and (_11293_, _11046_, _23583_);
  and (_11295_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or (_04159_, _11295_, _11293_);
  and (_11297_, _10789_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_11299_, _10788_, _23996_);
  or (_04162_, _11299_, _11297_);
  and (_11301_, _11046_, _23887_);
  and (_11302_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or (_04165_, _11302_, _11301_);
  and (_11304_, _05460_, _24051_);
  and (_11306_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_04168_, _11306_, _11304_);
  and (_11307_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_11308_, _10773_, _23548_);
  or (_04171_, _11308_, _11307_);
  or (_11309_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_04174_, _11309_, _03408_);
  and (_11311_, _24372_, _24006_);
  and (_11312_, _11311_, _24219_);
  not (_11313_, _11311_);
  and (_11314_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  or (_04177_, _11314_, _11312_);
  and (_11316_, _24442_, _24051_);
  and (_11317_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  or (_27075_, _11317_, _11316_);
  and (_11318_, _11046_, _23548_);
  and (_11319_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or (_04185_, _11319_, _11318_);
  and (_11320_, _11311_, _23996_);
  and (_11321_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  or (_04187_, _11321_, _11320_);
  and (_11323_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and (_11324_, _10773_, _23887_);
  or (_04189_, _11324_, _11323_);
  and (_11325_, _11311_, _24089_);
  and (_11327_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  or (_04191_, _11327_, _11325_);
  and (_11329_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_11330_, _10773_, _24051_);
  or (_04194_, _11330_, _11329_);
  and (_11333_, _09717_, _23887_);
  and (_11335_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_04198_, _11335_, _11333_);
  and (_11337_, _07013_, _24089_);
  and (_11338_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_04200_, _11338_, _11337_);
  and (_11339_, _24889_, _24089_);
  and (_11340_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_04205_, _11340_, _11339_);
  and (_11341_, _10774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  and (_11342_, _10773_, _24134_);
  or (_04208_, _11342_, _11341_);
  and (_11343_, _24889_, _23887_);
  and (_11344_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_04218_, _11344_, _11343_);
  and (_11345_, _09774_, _23996_);
  and (_11346_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  or (_27242_, _11346_, _11345_);
  and (_11348_, _08578_, _23548_);
  and (_11349_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  or (_27076_, _11349_, _11348_);
  and (_11350_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  and (_11351_, _10769_, _23548_);
  or (_27109_, _11351_, _11350_);
  and (_11353_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  and (_11354_, _10769_, _23583_);
  or (_04254_, _11354_, _11353_);
  and (_11358_, _09774_, _24134_);
  and (_11359_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  or (_04262_, _11359_, _11358_);
  and (_11360_, _24056_, _24006_);
  and (_11361_, _11360_, _23583_);
  not (_11362_, _11360_);
  and (_11363_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_04269_, _11363_, _11361_);
  and (_11364_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  and (_11365_, _10769_, _24089_);
  or (_04271_, _11365_, _11364_);
  and (_11367_, _11264_, _23548_);
  and (_11368_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or (_04273_, _11368_, _11367_);
  and (_11370_, _11264_, _24219_);
  and (_11371_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or (_04279_, _11371_, _11370_);
  and (_11373_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  and (_11374_, _10769_, _24134_);
  or (_04282_, _11374_, _11373_);
  and (_11376_, _02964_, _23548_);
  and (_11377_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_04284_, _11377_, _11376_);
  and (_11378_, _11360_, _24134_);
  and (_11379_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  or (_04294_, _11379_, _11378_);
  and (_11381_, _02964_, _24219_);
  and (_11382_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_04296_, _11382_, _11381_);
  and (_11384_, _08523_, _23996_);
  and (_11385_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  or (_04299_, _11385_, _11384_);
  and (_11386_, _10770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  and (_11387_, _10769_, _23996_);
  or (_27110_, _11387_, _11386_);
  and (_11388_, _08523_, _24089_);
  and (_11389_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  or (_04307_, _11389_, _11388_);
  and (_11391_, _10762_, _24219_);
  and (_11392_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_04310_, _11392_, _11391_);
  and (_11393_, _06763_, _23583_);
  and (_11394_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_04313_, _11394_, _11393_);
  and (_11395_, _10762_, _23887_);
  and (_11396_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_04316_, _11396_, _11395_);
  and (_11397_, _24089_, _24008_);
  and (_11398_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_04318_, _11398_, _11397_);
  and (_11399_, _24008_, _23548_);
  and (_11400_, _24011_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_04321_, _11400_, _11399_);
  and (_11401_, _10762_, _24089_);
  and (_11402_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_04324_, _11402_, _11401_);
  and (_11403_, _02488_, _23583_);
  and (_11404_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  or (_04346_, _11404_, _11403_);
  and (_11405_, _02964_, _24134_);
  and (_11406_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  or (_04351_, _11406_, _11405_);
  and (_11409_, _02065_, _23887_);
  and (_11410_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  or (_04354_, _11410_, _11409_);
  and (_11412_, _10762_, _24051_);
  and (_11413_, _10765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_27112_, _11413_, _11412_);
  and (_11414_, _02488_, _23996_);
  and (_11415_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  or (_04359_, _11415_, _11414_);
  and (_11417_, _05442_, _23887_);
  and (_11418_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_04365_, _11418_, _11417_);
  and (_11419_, _24016_, _24006_);
  and (_11420_, _11419_, _23548_);
  not (_11421_, _11419_);
  and (_11422_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_04369_, _11422_, _11420_);
  and (_11423_, _05442_, _24089_);
  and (_11424_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_04371_, _11424_, _11423_);
  and (_11426_, _10751_, _23548_);
  and (_11427_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  or (_04381_, _11427_, _11426_);
  and (_11428_, _11264_, _24089_);
  and (_11429_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or (_04386_, _11429_, _11428_);
  and (_11430_, _02964_, _24089_);
  and (_11431_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_04391_, _11431_, _11430_);
  and (_11432_, _11264_, _23583_);
  and (_11433_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or (_26999_, _11433_, _11432_);
  and (_11434_, _11419_, _24051_);
  and (_11435_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or (_04398_, _11435_, _11434_);
  and (_11437_, _10751_, _23887_);
  and (_11438_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  or (_27114_, _11438_, _11437_);
  and (_11441_, _24297_, _24006_);
  and (_11443_, _11441_, _24089_);
  not (_11444_, _11441_);
  and (_11445_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_04408_, _11445_, _11443_);
  and (_11447_, _02964_, _23583_);
  and (_11448_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_04411_, _11448_, _11447_);
  and (_11449_, _02964_, _23887_);
  and (_11451_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_04415_, _11451_, _11449_);
  and (_11453_, _11441_, _23548_);
  and (_11454_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_04417_, _11454_, _11453_);
  and (_11456_, _23922_, _22737_);
  and (_11457_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_11458_, _11457_, _26680_);
  or (_11459_, _11458_, _11456_);
  and (_26852_[1], _11459_, _22731_);
  and (_11460_, _06763_, _24051_);
  and (_11461_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or (_04422_, _11461_, _11460_);
  and (_11464_, _10751_, _23583_);
  and (_11465_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  or (_04424_, _11465_, _11464_);
  and (_11467_, _11264_, _23887_);
  and (_11468_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or (_26998_, _11468_, _11467_);
  and (_11469_, _08435_, _24219_);
  and (_11470_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  or (_04432_, _11470_, _11469_);
  and (_11471_, _23890_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_11472_, _23819_, _23809_);
  or (_11473_, _04789_, _23929_);
  or (_11474_, _11473_, _23836_);
  or (_11476_, _11474_, _23828_);
  or (_11477_, _11476_, _03919_);
  or (_11478_, _04796_, _26731_);
  or (_11479_, _11478_, _24276_);
  or (_11480_, _11479_, _24262_);
  or (_11481_, _11480_, _11477_);
  or (_11482_, _11481_, _11472_);
  and (_11483_, _11482_, _23855_);
  or (_26851_[3], _11483_, _11471_);
  and (_11484_, _06204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_11485_, _06203_, _24219_);
  or (_04445_, _11485_, _11484_);
  and (_11488_, _10751_, _24051_);
  and (_11489_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  or (_27115_, _11489_, _11488_);
  and (_11490_, _05438_, _23548_);
  and (_11491_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_04453_, _11491_, _11490_);
  and (_11492_, _10751_, _24134_);
  and (_11493_, _10754_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  or (_04455_, _11493_, _11492_);
  and (_11494_, _05438_, _23887_);
  and (_11495_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_04457_, _11495_, _11494_);
  and (_11497_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  and (_11498_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_11499_, _11498_, _11497_);
  and (_11500_, _11499_, _09792_);
  and (_11501_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  and (_11502_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_11503_, _11502_, _11501_);
  and (_11504_, _11503_, _05549_);
  or (_11505_, _11504_, _11500_);
  or (_11506_, _11505_, _09791_);
  and (_11507_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  and (_11508_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_11509_, _11508_, _11507_);
  and (_11511_, _11509_, _09792_);
  and (_11513_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  and (_11515_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  or (_11516_, _11515_, _11513_);
  and (_11518_, _11516_, _05549_);
  or (_11520_, _11518_, _11511_);
  or (_11521_, _11520_, _05535_);
  and (_11522_, _11521_, _09805_);
  and (_11523_, _11522_, _11506_);
  or (_11524_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_11525_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  and (_11527_, _11525_, _11524_);
  and (_11529_, _11527_, _09792_);
  or (_11530_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_11531_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  and (_11532_, _11531_, _11530_);
  and (_11533_, _11532_, _05549_);
  or (_11534_, _11533_, _11529_);
  or (_11535_, _11534_, _09791_);
  or (_11536_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  or (_11537_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  and (_11538_, _11537_, _11536_);
  and (_11540_, _11538_, _09792_);
  or (_11541_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  or (_11542_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  and (_11543_, _11542_, _11541_);
  and (_11544_, _11543_, _05549_);
  or (_11545_, _11544_, _11540_);
  or (_11546_, _11545_, _05535_);
  and (_11547_, _11546_, _05542_);
  and (_11548_, _11547_, _11535_);
  or (_11549_, _11548_, _11523_);
  and (_11551_, _11549_, _05518_);
  and (_11552_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  and (_11554_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  or (_11555_, _11554_, _11552_);
  and (_11556_, _11555_, _09792_);
  and (_11557_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  and (_11558_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  or (_11559_, _11558_, _11557_);
  and (_11560_, _11559_, _05549_);
  or (_11561_, _11560_, _11556_);
  or (_11562_, _11561_, _09791_);
  and (_11564_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  and (_11565_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  or (_11566_, _11565_, _11564_);
  and (_11567_, _11566_, _09792_);
  and (_11568_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  and (_11569_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_11570_, _11569_, _11568_);
  and (_11571_, _11570_, _05549_);
  or (_11572_, _11571_, _11567_);
  or (_11573_, _11572_, _05535_);
  and (_11574_, _11573_, _09805_);
  and (_11575_, _11574_, _11562_);
  or (_11576_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_11577_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  and (_11578_, _11577_, _05549_);
  and (_11579_, _11578_, _11576_);
  or (_11580_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  or (_11581_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  and (_11582_, _11581_, _09792_);
  and (_11583_, _11582_, _11580_);
  or (_11584_, _11583_, _11579_);
  or (_11585_, _11584_, _09791_);
  or (_11586_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_11587_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  and (_11588_, _11587_, _05549_);
  and (_11590_, _11588_, _11586_);
  or (_11591_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  or (_11593_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  and (_11595_, _11593_, _09792_);
  and (_11597_, _11595_, _11591_);
  or (_11598_, _11597_, _11590_);
  or (_11599_, _11598_, _05535_);
  and (_11600_, _11599_, _05542_);
  and (_11602_, _11600_, _11585_);
  or (_11604_, _11602_, _11575_);
  and (_11606_, _11604_, _09850_);
  or (_11607_, _11606_, _11551_);
  and (_11608_, _11607_, _09790_);
  and (_11609_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_11610_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_11612_, _11610_, _11609_);
  and (_11613_, _11612_, _09792_);
  and (_11615_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_11616_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_11617_, _11616_, _11615_);
  and (_11619_, _11617_, _05549_);
  or (_11620_, _11619_, _11613_);
  and (_11621_, _11620_, _05535_);
  and (_11622_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_11623_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_11624_, _11623_, _11622_);
  and (_11625_, _11624_, _09792_);
  and (_11626_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and (_11628_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_11629_, _11628_, _11626_);
  and (_11631_, _11629_, _05549_);
  or (_11633_, _11631_, _11625_);
  and (_11634_, _11633_, _09791_);
  or (_11635_, _11634_, _11621_);
  and (_11636_, _11635_, _09805_);
  or (_11637_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_11639_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_11640_, _11639_, _05549_);
  and (_11642_, _11640_, _11637_);
  or (_11643_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  or (_11645_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_11646_, _11645_, _09792_);
  and (_11647_, _11646_, _11643_);
  or (_11648_, _11647_, _11642_);
  and (_11649_, _11648_, _05535_);
  or (_11650_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_11651_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_11652_, _11651_, _05549_);
  and (_11653_, _11652_, _11650_);
  or (_11655_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_11657_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_11659_, _11657_, _09792_);
  and (_11660_, _11659_, _11655_);
  or (_11662_, _11660_, _11653_);
  and (_11663_, _11662_, _09791_);
  or (_11664_, _11663_, _11649_);
  and (_11665_, _11664_, _05542_);
  or (_11666_, _11665_, _11636_);
  and (_11667_, _11666_, _09850_);
  and (_11668_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  and (_11670_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  or (_11671_, _11670_, _11668_);
  and (_11672_, _11671_, _09792_);
  and (_11673_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  and (_11674_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  or (_11675_, _11674_, _11673_);
  and (_11676_, _11675_, _05549_);
  or (_11677_, _11676_, _11672_);
  and (_11678_, _11677_, _05535_);
  and (_11679_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  and (_11680_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_11681_, _11680_, _11679_);
  and (_11682_, _11681_, _09792_);
  and (_11683_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  and (_11684_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  or (_11686_, _11684_, _11683_);
  and (_11687_, _11686_, _05549_);
  or (_11689_, _11687_, _11682_);
  and (_11690_, _11689_, _09791_);
  or (_11692_, _11690_, _11678_);
  and (_11693_, _11692_, _09805_);
  or (_11695_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_11697_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  and (_11698_, _11697_, _11695_);
  and (_11700_, _11698_, _09792_);
  or (_11701_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_11702_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  and (_11703_, _11702_, _11701_);
  and (_11704_, _11703_, _05549_);
  or (_11705_, _11704_, _11700_);
  and (_11706_, _11705_, _05535_);
  or (_11707_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_11709_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  and (_11710_, _11709_, _11707_);
  and (_11712_, _11710_, _09792_);
  or (_11713_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_11715_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  and (_11717_, _11715_, _11713_);
  and (_11718_, _11717_, _05549_);
  or (_11719_, _11718_, _11712_);
  and (_11720_, _11719_, _09791_);
  or (_11722_, _11720_, _11706_);
  and (_11724_, _11722_, _05542_);
  or (_11725_, _11724_, _11693_);
  and (_11727_, _11725_, _05518_);
  or (_11729_, _11727_, _11667_);
  and (_11731_, _11729_, _05520_);
  or (_11732_, _11731_, _11608_);
  or (_11733_, _11732_, _05526_);
  and (_11735_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  and (_11737_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_11739_, _11737_, _11735_);
  and (_11741_, _11739_, _09792_);
  and (_11743_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  and (_11744_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_11745_, _11744_, _11743_);
  and (_11747_, _11745_, _05549_);
  or (_11748_, _11747_, _11741_);
  or (_11749_, _11748_, _09791_);
  and (_11751_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  and (_11753_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_11755_, _11753_, _11751_);
  and (_11756_, _11755_, _09792_);
  and (_11758_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  and (_11760_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_11762_, _11760_, _11758_);
  and (_11763_, _11762_, _05549_);
  or (_11764_, _11763_, _11756_);
  or (_11765_, _11764_, _05535_);
  and (_11766_, _11765_, _09805_);
  and (_11767_, _11766_, _11749_);
  or (_11768_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_11769_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  and (_11770_, _11769_, _05549_);
  and (_11771_, _11770_, _11768_);
  or (_11772_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_11773_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  and (_11774_, _11773_, _09792_);
  and (_11775_, _11774_, _11772_);
  or (_11777_, _11775_, _11771_);
  or (_11779_, _11777_, _09791_);
  or (_11780_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_11781_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  and (_11782_, _11781_, _05549_);
  and (_11783_, _11782_, _11780_);
  or (_11784_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_11785_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  and (_11786_, _11785_, _09792_);
  and (_11787_, _11786_, _11784_);
  or (_11788_, _11787_, _11783_);
  or (_11789_, _11788_, _05535_);
  and (_11790_, _11789_, _05542_);
  and (_11791_, _11790_, _11779_);
  or (_11793_, _11791_, _11767_);
  and (_11794_, _11793_, _09850_);
  and (_11796_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  and (_11797_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  or (_11798_, _11797_, _11796_);
  and (_11799_, _11798_, _09792_);
  and (_11800_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  and (_11801_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_11802_, _11801_, _11800_);
  and (_11803_, _11802_, _05549_);
  or (_11804_, _11803_, _11799_);
  or (_11805_, _11804_, _09791_);
  and (_11806_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  and (_11807_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_11808_, _11807_, _11806_);
  and (_11809_, _11808_, _09792_);
  and (_11810_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  and (_11811_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_11812_, _11811_, _11810_);
  and (_11813_, _11812_, _05549_);
  or (_11814_, _11813_, _11809_);
  or (_11815_, _11814_, _05535_);
  and (_11816_, _11815_, _09805_);
  and (_11817_, _11816_, _11805_);
  or (_11818_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_11819_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  and (_11820_, _11819_, _11818_);
  and (_11821_, _11820_, _09792_);
  or (_11822_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_11823_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  and (_11824_, _11823_, _11822_);
  and (_11825_, _11824_, _05549_);
  or (_11826_, _11825_, _11821_);
  or (_11827_, _11826_, _09791_);
  or (_11828_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_11829_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  and (_11830_, _11829_, _11828_);
  and (_11831_, _11830_, _09792_);
  or (_11832_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_11833_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  and (_11834_, _11833_, _11832_);
  and (_11835_, _11834_, _05549_);
  or (_11836_, _11835_, _11831_);
  or (_11837_, _11836_, _05535_);
  and (_11838_, _11837_, _05542_);
  and (_11839_, _11838_, _11827_);
  or (_11840_, _11839_, _11817_);
  and (_11841_, _11840_, _05518_);
  or (_11842_, _11841_, _11794_);
  and (_11843_, _11842_, _09790_);
  or (_11844_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_11845_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  and (_11846_, _11845_, _11844_);
  and (_11847_, _11846_, _09792_);
  or (_11848_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_11849_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  and (_11850_, _11849_, _11848_);
  and (_11851_, _11850_, _05549_);
  or (_11852_, _11851_, _11847_);
  and (_11853_, _11852_, _09791_);
  or (_11854_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_11855_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  and (_11856_, _11855_, _11854_);
  and (_11857_, _11856_, _09792_);
  or (_11858_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_11859_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  and (_11860_, _11859_, _11858_);
  and (_11861_, _11860_, _05549_);
  or (_11862_, _11861_, _11857_);
  and (_11863_, _11862_, _05535_);
  or (_11864_, _11863_, _11853_);
  and (_11865_, _11864_, _05542_);
  and (_11866_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  and (_11867_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_11868_, _11867_, _11866_);
  and (_11869_, _11868_, _09792_);
  and (_11870_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  and (_11871_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  or (_11872_, _11871_, _11870_);
  and (_11873_, _11872_, _05549_);
  or (_11874_, _11873_, _11869_);
  and (_11875_, _11874_, _09791_);
  and (_11876_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  and (_11877_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  or (_11878_, _11877_, _11876_);
  and (_11879_, _11878_, _09792_);
  and (_11880_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  and (_11881_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  or (_11882_, _11881_, _11880_);
  and (_11883_, _11882_, _05549_);
  or (_11884_, _11883_, _11879_);
  and (_11885_, _11884_, _05535_);
  or (_11886_, _11885_, _11875_);
  and (_11887_, _11886_, _09805_);
  or (_11888_, _11887_, _11865_);
  and (_11889_, _11888_, _05518_);
  or (_11890_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or (_11892_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  and (_11893_, _11892_, _05549_);
  and (_11894_, _11893_, _11890_);
  or (_11895_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_11896_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  and (_11897_, _11896_, _09792_);
  and (_11898_, _11897_, _11895_);
  or (_11899_, _11898_, _11894_);
  and (_11900_, _11899_, _09791_);
  or (_11901_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  or (_11903_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  and (_11904_, _11903_, _05549_);
  and (_11905_, _11904_, _11901_);
  or (_11907_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  or (_11908_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  and (_11910_, _11908_, _09792_);
  and (_11911_, _11910_, _11907_);
  or (_11912_, _11911_, _11905_);
  and (_11913_, _11912_, _05535_);
  or (_11915_, _11913_, _11900_);
  and (_11917_, _11915_, _05542_);
  and (_11918_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  and (_11919_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_11921_, _11919_, _11918_);
  and (_11922_, _11921_, _09792_);
  and (_11923_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  and (_11924_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_11926_, _11924_, _11923_);
  and (_11928_, _11926_, _05549_);
  or (_11929_, _11928_, _11922_);
  and (_11930_, _11929_, _09791_);
  and (_11931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  and (_11933_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_11935_, _11933_, _11931_);
  and (_11936_, _11935_, _09792_);
  and (_11938_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  and (_11939_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_11940_, _11939_, _11938_);
  and (_11941_, _11940_, _05549_);
  or (_11942_, _11941_, _11936_);
  and (_11943_, _11942_, _05535_);
  or (_11944_, _11943_, _11930_);
  and (_11945_, _11944_, _09805_);
  or (_11946_, _11945_, _11917_);
  and (_11947_, _11946_, _09850_);
  or (_11948_, _11947_, _11889_);
  and (_11949_, _11948_, _05520_);
  or (_11950_, _11949_, _11843_);
  or (_11951_, _11950_, _10033_);
  and (_11952_, _11951_, _11733_);
  or (_11953_, _11952_, _00143_);
  and (_11954_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  and (_11955_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  or (_11956_, _11955_, _11954_);
  and (_11957_, _11956_, _09792_);
  and (_11958_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  and (_11959_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  or (_11960_, _11959_, _11958_);
  and (_11961_, _11960_, _05549_);
  or (_11962_, _11961_, _11957_);
  or (_11963_, _11962_, _09791_);
  and (_11964_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  and (_11965_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  or (_11966_, _11965_, _11964_);
  and (_11967_, _11966_, _09792_);
  and (_11968_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  and (_11969_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  or (_11970_, _11969_, _11968_);
  and (_11971_, _11970_, _05549_);
  or (_11972_, _11971_, _11967_);
  or (_11974_, _11972_, _05535_);
  and (_11975_, _11974_, _09805_);
  and (_11976_, _11975_, _11963_);
  or (_11977_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  or (_11978_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  and (_11979_, _11978_, _11977_);
  and (_11980_, _11979_, _09792_);
  or (_11981_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  or (_11982_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  and (_11983_, _11982_, _11981_);
  and (_11984_, _11983_, _05549_);
  or (_11985_, _11984_, _11980_);
  or (_11986_, _11985_, _09791_);
  or (_11987_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  or (_11988_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  and (_11989_, _11988_, _11987_);
  and (_11990_, _11989_, _09792_);
  or (_11991_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_11992_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  and (_11993_, _11992_, _11991_);
  and (_11995_, _11993_, _05549_);
  or (_11996_, _11995_, _11990_);
  or (_11997_, _11996_, _05535_);
  and (_11998_, _11997_, _05542_);
  and (_11999_, _11998_, _11986_);
  or (_12000_, _11999_, _11976_);
  and (_12001_, _12000_, _05518_);
  and (_12002_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_12003_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  or (_12004_, _12003_, _12002_);
  and (_12005_, _12004_, _09792_);
  and (_12006_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  and (_12007_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  or (_12008_, _12007_, _12006_);
  and (_12009_, _12008_, _05549_);
  or (_12010_, _12009_, _12005_);
  or (_12011_, _12010_, _09791_);
  and (_12012_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  and (_12013_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  or (_12014_, _12013_, _12012_);
  and (_12015_, _12014_, _09792_);
  and (_12016_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  and (_12017_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  or (_12018_, _12017_, _12016_);
  and (_12019_, _12018_, _05549_);
  or (_12020_, _12019_, _12015_);
  or (_12021_, _12020_, _05535_);
  and (_12022_, _12021_, _09805_);
  and (_12023_, _12022_, _12011_);
  or (_12024_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  or (_12025_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  and (_12026_, _12025_, _05549_);
  and (_12027_, _12026_, _12024_);
  or (_12028_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  or (_12029_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_12030_, _12029_, _09792_);
  and (_12031_, _12030_, _12028_);
  or (_12032_, _12031_, _12027_);
  or (_12033_, _12032_, _09791_);
  or (_12034_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  or (_12035_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  and (_12036_, _12035_, _05549_);
  and (_12037_, _12036_, _12034_);
  or (_12038_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  or (_12039_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_12040_, _12039_, _09792_);
  and (_12041_, _12040_, _12038_);
  or (_12042_, _12041_, _12037_);
  or (_12043_, _12042_, _05535_);
  and (_12044_, _12043_, _05542_);
  and (_12045_, _12044_, _12033_);
  or (_12046_, _12045_, _12023_);
  and (_12047_, _12046_, _09850_);
  or (_12048_, _12047_, _12001_);
  and (_12049_, _12048_, _09790_);
  and (_12050_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  and (_12051_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or (_12052_, _12051_, _12050_);
  and (_12053_, _12052_, _09792_);
  and (_12054_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  and (_12055_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_12056_, _12055_, _12054_);
  and (_12057_, _12056_, _05549_);
  or (_12058_, _12057_, _12053_);
  and (_12059_, _12058_, _05535_);
  and (_12060_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  and (_12061_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or (_12062_, _12061_, _12060_);
  and (_12063_, _12062_, _09792_);
  and (_12064_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  and (_12066_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  or (_12067_, _12066_, _12064_);
  and (_12068_, _12067_, _05549_);
  or (_12069_, _12068_, _12063_);
  and (_12070_, _12069_, _09791_);
  or (_12071_, _12070_, _12059_);
  and (_12072_, _12071_, _09805_);
  or (_12073_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_12074_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  and (_12075_, _12074_, _05549_);
  and (_12076_, _12075_, _12073_);
  or (_12077_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_12078_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  and (_12079_, _12078_, _09792_);
  and (_12080_, _12079_, _12077_);
  or (_12081_, _12080_, _12076_);
  and (_12082_, _12081_, _05535_);
  or (_12083_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_12084_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  and (_12085_, _12084_, _05549_);
  and (_12086_, _12085_, _12083_);
  or (_12087_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or (_12088_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  and (_12089_, _12088_, _09792_);
  and (_12090_, _12089_, _12087_);
  or (_12091_, _12090_, _12086_);
  and (_12093_, _12091_, _09791_);
  or (_12094_, _12093_, _12082_);
  and (_12095_, _12094_, _05542_);
  or (_12096_, _12095_, _12072_);
  and (_12097_, _12096_, _09850_);
  and (_12098_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  and (_12099_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or (_12100_, _12099_, _12098_);
  and (_12101_, _12100_, _09792_);
  and (_12102_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  and (_12103_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or (_12104_, _12103_, _12102_);
  and (_12105_, _12104_, _05549_);
  or (_12106_, _12105_, _12101_);
  and (_12107_, _12106_, _05535_);
  and (_12108_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  and (_12109_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or (_12110_, _12109_, _12108_);
  and (_12111_, _12110_, _09792_);
  and (_12112_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  and (_12113_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_12114_, _12113_, _12112_);
  and (_12115_, _12114_, _05549_);
  or (_12116_, _12115_, _12111_);
  and (_12117_, _12116_, _09791_);
  or (_12118_, _12117_, _12107_);
  and (_12119_, _12118_, _09805_);
  or (_12120_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_12121_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  and (_12122_, _12121_, _12120_);
  and (_12123_, _12122_, _09792_);
  or (_12124_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or (_12125_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  and (_12126_, _12125_, _12124_);
  and (_12127_, _12126_, _05549_);
  or (_12128_, _12127_, _12123_);
  and (_12129_, _12128_, _05535_);
  or (_12130_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or (_12131_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  and (_12132_, _12131_, _12130_);
  and (_12133_, _12132_, _09792_);
  or (_12134_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or (_12135_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  and (_12136_, _12135_, _12134_);
  and (_12137_, _12136_, _05549_);
  or (_12138_, _12137_, _12133_);
  and (_12139_, _12138_, _09791_);
  or (_12141_, _12139_, _12129_);
  and (_12143_, _12141_, _05542_);
  or (_12144_, _12143_, _12119_);
  and (_12145_, _12144_, _05518_);
  or (_12146_, _12145_, _12097_);
  and (_12147_, _12146_, _05520_);
  or (_12149_, _12147_, _12049_);
  or (_12150_, _12149_, _05526_);
  and (_12151_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  and (_12152_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  or (_12153_, _12152_, _12151_);
  and (_12155_, _12153_, _09792_);
  and (_12156_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  and (_12157_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_12158_, _12157_, _12156_);
  and (_12159_, _12158_, _05549_);
  or (_12160_, _12159_, _12155_);
  or (_12161_, _12160_, _09791_);
  and (_12162_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  and (_12163_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  or (_12164_, _12163_, _12162_);
  and (_12165_, _12164_, _09792_);
  and (_12166_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  and (_12167_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  or (_12168_, _12167_, _12166_);
  and (_12169_, _12168_, _05549_);
  or (_12170_, _12169_, _12165_);
  or (_12171_, _12170_, _05535_);
  and (_12172_, _12171_, _09805_);
  and (_12173_, _12172_, _12161_);
  or (_12174_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  or (_12175_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  and (_12176_, _12175_, _05549_);
  and (_12177_, _12176_, _12174_);
  or (_12178_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  or (_12179_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  and (_12180_, _12179_, _09792_);
  and (_12181_, _12180_, _12178_);
  or (_12182_, _12181_, _12177_);
  or (_12183_, _12182_, _09791_);
  or (_12184_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  or (_12185_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  and (_12186_, _12185_, _05549_);
  and (_12187_, _12186_, _12184_);
  or (_12188_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  or (_12189_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  and (_12190_, _12189_, _09792_);
  and (_12191_, _12190_, _12188_);
  or (_12192_, _12191_, _12187_);
  or (_12193_, _12192_, _05535_);
  and (_12194_, _12193_, _05542_);
  and (_12195_, _12194_, _12183_);
  or (_12196_, _12195_, _12173_);
  and (_12197_, _12196_, _09850_);
  and (_12198_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  and (_12199_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  or (_12200_, _12199_, _12198_);
  and (_12201_, _12200_, _09792_);
  and (_12203_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  and (_12204_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  or (_12205_, _12204_, _12203_);
  and (_12206_, _12205_, _05549_);
  or (_12207_, _12206_, _12201_);
  or (_12208_, _12207_, _09791_);
  and (_12209_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  and (_12210_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or (_12211_, _12210_, _12209_);
  and (_12212_, _12211_, _09792_);
  and (_12213_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  and (_12214_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_12215_, _12214_, _12213_);
  and (_12216_, _12215_, _05549_);
  or (_12217_, _12216_, _12212_);
  or (_12218_, _12217_, _05535_);
  and (_12219_, _12218_, _09805_);
  and (_12220_, _12219_, _12208_);
  or (_12221_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_12222_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  and (_12223_, _12222_, _12221_);
  and (_12225_, _12223_, _09792_);
  or (_12226_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  or (_12227_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  and (_12228_, _12227_, _12226_);
  and (_12229_, _12228_, _05549_);
  or (_12230_, _12229_, _12225_);
  or (_12231_, _12230_, _09791_);
  or (_12232_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  or (_12233_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  and (_12234_, _12233_, _12232_);
  and (_12235_, _12234_, _09792_);
  or (_12236_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_12237_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  and (_12238_, _12237_, _12236_);
  and (_12239_, _12238_, _05549_);
  or (_12240_, _12239_, _12235_);
  or (_12241_, _12240_, _05535_);
  and (_12242_, _12241_, _05542_);
  and (_12244_, _12242_, _12231_);
  or (_12245_, _12244_, _12220_);
  and (_12246_, _12245_, _05518_);
  or (_12247_, _12246_, _12197_);
  and (_12248_, _12247_, _09790_);
  or (_12249_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  or (_12250_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  and (_12252_, _12250_, _12249_);
  and (_12253_, _12252_, _09792_);
  or (_12254_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  or (_12255_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  and (_12256_, _12255_, _12254_);
  and (_12257_, _12256_, _05549_);
  or (_12258_, _12257_, _12253_);
  and (_12259_, _12258_, _09791_);
  or (_12260_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  or (_12262_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  and (_12263_, _12262_, _12260_);
  and (_12264_, _12263_, _09792_);
  or (_12265_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  or (_12267_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  and (_12269_, _12267_, _12265_);
  and (_12270_, _12269_, _05549_);
  or (_12271_, _12270_, _12264_);
  and (_12272_, _12271_, _05535_);
  or (_12273_, _12272_, _12259_);
  and (_12275_, _12273_, _05542_);
  and (_12276_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and (_12277_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  or (_12278_, _12277_, _12276_);
  and (_12279_, _12278_, _09792_);
  and (_12281_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  and (_12282_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  or (_12283_, _12282_, _12281_);
  and (_12284_, _12283_, _05549_);
  or (_12285_, _12284_, _12279_);
  and (_12286_, _12285_, _09791_);
  and (_12287_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  and (_12288_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  or (_12289_, _12288_, _12287_);
  and (_12290_, _12289_, _09792_);
  and (_12291_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  and (_12292_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  or (_12294_, _12292_, _12291_);
  and (_12295_, _12294_, _05549_);
  or (_12296_, _12295_, _12290_);
  and (_12297_, _12296_, _05535_);
  or (_12298_, _12297_, _12286_);
  and (_12299_, _12298_, _09805_);
  or (_12300_, _12299_, _12275_);
  and (_12302_, _12300_, _05518_);
  or (_12303_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or (_12304_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  and (_12305_, _12304_, _05549_);
  and (_12306_, _12305_, _12303_);
  or (_12307_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  or (_12308_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  and (_12309_, _12308_, _09792_);
  and (_12310_, _12309_, _12307_);
  or (_12311_, _12310_, _12306_);
  and (_12312_, _12311_, _09791_);
  or (_12313_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  or (_12314_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  and (_12315_, _12314_, _05549_);
  and (_12317_, _12315_, _12313_);
  or (_12318_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  or (_12319_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  and (_12320_, _12319_, _09792_);
  and (_12321_, _12320_, _12318_);
  or (_12322_, _12321_, _12317_);
  and (_12323_, _12322_, _05535_);
  or (_12324_, _12323_, _12312_);
  and (_12326_, _12324_, _05542_);
  and (_12327_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  and (_12328_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  or (_12329_, _12328_, _12327_);
  and (_12330_, _12329_, _09792_);
  and (_12331_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  and (_12333_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or (_12335_, _12333_, _12331_);
  and (_12336_, _12335_, _05549_);
  or (_12337_, _12336_, _12330_);
  and (_12338_, _12337_, _09791_);
  and (_12339_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  and (_12341_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  or (_12343_, _12341_, _12339_);
  and (_12345_, _12343_, _09792_);
  and (_12346_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  and (_12347_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or (_12349_, _12347_, _12346_);
  and (_12350_, _12349_, _05549_);
  or (_12352_, _12350_, _12345_);
  and (_12354_, _12352_, _05535_);
  or (_12356_, _12354_, _12338_);
  and (_12358_, _12356_, _09805_);
  or (_12359_, _12358_, _12326_);
  and (_12360_, _12359_, _09850_);
  or (_12361_, _12360_, _12302_);
  and (_12362_, _12361_, _05520_);
  or (_12363_, _12362_, _12248_);
  or (_12364_, _12363_, _10033_);
  and (_12365_, _12364_, _12150_);
  or (_12366_, _12365_, _04413_);
  and (_12367_, _12366_, _11953_);
  or (_12368_, _12367_, _05563_);
  or (_12370_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_12371_, _12370_, _22731_);
  and (_04460_, _12371_, _12368_);
  and (_12372_, _09779_, _23941_);
  and (_12373_, _12372_, _23887_);
  not (_12374_, _12372_);
  and (_12375_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  or (_04471_, _12375_, _12373_);
  and (_12376_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  and (_12377_, _02513_, _23583_);
  or (_04473_, _12377_, _12376_);
  and (_12378_, _10746_, _23548_);
  and (_12379_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  or (_04487_, _12379_, _12378_);
  and (_12380_, _06763_, _24089_);
  and (_12381_, _06765_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_04490_, _12381_, _12380_);
  and (_12382_, _12372_, _23548_);
  and (_12383_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  or (_04492_, _12383_, _12382_);
  and (_12385_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  and (_12386_, _02513_, _24134_);
  or (_27089_, _12386_, _12385_);
  and (_12388_, _07038_, _23548_);
  and (_12389_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_04504_, _12389_, _12388_);
  and (_12392_, _07038_, _23583_);
  and (_12394_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_04506_, _12394_, _12392_);
  and (_12395_, _05438_, _24089_);
  and (_12396_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_04509_, _12396_, _12395_);
  and (_12398_, _05438_, _24134_);
  and (_12400_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  or (_04511_, _12400_, _12398_);
  and (_12401_, _07013_, _24051_);
  and (_12402_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  or (_04515_, _12402_, _12401_);
  and (_12403_, _07038_, _23887_);
  and (_12405_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_04525_, _12405_, _12403_);
  and (_12406_, _05438_, _24051_);
  and (_12407_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  or (_04546_, _12407_, _12406_);
  and (_12408_, _24409_, _24089_);
  and (_12409_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  or (_04562_, _12409_, _12408_);
  and (_12410_, _12372_, _23583_);
  and (_12411_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  or (_26996_, _12411_, _12410_);
  and (_12414_, _12372_, _24051_);
  and (_12415_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  or (_04571_, _12415_, _12414_);
  and (_12418_, _12372_, _24089_);
  and (_12419_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  or (_04576_, _12419_, _12418_);
  and (_12421_, _05442_, _24051_);
  and (_12423_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  or (_04588_, _12423_, _12421_);
  and (_12425_, _05442_, _23996_);
  and (_12426_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_04591_, _12426_, _12425_);
  and (_12427_, _07013_, _23996_);
  and (_12428_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_04600_, _12428_, _12427_);
  and (_12429_, _24476_, _23941_);
  and (_12430_, _12429_, _23996_);
  not (_12431_, _12429_);
  and (_12433_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  or (_04618_, _12433_, _12430_);
  and (_12434_, _24510_, _23887_);
  and (_12435_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_04621_, _12435_, _12434_);
  and (_12436_, _24510_, _23548_);
  and (_12437_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_04624_, _12437_, _12436_);
  and (_12438_, _24476_, _24297_);
  and (_12439_, _12438_, _23887_);
  not (_12440_, _12438_);
  and (_12441_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  or (_04655_, _12441_, _12439_);
  and (_12442_, _09779_, _24899_);
  and (_12443_, _12442_, _24089_);
  not (_12444_, _12442_);
  and (_12445_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  or (_04664_, _12445_, _12443_);
  and (_12446_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  and (_12447_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_12448_, _12447_, _12446_);
  and (_12449_, _12448_, _09792_);
  and (_12450_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  and (_12451_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  or (_12452_, _12451_, _12450_);
  and (_12453_, _12452_, _05549_);
  or (_12454_, _12453_, _12449_);
  or (_12455_, _12454_, _09791_);
  and (_12456_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  and (_12457_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_12458_, _12457_, _12456_);
  and (_12459_, _12458_, _09792_);
  and (_12460_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  and (_12461_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_12462_, _12461_, _12460_);
  and (_12463_, _12462_, _05549_);
  or (_12464_, _12463_, _12459_);
  or (_12465_, _12464_, _05535_);
  and (_12466_, _12465_, _09805_);
  and (_12467_, _12466_, _12455_);
  or (_12468_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_12469_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  and (_12470_, _12469_, _12468_);
  and (_12471_, _12470_, _09792_);
  or (_12472_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  or (_12473_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  and (_12474_, _12473_, _12472_);
  and (_12475_, _12474_, _05549_);
  or (_12476_, _12475_, _12471_);
  or (_12477_, _12476_, _09791_);
  or (_12478_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_12479_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  and (_12480_, _12479_, _12478_);
  and (_12481_, _12480_, _09792_);
  or (_12482_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  or (_12483_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  and (_12484_, _12483_, _12482_);
  and (_12485_, _12484_, _05549_);
  or (_12486_, _12485_, _12481_);
  or (_12487_, _12486_, _05535_);
  and (_12488_, _12487_, _05542_);
  and (_12489_, _12488_, _12477_);
  or (_12490_, _12489_, _12467_);
  and (_12491_, _12490_, _05518_);
  and (_12492_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  and (_12493_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  or (_12494_, _12493_, _12492_);
  and (_12495_, _12494_, _09792_);
  and (_12496_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  and (_12497_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_12498_, _12497_, _12496_);
  and (_12499_, _12498_, _05549_);
  or (_12500_, _12499_, _12495_);
  or (_12501_, _12500_, _09791_);
  and (_12502_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  and (_12503_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  or (_12504_, _12503_, _12502_);
  and (_12505_, _12504_, _09792_);
  and (_12506_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  and (_12507_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_12508_, _12507_, _12506_);
  and (_12509_, _12508_, _05549_);
  or (_12510_, _12509_, _12505_);
  or (_12511_, _12510_, _05535_);
  and (_12512_, _12511_, _09805_);
  and (_12513_, _12512_, _12501_);
  or (_12514_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  or (_12516_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  and (_12517_, _12516_, _05549_);
  and (_12518_, _12517_, _12514_);
  or (_12519_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  or (_12520_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  and (_12521_, _12520_, _09792_);
  and (_12522_, _12521_, _12519_);
  or (_12523_, _12522_, _12518_);
  or (_12524_, _12523_, _09791_);
  or (_12525_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_12526_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  and (_12527_, _12526_, _05549_);
  and (_12528_, _12527_, _12525_);
  or (_12529_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  or (_12530_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  and (_12531_, _12530_, _09792_);
  and (_12532_, _12531_, _12529_);
  or (_12533_, _12532_, _12528_);
  or (_12534_, _12533_, _05535_);
  and (_12535_, _12534_, _05542_);
  and (_12536_, _12535_, _12524_);
  or (_12537_, _12536_, _12513_);
  and (_12538_, _12537_, _09850_);
  or (_12539_, _12538_, _12491_);
  and (_12540_, _12539_, _09790_);
  and (_12541_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_12542_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or (_12543_, _12542_, _12541_);
  and (_12544_, _12543_, _09792_);
  and (_12545_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_12546_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_12547_, _12546_, _12545_);
  and (_12548_, _12547_, _05549_);
  or (_12549_, _12548_, _12544_);
  and (_12550_, _12549_, _05535_);
  and (_12551_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_12552_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_12553_, _12552_, _12551_);
  and (_12554_, _12553_, _09792_);
  and (_12555_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_12556_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_12557_, _12556_, _12555_);
  and (_12558_, _12557_, _05549_);
  or (_12559_, _12558_, _12554_);
  and (_12560_, _12559_, _09791_);
  or (_12561_, _12560_, _12550_);
  and (_12562_, _12561_, _09805_);
  or (_12563_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_12564_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and (_12565_, _12564_, _05549_);
  and (_12566_, _12565_, _12563_);
  or (_12567_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_12568_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  and (_12569_, _12568_, _09792_);
  and (_12570_, _12569_, _12567_);
  or (_12571_, _12570_, _12566_);
  and (_12572_, _12571_, _05535_);
  or (_12573_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_12574_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_12575_, _12574_, _05549_);
  and (_12576_, _12575_, _12573_);
  or (_12577_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_12578_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  and (_12579_, _12578_, _09792_);
  and (_12580_, _12579_, _12577_);
  or (_12581_, _12580_, _12576_);
  and (_12582_, _12581_, _09791_);
  or (_12583_, _12582_, _12572_);
  and (_12584_, _12583_, _05542_);
  or (_12585_, _12584_, _12562_);
  and (_12586_, _12585_, _09850_);
  and (_12587_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  and (_12588_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  or (_12589_, _12588_, _12587_);
  and (_12590_, _12589_, _09792_);
  and (_12591_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  and (_12592_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_12593_, _12592_, _12591_);
  and (_12594_, _12593_, _05549_);
  or (_12595_, _12594_, _12590_);
  and (_12596_, _12595_, _05535_);
  and (_12597_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  and (_12598_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_12599_, _12598_, _12597_);
  and (_12600_, _12599_, _09792_);
  and (_12601_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  and (_12602_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  or (_12603_, _12602_, _12601_);
  and (_12604_, _12603_, _05549_);
  or (_12605_, _12604_, _12600_);
  and (_12606_, _12605_, _09791_);
  or (_12607_, _12606_, _12596_);
  and (_12608_, _12607_, _09805_);
  or (_12609_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  or (_12610_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  and (_12611_, _12610_, _12609_);
  and (_12612_, _12611_, _09792_);
  or (_12613_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  or (_12614_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  and (_12615_, _12614_, _12613_);
  and (_12617_, _12615_, _05549_);
  or (_12618_, _12617_, _12612_);
  and (_12619_, _12618_, _05535_);
  or (_12620_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  or (_12621_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  and (_12622_, _12621_, _12620_);
  and (_12623_, _12622_, _09792_);
  or (_12624_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  or (_12625_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  and (_12626_, _12625_, _12624_);
  and (_12627_, _12626_, _05549_);
  or (_12628_, _12627_, _12623_);
  and (_12629_, _12628_, _09791_);
  or (_12630_, _12629_, _12619_);
  and (_12631_, _12630_, _05542_);
  or (_12632_, _12631_, _12608_);
  and (_12633_, _12632_, _05518_);
  or (_12634_, _12633_, _12586_);
  and (_12635_, _12634_, _05520_);
  or (_12636_, _12635_, _12540_);
  or (_12638_, _12636_, _05526_);
  and (_12639_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  and (_12640_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_12641_, _12640_, _12639_);
  and (_12642_, _12641_, _09792_);
  and (_12643_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  and (_12644_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_12645_, _12644_, _12643_);
  and (_12646_, _12645_, _05549_);
  or (_12647_, _12646_, _12642_);
  or (_12648_, _12647_, _09791_);
  and (_12649_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  and (_12650_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_12651_, _12650_, _12649_);
  and (_12652_, _12651_, _09792_);
  and (_12653_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  and (_12654_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_12655_, _12654_, _12653_);
  and (_12656_, _12655_, _05549_);
  or (_12657_, _12656_, _12652_);
  or (_12658_, _12657_, _05535_);
  and (_12659_, _12658_, _09805_);
  and (_12660_, _12659_, _12648_);
  or (_12661_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_12662_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  and (_12663_, _12662_, _05549_);
  and (_12664_, _12663_, _12661_);
  or (_12665_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_12666_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  and (_12667_, _12666_, _09792_);
  and (_12668_, _12667_, _12665_);
  or (_12669_, _12668_, _12664_);
  or (_12670_, _12669_, _09791_);
  or (_12671_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_12672_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  and (_12673_, _12672_, _05549_);
  and (_12674_, _12673_, _12671_);
  or (_12675_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_12676_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  and (_12677_, _12676_, _09792_);
  and (_12678_, _12677_, _12675_);
  or (_12679_, _12678_, _12674_);
  or (_12680_, _12679_, _05535_);
  and (_12681_, _12680_, _05542_);
  and (_12682_, _12681_, _12670_);
  or (_12683_, _12682_, _12660_);
  and (_12684_, _12683_, _09850_);
  and (_12685_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  and (_12686_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  or (_12687_, _12686_, _12685_);
  and (_12688_, _12687_, _09792_);
  and (_12689_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  and (_12690_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_12691_, _12690_, _12689_);
  and (_12692_, _12691_, _05549_);
  or (_12693_, _12692_, _12688_);
  or (_12694_, _12693_, _09791_);
  and (_12695_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  and (_12696_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_12697_, _12696_, _12695_);
  and (_12698_, _12697_, _09792_);
  and (_12699_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  and (_12700_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_12701_, _12700_, _12699_);
  and (_12702_, _12701_, _05549_);
  or (_12703_, _12702_, _12698_);
  or (_12704_, _12703_, _05535_);
  and (_12705_, _12704_, _09805_);
  and (_12706_, _12705_, _12694_);
  or (_12707_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_12708_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  and (_12709_, _12708_, _12707_);
  and (_12710_, _12709_, _09792_);
  or (_12711_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_12712_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  and (_12713_, _12712_, _12711_);
  and (_12714_, _12713_, _05549_);
  or (_12715_, _12714_, _12710_);
  or (_12716_, _12715_, _09791_);
  or (_12717_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_12718_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  and (_12719_, _12718_, _12717_);
  and (_12720_, _12719_, _09792_);
  or (_12721_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  or (_12722_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  and (_12723_, _12722_, _12721_);
  and (_12724_, _12723_, _05549_);
  or (_12725_, _12724_, _12720_);
  or (_12726_, _12725_, _05535_);
  and (_12727_, _12726_, _05542_);
  and (_12728_, _12727_, _12716_);
  or (_12729_, _12728_, _12706_);
  and (_12730_, _12729_, _05518_);
  or (_12731_, _12730_, _12684_);
  and (_12732_, _12731_, _09790_);
  or (_12733_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_12734_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  and (_12735_, _12734_, _12733_);
  and (_12736_, _12735_, _09792_);
  or (_12737_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_12738_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  and (_12739_, _12738_, _12737_);
  and (_12740_, _12739_, _05549_);
  or (_12741_, _12740_, _12736_);
  and (_12742_, _12741_, _09791_);
  or (_12743_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_12744_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  and (_12745_, _12744_, _12743_);
  and (_12746_, _12745_, _09792_);
  or (_12747_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_12749_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  and (_12750_, _12749_, _12747_);
  and (_12751_, _12750_, _05549_);
  or (_12752_, _12751_, _12746_);
  and (_12753_, _12752_, _05535_);
  or (_12754_, _12753_, _12742_);
  and (_12755_, _12754_, _05542_);
  and (_12756_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  and (_12757_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_12758_, _12757_, _12756_);
  and (_12759_, _12758_, _09792_);
  and (_12760_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  and (_12761_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  or (_12762_, _12761_, _12760_);
  and (_12763_, _12762_, _05549_);
  or (_12764_, _12763_, _12759_);
  and (_12765_, _12764_, _09791_);
  and (_12766_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  and (_12767_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_12768_, _12767_, _12766_);
  and (_12769_, _12768_, _09792_);
  and (_12770_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  and (_12771_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  or (_12772_, _12771_, _12770_);
  and (_12773_, _12772_, _05549_);
  or (_12774_, _12773_, _12769_);
  and (_12775_, _12774_, _05535_);
  or (_12776_, _12775_, _12765_);
  and (_12777_, _12776_, _09805_);
  or (_12778_, _12777_, _12755_);
  and (_12779_, _12778_, _05518_);
  or (_12780_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or (_12781_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  and (_12782_, _12781_, _05549_);
  and (_12783_, _12782_, _12780_);
  or (_12784_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or (_12785_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  and (_12786_, _12785_, _09792_);
  and (_12787_, _12786_, _12784_);
  or (_12788_, _12787_, _12783_);
  and (_12789_, _12788_, _09791_);
  or (_12790_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or (_12791_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  and (_12792_, _12791_, _05549_);
  and (_12793_, _12792_, _12790_);
  or (_12794_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or (_12795_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  and (_12796_, _12795_, _09792_);
  and (_12797_, _12796_, _12794_);
  or (_12798_, _12797_, _12793_);
  and (_12799_, _12798_, _05535_);
  or (_12800_, _12799_, _12789_);
  and (_12801_, _12800_, _05542_);
  and (_12802_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  and (_12803_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or (_12804_, _12803_, _12802_);
  and (_12805_, _12804_, _09792_);
  and (_12806_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  and (_12807_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or (_12808_, _12807_, _12806_);
  and (_12809_, _12808_, _05549_);
  or (_12810_, _12809_, _12805_);
  and (_12811_, _12810_, _09791_);
  and (_12812_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  and (_12813_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or (_12814_, _12813_, _12812_);
  and (_12815_, _12814_, _09792_);
  and (_12816_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  and (_12817_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or (_12818_, _12817_, _12816_);
  and (_12819_, _12818_, _05549_);
  or (_12820_, _12819_, _12815_);
  and (_12821_, _12820_, _05535_);
  or (_12822_, _12821_, _12811_);
  and (_12823_, _12822_, _09805_);
  or (_12824_, _12823_, _12801_);
  and (_12825_, _12824_, _09850_);
  or (_12826_, _12825_, _12779_);
  and (_12827_, _12826_, _05520_);
  or (_12828_, _12827_, _12732_);
  or (_12829_, _12828_, _10033_);
  and (_12830_, _12829_, _12638_);
  or (_12831_, _12830_, _00143_);
  and (_12832_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  and (_12833_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  or (_12834_, _12833_, _12832_);
  and (_12835_, _12834_, _09792_);
  and (_12836_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  and (_12837_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  or (_12838_, _12837_, _12836_);
  and (_12839_, _12838_, _05549_);
  or (_12840_, _12839_, _12835_);
  or (_12841_, _12840_, _09791_);
  and (_12842_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  and (_12843_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  or (_12844_, _12843_, _12842_);
  and (_12845_, _12844_, _09792_);
  and (_12846_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  and (_12847_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  or (_12848_, _12847_, _12846_);
  and (_12849_, _12848_, _05549_);
  or (_12850_, _12849_, _12845_);
  or (_12851_, _12850_, _05535_);
  and (_12852_, _12851_, _09805_);
  and (_12853_, _12852_, _12841_);
  or (_12854_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  or (_12855_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  and (_12856_, _12855_, _12854_);
  and (_12857_, _12856_, _09792_);
  or (_12858_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_12859_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  and (_12860_, _12859_, _12858_);
  and (_12861_, _12860_, _05549_);
  or (_12862_, _12861_, _12857_);
  or (_12863_, _12862_, _09791_);
  or (_12864_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_12865_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  and (_12866_, _12865_, _12864_);
  and (_12867_, _12866_, _09792_);
  or (_12868_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  or (_12869_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  and (_12870_, _12869_, _12868_);
  and (_12871_, _12870_, _05549_);
  or (_12872_, _12871_, _12867_);
  or (_12873_, _12872_, _05535_);
  and (_12874_, _12873_, _05542_);
  and (_12875_, _12874_, _12863_);
  or (_12876_, _12875_, _12853_);
  and (_12877_, _12876_, _05518_);
  and (_12878_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_12879_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  or (_12880_, _12879_, _12878_);
  and (_12881_, _12880_, _09792_);
  and (_12882_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  and (_12883_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  or (_12884_, _12883_, _12882_);
  and (_12885_, _12884_, _05549_);
  or (_12886_, _12885_, _12881_);
  or (_12887_, _12886_, _09791_);
  and (_12888_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  and (_12889_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  or (_12890_, _12889_, _12888_);
  and (_12891_, _12890_, _09792_);
  and (_12892_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  and (_12893_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  or (_12894_, _12893_, _12892_);
  and (_12895_, _12894_, _05549_);
  or (_12896_, _12895_, _12891_);
  or (_12897_, _12896_, _05535_);
  and (_12898_, _12897_, _09805_);
  and (_12899_, _12898_, _12887_);
  or (_12900_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  or (_12901_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  and (_12902_, _12901_, _05549_);
  and (_12903_, _12902_, _12900_);
  or (_12904_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  or (_12905_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_12906_, _12905_, _09792_);
  and (_12907_, _12906_, _12904_);
  or (_12908_, _12907_, _12903_);
  or (_12909_, _12908_, _09791_);
  or (_12910_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  or (_12911_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  and (_12912_, _12911_, _05549_);
  and (_12913_, _12912_, _12910_);
  or (_12914_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  or (_12915_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_12916_, _12915_, _09792_);
  and (_12917_, _12916_, _12914_);
  or (_12918_, _12917_, _12913_);
  or (_12919_, _12918_, _05535_);
  and (_12920_, _12919_, _05542_);
  and (_12921_, _12920_, _12909_);
  or (_12922_, _12921_, _12899_);
  and (_12923_, _12922_, _09850_);
  or (_12924_, _12923_, _12877_);
  and (_12925_, _12924_, _09790_);
  and (_12926_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  and (_12927_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or (_12928_, _12927_, _12926_);
  and (_12929_, _12928_, _09792_);
  and (_12930_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  and (_12931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or (_12932_, _12931_, _12930_);
  and (_12933_, _12932_, _05549_);
  or (_12934_, _12933_, _12929_);
  and (_12935_, _12934_, _05535_);
  and (_12936_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  and (_12937_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or (_12938_, _12937_, _12936_);
  and (_12939_, _12938_, _09792_);
  and (_12940_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  and (_12941_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or (_12942_, _12941_, _12940_);
  and (_12943_, _12942_, _05549_);
  or (_12944_, _12943_, _12939_);
  and (_12945_, _12944_, _09791_);
  or (_12946_, _12945_, _12935_);
  and (_12947_, _12946_, _09805_);
  or (_12948_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or (_12949_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  and (_12950_, _12949_, _05549_);
  and (_12951_, _12950_, _12948_);
  or (_12952_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or (_12953_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  and (_12954_, _12953_, _09792_);
  and (_12955_, _12954_, _12952_);
  or (_12956_, _12955_, _12951_);
  and (_12957_, _12956_, _05535_);
  or (_12958_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or (_12959_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  and (_12960_, _12959_, _05549_);
  and (_12961_, _12960_, _12958_);
  or (_12962_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or (_12963_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  and (_12964_, _12963_, _09792_);
  and (_12965_, _12964_, _12962_);
  or (_12966_, _12965_, _12961_);
  and (_12967_, _12966_, _09791_);
  or (_12968_, _12967_, _12957_);
  and (_12969_, _12968_, _05542_);
  or (_12970_, _12969_, _12947_);
  and (_12971_, _12970_, _09850_);
  and (_12972_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  and (_12973_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or (_12974_, _12973_, _12972_);
  and (_12975_, _12974_, _09792_);
  and (_12976_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  and (_12977_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or (_12978_, _12977_, _12976_);
  and (_12979_, _12978_, _05549_);
  or (_12980_, _12979_, _12975_);
  and (_12981_, _12980_, _05535_);
  and (_12982_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  and (_12983_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or (_12984_, _12983_, _12982_);
  and (_12985_, _12984_, _09792_);
  and (_12986_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  and (_12987_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or (_12988_, _12987_, _12986_);
  and (_12989_, _12988_, _05549_);
  or (_12990_, _12989_, _12985_);
  and (_12991_, _12990_, _09791_);
  or (_12992_, _12991_, _12981_);
  and (_12993_, _12992_, _09805_);
  or (_12994_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or (_12995_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  and (_12996_, _12995_, _12994_);
  and (_12997_, _12996_, _09792_);
  or (_12998_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  or (_12999_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  and (_13000_, _12999_, _12998_);
  and (_13001_, _13000_, _05549_);
  or (_13002_, _13001_, _12997_);
  and (_13003_, _13002_, _05535_);
  or (_13004_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  or (_13005_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  and (_13006_, _13005_, _13004_);
  and (_13007_, _13006_, _09792_);
  or (_13008_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  or (_13009_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  and (_13010_, _13009_, _13008_);
  and (_13011_, _13010_, _05549_);
  or (_13012_, _13011_, _13007_);
  and (_13013_, _13012_, _09791_);
  or (_13014_, _13013_, _13003_);
  and (_13015_, _13014_, _05542_);
  or (_13016_, _13015_, _12993_);
  and (_13017_, _13016_, _05518_);
  or (_13018_, _13017_, _12971_);
  and (_13019_, _13018_, _05520_);
  or (_13020_, _13019_, _12925_);
  or (_13021_, _13020_, _05526_);
  and (_13022_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  and (_13023_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  or (_13024_, _13023_, _13022_);
  and (_13025_, _13024_, _09792_);
  and (_13026_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  and (_13027_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_13028_, _13027_, _13026_);
  and (_13029_, _13028_, _05549_);
  or (_13030_, _13029_, _13025_);
  or (_13031_, _13030_, _09791_);
  and (_13032_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  and (_13033_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_13034_, _13033_, _13032_);
  and (_13035_, _13034_, _09792_);
  and (_13036_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  and (_13037_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  or (_13038_, _13037_, _13036_);
  and (_13039_, _13038_, _05549_);
  or (_13040_, _13039_, _13035_);
  or (_13041_, _13040_, _05535_);
  and (_13042_, _13041_, _09805_);
  and (_13043_, _13042_, _13031_);
  or (_13044_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  or (_13045_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  and (_13046_, _13045_, _05549_);
  and (_13047_, _13046_, _13044_);
  or (_13048_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_13049_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  and (_13050_, _13049_, _09792_);
  and (_13051_, _13050_, _13048_);
  or (_13052_, _13051_, _13047_);
  or (_13053_, _13052_, _09791_);
  or (_13054_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  or (_13055_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  and (_13056_, _13055_, _05549_);
  and (_13057_, _13056_, _13054_);
  or (_13058_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  or (_13059_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  and (_13060_, _13059_, _09792_);
  and (_13061_, _13060_, _13058_);
  or (_13062_, _13061_, _13057_);
  or (_13063_, _13062_, _05535_);
  and (_13064_, _13063_, _05542_);
  and (_13065_, _13064_, _13053_);
  or (_13066_, _13065_, _13043_);
  and (_13067_, _13066_, _09850_);
  and (_13068_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  and (_13069_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  or (_13070_, _13069_, _13068_);
  and (_13071_, _13070_, _09792_);
  and (_13072_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  and (_13073_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  or (_13074_, _13073_, _13072_);
  and (_13075_, _13074_, _05549_);
  or (_13076_, _13075_, _13071_);
  or (_13077_, _13076_, _09791_);
  and (_13078_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  and (_13079_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or (_13080_, _13079_, _13078_);
  and (_13081_, _13080_, _09792_);
  and (_13082_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  and (_13083_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_13084_, _13083_, _13082_);
  and (_13085_, _13084_, _05549_);
  or (_13086_, _13085_, _13081_);
  or (_13087_, _13086_, _05535_);
  and (_13088_, _13087_, _09805_);
  and (_13089_, _13088_, _13077_);
  or (_13090_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_13091_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  and (_13092_, _13091_, _13090_);
  and (_13093_, _13092_, _09792_);
  or (_13094_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_13095_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  and (_13096_, _13095_, _13094_);
  and (_13097_, _13096_, _05549_);
  or (_13098_, _13097_, _13093_);
  or (_13099_, _13098_, _09791_);
  or (_13100_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or (_13101_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  and (_13102_, _13101_, _13100_);
  and (_13103_, _13102_, _09792_);
  or (_13104_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_13105_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  and (_13106_, _13105_, _13104_);
  and (_13107_, _13106_, _05549_);
  or (_13108_, _13107_, _13103_);
  or (_13110_, _13108_, _05535_);
  and (_13111_, _13110_, _05542_);
  and (_13112_, _13111_, _13099_);
  or (_13113_, _13112_, _13089_);
  and (_13114_, _13113_, _05518_);
  or (_13115_, _13114_, _13067_);
  and (_13116_, _13115_, _09790_);
  or (_13117_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  or (_13118_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  and (_13119_, _13118_, _13117_);
  and (_13120_, _13119_, _09792_);
  or (_13121_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  or (_13122_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  and (_13123_, _13122_, _13121_);
  and (_13124_, _13123_, _05549_);
  or (_13125_, _13124_, _13120_);
  and (_13126_, _13125_, _09791_);
  or (_13127_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  or (_13128_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  and (_13129_, _13128_, _13127_);
  and (_13130_, _13129_, _09792_);
  or (_13131_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  or (_13132_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  and (_13133_, _13132_, _13131_);
  and (_13134_, _13133_, _05549_);
  or (_13135_, _13134_, _13130_);
  and (_13136_, _13135_, _05535_);
  or (_13137_, _13136_, _13126_);
  and (_13138_, _13137_, _05542_);
  and (_13139_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  and (_13140_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  or (_13141_, _13140_, _13139_);
  and (_13142_, _13141_, _09792_);
  and (_13143_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  and (_13144_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  or (_13145_, _13144_, _13143_);
  and (_13146_, _13145_, _05549_);
  or (_13147_, _13146_, _13142_);
  and (_13148_, _13147_, _09791_);
  and (_13149_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  and (_13150_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  or (_13151_, _13150_, _13149_);
  and (_13152_, _13151_, _09792_);
  and (_13153_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and (_13154_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  or (_13155_, _13154_, _13153_);
  and (_13156_, _13155_, _05549_);
  or (_13157_, _13156_, _13152_);
  and (_13158_, _13157_, _05535_);
  or (_13159_, _13158_, _13148_);
  and (_13160_, _13159_, _09805_);
  or (_13161_, _13160_, _13138_);
  and (_13162_, _13161_, _05518_);
  or (_13163_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  or (_13164_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  and (_13165_, _13164_, _05549_);
  and (_13166_, _13165_, _13163_);
  or (_13167_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  or (_13168_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  and (_13169_, _13168_, _09792_);
  and (_13170_, _13169_, _13167_);
  or (_13171_, _13170_, _13166_);
  and (_13172_, _13171_, _09791_);
  or (_13173_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  or (_13174_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  and (_13175_, _13174_, _05549_);
  and (_13176_, _13175_, _13173_);
  or (_13177_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  or (_13178_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  and (_13179_, _13178_, _09792_);
  and (_13180_, _13179_, _13177_);
  or (_13181_, _13180_, _13176_);
  and (_13182_, _13181_, _05535_);
  or (_13183_, _13182_, _13172_);
  and (_13184_, _13183_, _05542_);
  and (_13185_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  and (_13186_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_13187_, _13186_, _13185_);
  and (_13188_, _13187_, _09792_);
  and (_13189_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  and (_13190_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_13191_, _13190_, _13189_);
  and (_13192_, _13191_, _05549_);
  or (_13193_, _13192_, _13188_);
  and (_13194_, _13193_, _09791_);
  and (_13195_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  and (_13196_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  or (_13197_, _13196_, _13195_);
  and (_13198_, _13197_, _09792_);
  and (_13199_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  and (_13200_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  or (_13201_, _13200_, _13199_);
  and (_13202_, _13201_, _05549_);
  or (_13203_, _13202_, _13198_);
  and (_13204_, _13203_, _05535_);
  or (_13205_, _13204_, _13194_);
  and (_13206_, _13205_, _09805_);
  or (_13207_, _13206_, _13184_);
  and (_13208_, _13207_, _09850_);
  or (_13209_, _13208_, _13162_);
  and (_13210_, _13209_, _05520_);
  or (_13211_, _13210_, _13116_);
  or (_13212_, _13211_, _10033_);
  and (_13213_, _13212_, _13021_);
  or (_13214_, _13213_, _04413_);
  and (_13215_, _13214_, _12831_);
  or (_13216_, _13215_, _05563_);
  or (_13217_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_13218_, _13217_, _22731_);
  and (_04666_, _13218_, _13216_);
  and (_13219_, _12438_, _23548_);
  and (_13220_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  or (_27191_, _13220_, _13219_);
  and (_13221_, _12442_, _23583_);
  and (_13222_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  or (_04679_, _13222_, _13221_);
  and (_13223_, _05465_, _24089_);
  and (_13224_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  or (_27069_, _13224_, _13223_);
  and (_13225_, _12442_, _23887_);
  and (_13226_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  or (_26994_, _13226_, _13225_);
  and (_13227_, _12438_, _24134_);
  and (_13228_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  or (_04713_, _13228_, _13227_);
  and (_13229_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  and (_13230_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_13231_, _13230_, _13229_);
  and (_13232_, _13231_, _09792_);
  and (_13233_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  and (_13234_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_13235_, _13234_, _13233_);
  and (_13236_, _13235_, _05549_);
  or (_13237_, _13236_, _13232_);
  or (_13238_, _13237_, _09791_);
  and (_13239_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  and (_13240_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_13241_, _13240_, _13239_);
  and (_13242_, _13241_, _09792_);
  and (_13243_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  and (_13244_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_13245_, _13244_, _13243_);
  and (_13246_, _13245_, _05549_);
  or (_13247_, _13246_, _13242_);
  or (_13248_, _13247_, _05535_);
  and (_13249_, _13248_, _09805_);
  and (_13250_, _13249_, _13238_);
  or (_13251_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_13252_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  and (_13253_, _13252_, _13251_);
  and (_13254_, _13253_, _09792_);
  or (_13255_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_13256_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  and (_13257_, _13256_, _13255_);
  and (_13258_, _13257_, _05549_);
  or (_13259_, _13258_, _13254_);
  or (_13260_, _13259_, _09791_);
  or (_13261_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_13262_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  and (_13263_, _13262_, _13261_);
  and (_13264_, _13263_, _09792_);
  or (_13265_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  or (_13266_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  and (_13267_, _13266_, _13265_);
  and (_13268_, _13267_, _05549_);
  or (_13269_, _13268_, _13264_);
  or (_13270_, _13269_, _05535_);
  and (_13271_, _13270_, _05542_);
  and (_13272_, _13271_, _13260_);
  or (_13273_, _13272_, _13250_);
  and (_13274_, _13273_, _05518_);
  and (_13275_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  and (_13276_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  or (_13277_, _13276_, _13275_);
  and (_13278_, _13277_, _09792_);
  and (_13279_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  and (_13280_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  or (_13281_, _13280_, _13279_);
  and (_13282_, _13281_, _05549_);
  or (_13283_, _13282_, _13278_);
  or (_13284_, _13283_, _09791_);
  and (_13285_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  and (_13286_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_13287_, _13286_, _13285_);
  and (_13288_, _13287_, _09792_);
  and (_13289_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  and (_13290_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  or (_13291_, _13290_, _13289_);
  and (_13292_, _13291_, _05549_);
  or (_13293_, _13292_, _13288_);
  or (_13294_, _13293_, _05535_);
  and (_13295_, _13294_, _09805_);
  and (_13296_, _13295_, _13284_);
  or (_13297_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  or (_13298_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  and (_13299_, _13298_, _05549_);
  and (_13300_, _13299_, _13297_);
  or (_13301_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_13302_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  and (_13303_, _13302_, _09792_);
  and (_13304_, _13303_, _13301_);
  or (_13305_, _13304_, _13300_);
  or (_13306_, _13305_, _09791_);
  or (_13307_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  or (_13308_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  and (_13309_, _13308_, _05549_);
  and (_13310_, _13309_, _13307_);
  or (_13311_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_13312_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  and (_13313_, _13312_, _09792_);
  and (_13314_, _13313_, _13311_);
  or (_13315_, _13314_, _13310_);
  or (_13316_, _13315_, _05535_);
  and (_13317_, _13316_, _05542_);
  and (_13318_, _13317_, _13306_);
  or (_13319_, _13318_, _13296_);
  and (_13320_, _13319_, _09850_);
  or (_13321_, _13320_, _13274_);
  and (_13322_, _13321_, _09790_);
  and (_13323_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_13324_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_13325_, _13324_, _13323_);
  and (_13326_, _13325_, _09792_);
  and (_13327_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_13328_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_13329_, _13328_, _13327_);
  and (_13330_, _13329_, _05549_);
  or (_13331_, _13330_, _13326_);
  and (_13332_, _13331_, _05535_);
  and (_13333_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_13334_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_13335_, _13334_, _13333_);
  and (_13336_, _13335_, _09792_);
  and (_13337_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_13338_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_13339_, _13338_, _13337_);
  and (_13340_, _13339_, _05549_);
  or (_13341_, _13340_, _13336_);
  and (_13342_, _13341_, _09791_);
  or (_13343_, _13342_, _13332_);
  and (_13344_, _13343_, _09805_);
  or (_13345_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or (_13346_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_13347_, _13346_, _05549_);
  and (_13348_, _13347_, _13345_);
  or (_13349_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  or (_13350_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_13351_, _13350_, _09792_);
  and (_13352_, _13351_, _13349_);
  or (_13353_, _13352_, _13348_);
  and (_13354_, _13353_, _05535_);
  or (_13355_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or (_13356_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_13357_, _13356_, _05549_);
  and (_13358_, _13357_, _13355_);
  or (_13359_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_13360_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_13361_, _13360_, _09792_);
  and (_13362_, _13361_, _13359_);
  or (_13363_, _13362_, _13358_);
  and (_13364_, _13363_, _09791_);
  or (_13365_, _13364_, _13354_);
  and (_13366_, _13365_, _05542_);
  or (_13367_, _13366_, _13344_);
  and (_13368_, _13367_, _09850_);
  and (_13369_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  and (_13370_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  or (_13371_, _13370_, _13369_);
  and (_13372_, _13371_, _09792_);
  and (_13373_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  and (_13374_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  or (_13375_, _13374_, _13373_);
  and (_13376_, _13375_, _05549_);
  or (_13377_, _13376_, _13372_);
  and (_13378_, _13377_, _05535_);
  and (_13379_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  and (_13380_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_13381_, _13380_, _13379_);
  and (_13382_, _13381_, _09792_);
  and (_13383_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  and (_13384_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  or (_13385_, _13384_, _13383_);
  and (_13386_, _13385_, _05549_);
  or (_13387_, _13386_, _13382_);
  and (_13388_, _13387_, _09791_);
  or (_13389_, _13388_, _13378_);
  and (_13390_, _13389_, _09805_);
  or (_13391_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_13392_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  and (_13393_, _13392_, _13391_);
  and (_13394_, _13393_, _09792_);
  or (_13395_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  or (_13396_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  and (_13397_, _13396_, _13395_);
  and (_13398_, _13397_, _05549_);
  or (_13399_, _13398_, _13394_);
  and (_13400_, _13399_, _05535_);
  or (_13401_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  or (_13402_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  and (_13403_, _13402_, _13401_);
  and (_13404_, _13403_, _09792_);
  or (_13405_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  or (_13406_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  and (_13407_, _13406_, _13405_);
  and (_13408_, _13407_, _05549_);
  or (_13409_, _13408_, _13404_);
  and (_13410_, _13409_, _09791_);
  or (_13411_, _13410_, _13400_);
  and (_13412_, _13411_, _05542_);
  or (_13413_, _13412_, _13390_);
  and (_13414_, _13413_, _05518_);
  or (_13415_, _13414_, _13368_);
  and (_13416_, _13415_, _05520_);
  or (_13417_, _13416_, _13322_);
  or (_13418_, _13417_, _05526_);
  and (_13419_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  and (_13420_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_13421_, _13420_, _13419_);
  and (_13422_, _13421_, _09792_);
  and (_13423_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  and (_13424_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_13425_, _13424_, _13423_);
  and (_13426_, _13425_, _05549_);
  or (_13427_, _13426_, _13422_);
  or (_13428_, _13427_, _09791_);
  and (_13429_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  and (_13430_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_13431_, _13430_, _13429_);
  and (_13432_, _13431_, _09792_);
  and (_13433_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  and (_13434_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_13435_, _13434_, _13433_);
  and (_13436_, _13435_, _05549_);
  or (_13437_, _13436_, _13432_);
  or (_13438_, _13437_, _05535_);
  and (_13439_, _13438_, _09805_);
  and (_13440_, _13439_, _13428_);
  or (_13441_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_13442_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  and (_13443_, _13442_, _05549_);
  and (_13444_, _13443_, _13441_);
  or (_13445_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_13446_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  and (_13447_, _13446_, _09792_);
  and (_13448_, _13447_, _13445_);
  or (_13449_, _13448_, _13444_);
  or (_13450_, _13449_, _09791_);
  or (_13451_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_13452_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  and (_13453_, _13452_, _05549_);
  and (_13454_, _13453_, _13451_);
  or (_13455_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_13456_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  and (_13457_, _13456_, _09792_);
  and (_13458_, _13457_, _13455_);
  or (_13459_, _13458_, _13454_);
  or (_13460_, _13459_, _05535_);
  and (_13461_, _13460_, _05542_);
  and (_13462_, _13461_, _13450_);
  or (_13463_, _13462_, _13440_);
  and (_13464_, _13463_, _09850_);
  and (_13465_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  and (_13466_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  or (_13467_, _13466_, _13465_);
  and (_13468_, _13467_, _09792_);
  and (_13469_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  and (_13470_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_13471_, _13470_, _13469_);
  and (_13472_, _13471_, _05549_);
  or (_13473_, _13472_, _13468_);
  or (_13474_, _13473_, _09791_);
  and (_13475_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  and (_13476_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_13477_, _13476_, _13475_);
  and (_13478_, _13477_, _09792_);
  and (_13479_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  and (_13480_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_13481_, _13480_, _13479_);
  and (_13482_, _13481_, _05549_);
  or (_13483_, _13482_, _13478_);
  or (_13484_, _13483_, _05535_);
  and (_13485_, _13484_, _09805_);
  and (_13486_, _13485_, _13474_);
  or (_13487_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_13488_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  and (_13489_, _13488_, _13487_);
  and (_13490_, _13489_, _09792_);
  or (_13491_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_13492_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  and (_13493_, _13492_, _13491_);
  and (_13494_, _13493_, _05549_);
  or (_13495_, _13494_, _13490_);
  or (_13496_, _13495_, _09791_);
  or (_13497_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_13498_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  and (_13499_, _13498_, _13497_);
  and (_13500_, _13499_, _09792_);
  or (_13501_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  or (_13502_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  and (_13503_, _13502_, _13501_);
  and (_13504_, _13503_, _05549_);
  or (_13505_, _13504_, _13500_);
  or (_13506_, _13505_, _05535_);
  and (_13507_, _13506_, _05542_);
  and (_13508_, _13507_, _13496_);
  or (_13509_, _13508_, _13486_);
  and (_13510_, _13509_, _05518_);
  or (_13511_, _13510_, _13464_);
  and (_13512_, _13511_, _09790_);
  or (_13513_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_13514_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  and (_13515_, _13514_, _13513_);
  and (_13516_, _13515_, _09792_);
  or (_13517_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_13518_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  and (_13519_, _13518_, _13517_);
  and (_13520_, _13519_, _05549_);
  or (_13521_, _13520_, _13516_);
  and (_13522_, _13521_, _09791_);
  or (_13523_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_13524_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  and (_13525_, _13524_, _13523_);
  and (_13526_, _13525_, _09792_);
  or (_13527_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_13528_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  and (_13529_, _13528_, _13527_);
  and (_13530_, _13529_, _05549_);
  or (_13531_, _13530_, _13526_);
  and (_13532_, _13531_, _05535_);
  or (_13533_, _13532_, _13522_);
  and (_13534_, _13533_, _05542_);
  and (_13535_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  and (_13536_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  or (_13537_, _13536_, _13535_);
  and (_13538_, _13537_, _09792_);
  and (_13539_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  and (_13540_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_13541_, _13540_, _13539_);
  and (_13542_, _13541_, _05549_);
  or (_13543_, _13542_, _13538_);
  and (_13544_, _13543_, _09791_);
  and (_13545_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  and (_13546_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  or (_13547_, _13546_, _13545_);
  and (_13548_, _13547_, _09792_);
  and (_13549_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  and (_13550_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  or (_13551_, _13550_, _13549_);
  and (_13552_, _13551_, _05549_);
  or (_13553_, _13552_, _13548_);
  and (_13554_, _13553_, _05535_);
  or (_13555_, _13554_, _13544_);
  and (_13556_, _13555_, _09805_);
  or (_13557_, _13556_, _13534_);
  and (_13558_, _13557_, _05518_);
  or (_13559_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or (_13560_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  and (_13561_, _13560_, _05549_);
  and (_13562_, _13561_, _13559_);
  or (_13563_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or (_13564_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  and (_13565_, _13564_, _09792_);
  and (_13566_, _13565_, _13563_);
  or (_13567_, _13566_, _13562_);
  and (_13568_, _13567_, _09791_);
  or (_13569_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  or (_13570_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  and (_13571_, _13570_, _05549_);
  and (_13572_, _13571_, _13569_);
  or (_13573_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  or (_13574_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  and (_13575_, _13574_, _09792_);
  and (_13576_, _13575_, _13573_);
  or (_13577_, _13576_, _13572_);
  and (_13578_, _13577_, _05535_);
  or (_13579_, _13578_, _13568_);
  and (_13580_, _13579_, _05542_);
  and (_13581_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  and (_13582_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or (_13583_, _13582_, _13581_);
  and (_13584_, _13583_, _09792_);
  and (_13585_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  and (_13586_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or (_13587_, _13586_, _13585_);
  and (_13588_, _13587_, _05549_);
  or (_13589_, _13588_, _13584_);
  and (_13590_, _13589_, _09791_);
  and (_13591_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  and (_13592_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or (_13593_, _13592_, _13591_);
  and (_13594_, _13593_, _09792_);
  and (_13595_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  and (_13596_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or (_13597_, _13596_, _13595_);
  and (_13598_, _13597_, _05549_);
  or (_13599_, _13598_, _13594_);
  and (_13600_, _13599_, _05535_);
  or (_13601_, _13600_, _13590_);
  and (_13602_, _13601_, _09805_);
  or (_13603_, _13602_, _13580_);
  and (_13604_, _13603_, _09850_);
  or (_13605_, _13604_, _13558_);
  and (_13606_, _13605_, _05520_);
  or (_13607_, _13606_, _13512_);
  or (_13608_, _13607_, _10033_);
  and (_13609_, _13608_, _13418_);
  or (_13610_, _13609_, _00143_);
  and (_13611_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  and (_13612_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  or (_13613_, _13612_, _13611_);
  and (_13614_, _13613_, _09792_);
  and (_13615_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  and (_13616_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  or (_13617_, _13616_, _13615_);
  and (_13618_, _13617_, _05549_);
  or (_13619_, _13618_, _13614_);
  or (_13620_, _13619_, _09791_);
  and (_13621_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  and (_13622_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  or (_13623_, _13622_, _13621_);
  and (_13624_, _13623_, _09792_);
  and (_13625_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  and (_13626_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  or (_13627_, _13626_, _13625_);
  and (_13628_, _13627_, _05549_);
  or (_13629_, _13628_, _13624_);
  or (_13630_, _13629_, _05535_);
  and (_13631_, _13630_, _09805_);
  and (_13632_, _13631_, _13620_);
  or (_13633_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  or (_13634_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  and (_13635_, _13634_, _13633_);
  and (_13636_, _13635_, _09792_);
  or (_13637_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  or (_13638_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  and (_13639_, _13638_, _13637_);
  and (_13640_, _13639_, _05549_);
  or (_13641_, _13640_, _13636_);
  or (_13642_, _13641_, _09791_);
  or (_13643_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  or (_13644_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  and (_13645_, _13644_, _13643_);
  and (_13646_, _13645_, _09792_);
  or (_13647_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  or (_13648_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  and (_13649_, _13648_, _13647_);
  and (_13650_, _13649_, _05549_);
  or (_13651_, _13650_, _13646_);
  or (_13652_, _13651_, _05535_);
  and (_13653_, _13652_, _05542_);
  and (_13654_, _13653_, _13642_);
  or (_13655_, _13654_, _13632_);
  and (_13656_, _13655_, _05518_);
  and (_13657_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  and (_13658_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  or (_13659_, _13658_, _13657_);
  and (_13660_, _13659_, _09792_);
  and (_13661_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_13662_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  or (_13663_, _13662_, _13661_);
  and (_13664_, _13663_, _05549_);
  or (_13665_, _13664_, _13660_);
  or (_13666_, _13665_, _09791_);
  and (_13667_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  and (_13668_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  or (_13669_, _13668_, _13667_);
  and (_13670_, _13669_, _09792_);
  and (_13671_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_13672_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  or (_13673_, _13672_, _13671_);
  and (_13674_, _13673_, _05549_);
  or (_13675_, _13674_, _13670_);
  or (_13676_, _13675_, _05535_);
  and (_13677_, _13676_, _09805_);
  and (_13678_, _13677_, _13666_);
  or (_13679_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  or (_13680_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  and (_13681_, _13680_, _05549_);
  and (_13682_, _13681_, _13679_);
  or (_13683_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  or (_13684_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_13685_, _13684_, _09792_);
  and (_13686_, _13685_, _13683_);
  or (_13687_, _13686_, _13682_);
  or (_13688_, _13687_, _09791_);
  or (_13689_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  or (_13690_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  and (_13691_, _13690_, _05549_);
  and (_13692_, _13691_, _13689_);
  or (_13693_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  or (_13694_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  and (_13695_, _13694_, _09792_);
  and (_13696_, _13695_, _13693_);
  or (_13697_, _13696_, _13692_);
  or (_13698_, _13697_, _05535_);
  and (_13699_, _13698_, _05542_);
  and (_13700_, _13699_, _13688_);
  or (_13701_, _13700_, _13678_);
  and (_13702_, _13701_, _09850_);
  or (_13703_, _13702_, _13656_);
  and (_13704_, _13703_, _09790_);
  and (_13705_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  and (_13706_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or (_13707_, _13706_, _13705_);
  and (_13708_, _13707_, _09792_);
  and (_13709_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  and (_13710_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or (_13711_, _13710_, _13709_);
  and (_13712_, _13711_, _05549_);
  or (_13713_, _13712_, _13708_);
  and (_13714_, _13713_, _05535_);
  and (_13715_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  and (_13716_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or (_13717_, _13716_, _13715_);
  and (_13718_, _13717_, _09792_);
  and (_13719_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  and (_13720_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or (_13721_, _13720_, _13719_);
  and (_13722_, _13721_, _05549_);
  or (_13723_, _13722_, _13718_);
  and (_13724_, _13723_, _09791_);
  or (_13725_, _13724_, _13714_);
  and (_13726_, _13725_, _09805_);
  or (_13727_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or (_13728_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  and (_13729_, _13728_, _05549_);
  and (_13730_, _13729_, _13727_);
  or (_13731_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or (_13732_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  and (_13733_, _13732_, _09792_);
  and (_13734_, _13733_, _13731_);
  or (_13735_, _13734_, _13730_);
  and (_13736_, _13735_, _05535_);
  or (_13737_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or (_13738_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  and (_13739_, _13738_, _05549_);
  and (_13740_, _13739_, _13737_);
  or (_13741_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or (_13742_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  and (_13743_, _13742_, _09792_);
  and (_13744_, _13743_, _13741_);
  or (_13745_, _13744_, _13740_);
  and (_13746_, _13745_, _09791_);
  or (_13747_, _13746_, _13736_);
  and (_13748_, _13747_, _05542_);
  or (_13749_, _13748_, _13726_);
  and (_13750_, _13749_, _09850_);
  and (_13751_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  and (_13752_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or (_13753_, _13752_, _13751_);
  and (_13754_, _13753_, _09792_);
  and (_13755_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  and (_13756_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or (_13757_, _13756_, _13755_);
  and (_13758_, _13757_, _05549_);
  or (_13759_, _13758_, _13754_);
  and (_13760_, _13759_, _05535_);
  and (_13761_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  and (_13762_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or (_13763_, _13762_, _13761_);
  and (_13764_, _13763_, _09792_);
  and (_13765_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  and (_13766_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or (_13767_, _13766_, _13765_);
  and (_13768_, _13767_, _05549_);
  or (_13769_, _13768_, _13764_);
  and (_13770_, _13769_, _09791_);
  or (_13771_, _13770_, _13760_);
  and (_13772_, _13771_, _09805_);
  or (_13773_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or (_13774_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  and (_13775_, _13774_, _13773_);
  and (_13776_, _13775_, _09792_);
  or (_13777_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  or (_13778_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  and (_13779_, _13778_, _13777_);
  and (_13780_, _13779_, _05549_);
  or (_13781_, _13780_, _13776_);
  and (_13782_, _13781_, _05535_);
  or (_13783_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or (_13784_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  and (_13785_, _13784_, _13783_);
  and (_13786_, _13785_, _09792_);
  or (_13787_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  or (_13788_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  and (_13789_, _13788_, _13787_);
  and (_13790_, _13789_, _05549_);
  or (_13791_, _13790_, _13786_);
  and (_13792_, _13791_, _09791_);
  or (_13793_, _13792_, _13782_);
  and (_13794_, _13793_, _05542_);
  or (_13795_, _13794_, _13772_);
  and (_13796_, _13795_, _05518_);
  or (_13797_, _13796_, _13750_);
  and (_13798_, _13797_, _05520_);
  or (_13799_, _13798_, _13704_);
  or (_13800_, _13799_, _05526_);
  and (_13801_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  and (_13802_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  or (_13803_, _13802_, _13801_);
  and (_13804_, _13803_, _09792_);
  and (_13805_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  and (_13806_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  or (_13807_, _13806_, _13805_);
  and (_13808_, _13807_, _05549_);
  or (_13809_, _13808_, _13804_);
  or (_13810_, _13809_, _09791_);
  and (_13811_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  and (_13812_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_13813_, _13812_, _13811_);
  and (_13814_, _13813_, _09792_);
  and (_13815_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  and (_13816_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  or (_13817_, _13816_, _13815_);
  and (_13818_, _13817_, _05549_);
  or (_13819_, _13818_, _13814_);
  or (_13820_, _13819_, _05535_);
  and (_13821_, _13820_, _09805_);
  and (_13822_, _13821_, _13810_);
  or (_13823_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  or (_13824_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  and (_13825_, _13824_, _05549_);
  and (_13826_, _13825_, _13823_);
  or (_13827_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  or (_13828_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  and (_13829_, _13828_, _09792_);
  and (_13830_, _13829_, _13827_);
  or (_13831_, _13830_, _13826_);
  or (_13832_, _13831_, _09791_);
  or (_13833_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  or (_13834_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  and (_13835_, _13834_, _05549_);
  and (_13836_, _13835_, _13833_);
  or (_13837_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  or (_13838_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  and (_13839_, _13838_, _09792_);
  and (_13840_, _13839_, _13837_);
  or (_13841_, _13840_, _13836_);
  or (_13842_, _13841_, _05535_);
  and (_13843_, _13842_, _05542_);
  and (_13844_, _13843_, _13832_);
  or (_13845_, _13844_, _13822_);
  and (_13846_, _13845_, _09850_);
  and (_13847_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  and (_13848_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  or (_13849_, _13848_, _13847_);
  and (_13850_, _13849_, _09792_);
  and (_13851_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  and (_13852_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  or (_13853_, _13852_, _13851_);
  and (_13854_, _13853_, _05549_);
  or (_13855_, _13854_, _13850_);
  or (_13856_, _13855_, _09791_);
  and (_13857_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  and (_13858_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or (_13859_, _13858_, _13857_);
  and (_13860_, _13859_, _09792_);
  and (_13861_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  and (_13862_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  or (_13863_, _13862_, _13861_);
  and (_13864_, _13863_, _05549_);
  or (_13865_, _13864_, _13860_);
  or (_13866_, _13865_, _05535_);
  and (_13867_, _13866_, _09805_);
  and (_13868_, _13867_, _13856_);
  or (_13869_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or (_13870_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  and (_13871_, _13870_, _13869_);
  and (_13872_, _13871_, _09792_);
  or (_13873_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  or (_13874_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  and (_13875_, _13874_, _13873_);
  and (_13876_, _13875_, _05549_);
  or (_13877_, _13876_, _13872_);
  or (_13878_, _13877_, _09791_);
  or (_13879_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  or (_13880_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  and (_13881_, _13880_, _13879_);
  and (_13882_, _13881_, _09792_);
  or (_13883_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  or (_13884_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  and (_13885_, _13884_, _13883_);
  and (_13886_, _13885_, _05549_);
  or (_13887_, _13886_, _13882_);
  or (_13888_, _13887_, _05535_);
  and (_13889_, _13888_, _05542_);
  and (_13890_, _13889_, _13878_);
  or (_13891_, _13890_, _13868_);
  and (_13892_, _13891_, _05518_);
  or (_13893_, _13892_, _13846_);
  and (_13894_, _13893_, _09790_);
  or (_13895_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  or (_13896_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  and (_13897_, _13896_, _13895_);
  and (_13898_, _13897_, _09792_);
  or (_13899_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  or (_13900_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  and (_13901_, _13900_, _13899_);
  and (_13902_, _13901_, _05549_);
  or (_13903_, _13902_, _13898_);
  and (_13904_, _13903_, _09791_);
  or (_13905_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  or (_13906_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  and (_13907_, _13906_, _13905_);
  and (_13908_, _13907_, _09792_);
  or (_13909_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  or (_13910_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  and (_13911_, _13910_, _13909_);
  and (_13912_, _13911_, _05549_);
  or (_13913_, _13912_, _13908_);
  and (_13914_, _13913_, _05535_);
  or (_13915_, _13914_, _13904_);
  and (_13916_, _13915_, _05542_);
  and (_13917_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  and (_13918_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  or (_13919_, _13918_, _13917_);
  and (_13920_, _13919_, _09792_);
  and (_13921_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  and (_13922_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  or (_13923_, _13922_, _13921_);
  and (_13924_, _13923_, _05549_);
  or (_13925_, _13924_, _13920_);
  and (_13926_, _13925_, _09791_);
  and (_13927_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  and (_13928_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  or (_13929_, _13928_, _13927_);
  and (_13930_, _13929_, _09792_);
  and (_13931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  and (_13932_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  or (_13933_, _13932_, _13931_);
  and (_13934_, _13933_, _05549_);
  or (_13935_, _13934_, _13930_);
  and (_13936_, _13935_, _05535_);
  or (_13937_, _13936_, _13926_);
  and (_13938_, _13937_, _09805_);
  or (_13939_, _13938_, _13916_);
  and (_13940_, _13939_, _05518_);
  or (_13941_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  or (_13942_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  and (_13943_, _13942_, _05549_);
  and (_13944_, _13943_, _13941_);
  or (_13945_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_13946_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  and (_13947_, _13946_, _09792_);
  and (_13948_, _13947_, _13945_);
  or (_13949_, _13948_, _13944_);
  and (_13950_, _13949_, _09791_);
  or (_13951_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  or (_13952_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  and (_13953_, _13952_, _05549_);
  and (_13954_, _13953_, _13951_);
  or (_13955_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  or (_13956_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  and (_13957_, _13956_, _09792_);
  and (_13958_, _13957_, _13955_);
  or (_13959_, _13958_, _13954_);
  and (_13960_, _13959_, _05535_);
  or (_13961_, _13960_, _13950_);
  and (_13962_, _13961_, _05542_);
  and (_13963_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  and (_13964_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  or (_13965_, _13964_, _13963_);
  and (_13966_, _13965_, _09792_);
  and (_13967_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  and (_13968_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_13969_, _13968_, _13967_);
  and (_13970_, _13969_, _05549_);
  or (_13971_, _13970_, _13966_);
  and (_13972_, _13971_, _09791_);
  and (_13973_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  and (_13974_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_13975_, _13974_, _13973_);
  and (_13976_, _13975_, _09792_);
  and (_13977_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  and (_13978_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  or (_13979_, _13978_, _13977_);
  and (_13980_, _13979_, _05549_);
  or (_13981_, _13980_, _13976_);
  and (_13982_, _13981_, _05535_);
  or (_13983_, _13982_, _13972_);
  and (_13984_, _13983_, _09805_);
  or (_13985_, _13984_, _13962_);
  and (_13986_, _13985_, _09850_);
  or (_13987_, _13986_, _13940_);
  and (_13988_, _13987_, _05520_);
  or (_13989_, _13988_, _13894_);
  or (_13990_, _13989_, _10033_);
  and (_13991_, _13990_, _13800_);
  or (_13992_, _13991_, _04413_);
  and (_13993_, _13992_, _13610_);
  or (_13994_, _13993_, _05563_);
  or (_13995_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_13996_, _13995_, _22731_);
  and (_04717_, _13996_, _13994_);
  and (_13997_, _12438_, _24051_);
  and (_13998_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  or (_04720_, _13998_, _13997_);
  and (_13999_, _12438_, _24089_);
  and (_14000_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  or (_04728_, _14000_, _13999_);
  and (_14001_, _07013_, _24134_);
  and (_14002_, _07015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  or (_04731_, _14002_, _14001_);
  and (_14003_, _12442_, _24051_);
  and (_14004_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  or (_04734_, _14004_, _14003_);
  and (_14005_, _12442_, _23996_);
  and (_14006_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  or (_04740_, _14006_, _14005_);
  and (_14007_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  and (_14008_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  or (_14009_, _14008_, _14007_);
  and (_14010_, _14009_, _09792_);
  and (_14011_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  and (_14012_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  or (_14013_, _14012_, _14011_);
  and (_14014_, _14013_, _05549_);
  or (_14015_, _14014_, _14010_);
  or (_14016_, _14015_, _09791_);
  and (_14017_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  and (_14018_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_14019_, _14018_, _14017_);
  and (_14020_, _14019_, _09792_);
  and (_14021_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  and (_14022_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_14023_, _14022_, _14021_);
  and (_14024_, _14023_, _05549_);
  or (_14025_, _14024_, _14020_);
  or (_14026_, _14025_, _05535_);
  and (_14027_, _14026_, _09805_);
  and (_14028_, _14027_, _14016_);
  or (_14029_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  or (_14030_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  and (_14031_, _14030_, _14029_);
  and (_14032_, _14031_, _09792_);
  or (_14033_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  or (_14034_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  and (_14035_, _14034_, _14033_);
  and (_14036_, _14035_, _05549_);
  or (_14037_, _14036_, _14032_);
  or (_14038_, _14037_, _09791_);
  or (_14039_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  or (_14040_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  and (_14041_, _14040_, _14039_);
  and (_14042_, _14041_, _09792_);
  or (_14043_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  or (_14044_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  and (_14045_, _14044_, _14043_);
  and (_14046_, _14045_, _05549_);
  or (_14047_, _14046_, _14042_);
  or (_14048_, _14047_, _05535_);
  and (_14049_, _14048_, _05542_);
  and (_14050_, _14049_, _14038_);
  or (_14051_, _14050_, _14028_);
  or (_14052_, _14051_, _09850_);
  and (_14053_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  and (_14054_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  or (_14055_, _14054_, _14053_);
  and (_14056_, _14055_, _09792_);
  and (_14057_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  and (_14058_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  or (_14059_, _14058_, _14057_);
  and (_14060_, _14059_, _05549_);
  or (_14061_, _14060_, _14056_);
  or (_14062_, _14061_, _09791_);
  and (_14063_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  and (_14064_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  or (_14065_, _14064_, _14063_);
  and (_14066_, _14065_, _09792_);
  and (_14067_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  and (_14068_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  or (_14069_, _14068_, _14067_);
  and (_14070_, _14069_, _05549_);
  or (_14071_, _14070_, _14066_);
  or (_14072_, _14071_, _05535_);
  and (_14073_, _14072_, _09805_);
  and (_14074_, _14073_, _14062_);
  or (_14075_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  or (_14076_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  and (_14077_, _14076_, _05549_);
  and (_14078_, _14077_, _14075_);
  or (_14079_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_14080_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  and (_14081_, _14080_, _09792_);
  and (_14082_, _14081_, _14079_);
  or (_14083_, _14082_, _14078_);
  or (_14084_, _14083_, _09791_);
  or (_14085_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_14086_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  and (_14087_, _14086_, _05549_);
  and (_14088_, _14087_, _14085_);
  or (_14089_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_14090_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  and (_14091_, _14090_, _09792_);
  and (_14092_, _14091_, _14089_);
  or (_14093_, _14092_, _14088_);
  or (_14094_, _14093_, _05535_);
  and (_14095_, _14094_, _05542_);
  and (_14096_, _14095_, _14084_);
  or (_14097_, _14096_, _14074_);
  or (_14098_, _14097_, _05518_);
  and (_14099_, _14098_, _09790_);
  and (_14100_, _14099_, _14052_);
  and (_14101_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_14102_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_14103_, _14102_, _14101_);
  and (_14104_, _14103_, _09792_);
  and (_14105_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_14106_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_14107_, _14106_, _14105_);
  and (_14108_, _14107_, _05549_);
  or (_14109_, _14108_, _14104_);
  and (_14110_, _14109_, _05535_);
  and (_14111_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_14112_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_14113_, _14112_, _14111_);
  and (_14114_, _14113_, _09792_);
  and (_14115_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and (_14116_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  or (_14117_, _14116_, _14115_);
  and (_14118_, _14117_, _05549_);
  or (_14119_, _14118_, _14114_);
  and (_14120_, _14119_, _09791_);
  or (_14121_, _14120_, _05542_);
  or (_14122_, _14121_, _14110_);
  or (_14123_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_14124_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and (_14125_, _14124_, _05549_);
  and (_14126_, _14125_, _14123_);
  or (_14127_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_14128_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_14129_, _14128_, _09792_);
  and (_14130_, _14129_, _14127_);
  or (_14131_, _14130_, _14126_);
  and (_14132_, _14131_, _05535_);
  or (_14133_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_14134_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_14135_, _14134_, _05549_);
  and (_14136_, _14135_, _14133_);
  or (_14137_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_14138_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_14139_, _14138_, _09792_);
  and (_14140_, _14139_, _14137_);
  or (_14141_, _14140_, _14136_);
  and (_14142_, _14141_, _09791_);
  or (_14143_, _14142_, _09805_);
  or (_14144_, _14143_, _14132_);
  and (_14145_, _14144_, _14122_);
  or (_14146_, _14145_, _05518_);
  and (_14147_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  and (_14148_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_14149_, _14148_, _14147_);
  and (_14150_, _14149_, _09792_);
  and (_14151_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  and (_14152_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_14153_, _14152_, _14151_);
  and (_14154_, _14153_, _05549_);
  or (_14155_, _14154_, _14150_);
  and (_14156_, _14155_, _05535_);
  and (_14157_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  and (_14158_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  or (_14159_, _14158_, _14157_);
  and (_14160_, _14159_, _09792_);
  and (_14161_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  and (_14162_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  or (_14163_, _14162_, _14161_);
  and (_14164_, _14163_, _05549_);
  or (_14165_, _14164_, _14160_);
  and (_14166_, _14165_, _09791_);
  or (_14167_, _14166_, _05542_);
  or (_14168_, _14167_, _14156_);
  or (_14169_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  or (_14170_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  and (_14171_, _14170_, _14169_);
  and (_14172_, _14171_, _09792_);
  or (_14173_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  or (_14174_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  and (_14175_, _14174_, _14173_);
  and (_14176_, _14175_, _05549_);
  or (_14177_, _14176_, _14172_);
  and (_14178_, _14177_, _05535_);
  or (_14179_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  or (_14180_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  and (_14181_, _14180_, _14179_);
  and (_14182_, _14181_, _09792_);
  or (_14183_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  or (_14184_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  and (_14185_, _14184_, _14183_);
  and (_14186_, _14185_, _05549_);
  or (_14187_, _14186_, _14182_);
  and (_14188_, _14187_, _09791_);
  or (_14189_, _14188_, _09805_);
  or (_14190_, _14189_, _14178_);
  and (_14191_, _14190_, _14168_);
  or (_14192_, _14191_, _09850_);
  and (_14193_, _14192_, _05520_);
  and (_14194_, _14193_, _14146_);
  or (_14195_, _14194_, _14100_);
  or (_14196_, _14195_, _05526_);
  and (_14197_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  and (_14198_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or (_14199_, _14198_, _14197_);
  and (_14200_, _14199_, _09792_);
  and (_14201_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  and (_14202_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or (_14203_, _14202_, _14201_);
  and (_14204_, _14203_, _05549_);
  or (_14205_, _14204_, _14200_);
  and (_14206_, _14205_, _05535_);
  and (_14207_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  and (_14208_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or (_14209_, _14208_, _14207_);
  and (_14210_, _14209_, _09792_);
  and (_14211_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  and (_14212_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  or (_14213_, _14212_, _14211_);
  and (_14214_, _14213_, _05549_);
  or (_14215_, _14214_, _14210_);
  and (_14216_, _14215_, _09791_);
  or (_14217_, _14216_, _05542_);
  or (_14218_, _14217_, _14206_);
  or (_14219_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  or (_14220_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  and (_14221_, _14220_, _14219_);
  and (_14222_, _14221_, _09792_);
  or (_14223_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or (_14224_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  and (_14225_, _14224_, _14223_);
  and (_14226_, _14225_, _05549_);
  or (_14227_, _14226_, _14222_);
  and (_14228_, _14227_, _05535_);
  or (_14229_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or (_14230_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  and (_14231_, _14230_, _14229_);
  and (_14232_, _14231_, _09792_);
  or (_14233_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or (_14234_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  and (_14235_, _14234_, _14233_);
  and (_14236_, _14235_, _05549_);
  or (_14237_, _14236_, _14232_);
  and (_14238_, _14237_, _09791_);
  or (_14239_, _14238_, _09805_);
  or (_14240_, _14239_, _14228_);
  and (_14241_, _14240_, _14218_);
  or (_14242_, _14241_, _05518_);
  and (_14243_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  and (_14244_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_14245_, _14244_, _14243_);
  and (_14246_, _14245_, _09792_);
  and (_14247_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  and (_14248_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  or (_14249_, _14248_, _14247_);
  and (_14250_, _14249_, _05549_);
  or (_14251_, _14250_, _14246_);
  and (_14252_, _14251_, _05535_);
  and (_14253_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  and (_14254_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_14255_, _14254_, _14253_);
  and (_14256_, _14255_, _09792_);
  and (_14257_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  and (_14258_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  or (_14259_, _14258_, _14257_);
  and (_14260_, _14259_, _05549_);
  or (_14261_, _14260_, _14256_);
  and (_14262_, _14261_, _09791_);
  or (_14263_, _14262_, _05542_);
  or (_14264_, _14263_, _14252_);
  or (_14265_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_14266_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  and (_14267_, _14266_, _14265_);
  and (_14269_, _14267_, _09792_);
  or (_14270_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_14271_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  and (_14272_, _14271_, _14270_);
  and (_14273_, _14272_, _05549_);
  or (_14274_, _14273_, _14269_);
  and (_14275_, _14274_, _05535_);
  or (_14276_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_14277_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  and (_14278_, _14277_, _14276_);
  and (_14279_, _14278_, _09792_);
  or (_14280_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_14281_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  and (_14282_, _14281_, _14280_);
  and (_14283_, _14282_, _05549_);
  or (_14284_, _14283_, _14279_);
  and (_14285_, _14284_, _09791_);
  or (_14286_, _14285_, _09805_);
  or (_14287_, _14286_, _14275_);
  and (_14288_, _14287_, _14264_);
  or (_14289_, _14288_, _09850_);
  and (_14290_, _14289_, _05520_);
  and (_14291_, _14290_, _14242_);
  and (_14292_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  and (_14293_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_14294_, _14293_, _14292_);
  and (_14295_, _14294_, _05549_);
  and (_14296_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  and (_14297_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_14298_, _14297_, _14296_);
  and (_14299_, _14298_, _09792_);
  or (_14300_, _14299_, _14295_);
  or (_14301_, _14300_, _09791_);
  and (_14302_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  and (_14303_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_14304_, _14303_, _14302_);
  and (_14305_, _14304_, _05549_);
  and (_14306_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  and (_14307_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_14308_, _14307_, _14306_);
  and (_14309_, _14308_, _09792_);
  or (_14310_, _14309_, _14305_);
  or (_14311_, _14310_, _05535_);
  and (_14312_, _14311_, _09805_);
  and (_14313_, _14312_, _14301_);
  or (_14314_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_14315_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  and (_14316_, _14315_, _09792_);
  and (_14317_, _14316_, _14314_);
  or (_14318_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_14319_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  and (_14320_, _14319_, _05549_);
  and (_14321_, _14320_, _14318_);
  or (_14322_, _14321_, _14317_);
  or (_14323_, _14322_, _09791_);
  or (_14324_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_14325_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  and (_14326_, _14325_, _09792_);
  and (_14327_, _14326_, _14324_);
  or (_14328_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_14329_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  and (_14330_, _14329_, _05549_);
  and (_14331_, _14330_, _14328_);
  or (_14332_, _14331_, _14327_);
  or (_14333_, _14332_, _05535_);
  and (_14334_, _14333_, _05542_);
  and (_14335_, _14334_, _14323_);
  or (_14336_, _14335_, _14313_);
  and (_14337_, _14336_, _09850_);
  and (_14338_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  and (_14339_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_14340_, _14339_, _09792_);
  or (_14341_, _14340_, _14338_);
  and (_14342_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  and (_14343_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  or (_14344_, _14343_, _05549_);
  or (_14345_, _14344_, _14342_);
  and (_14346_, _14345_, _14341_);
  or (_14347_, _14346_, _09791_);
  and (_14348_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  and (_14349_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_14350_, _14349_, _09792_);
  or (_14351_, _14350_, _14348_);
  and (_14352_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  and (_14353_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_14354_, _14353_, _05549_);
  or (_14355_, _14354_, _14352_);
  and (_14356_, _14355_, _14351_);
  or (_14357_, _14356_, _05535_);
  and (_14358_, _14357_, _09805_);
  and (_14359_, _14358_, _14347_);
  or (_14360_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_14361_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  and (_14362_, _14361_, _14360_);
  or (_14363_, _14362_, _05549_);
  or (_14364_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_14365_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  and (_14366_, _14365_, _14364_);
  or (_14367_, _14366_, _09792_);
  and (_14368_, _14367_, _14363_);
  or (_14369_, _14368_, _09791_);
  or (_14370_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_14371_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  and (_14372_, _14371_, _14370_);
  or (_14373_, _14372_, _05549_);
  or (_14374_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_14375_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  and (_14376_, _14375_, _14374_);
  or (_14377_, _14376_, _09792_);
  and (_14378_, _14377_, _14373_);
  or (_14379_, _14378_, _05535_);
  and (_14380_, _14379_, _05542_);
  and (_14381_, _14380_, _14369_);
  or (_14382_, _14381_, _14359_);
  and (_14383_, _14382_, _05518_);
  or (_14384_, _14383_, _14337_);
  and (_14385_, _14384_, _09790_);
  or (_14386_, _14385_, _14291_);
  or (_14387_, _14386_, _10033_);
  and (_14388_, _14387_, _14196_);
  or (_14389_, _14388_, _00143_);
  and (_14390_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  and (_14391_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  or (_14392_, _14391_, _14390_);
  and (_14393_, _14392_, _09792_);
  and (_14394_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  and (_14395_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  or (_14396_, _14395_, _14394_);
  and (_14397_, _14396_, _05549_);
  or (_14398_, _14397_, _14393_);
  or (_14399_, _14398_, _09791_);
  and (_14400_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  and (_14401_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  or (_14402_, _14401_, _14400_);
  and (_14403_, _14402_, _09792_);
  and (_14404_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  and (_14405_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  or (_14406_, _14405_, _14404_);
  and (_14407_, _14406_, _05549_);
  or (_14408_, _14407_, _14403_);
  or (_14409_, _14408_, _05535_);
  and (_14410_, _14409_, _09805_);
  and (_14411_, _14410_, _14399_);
  or (_14412_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  or (_14413_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  and (_14414_, _14413_, _14412_);
  and (_14415_, _14414_, _09792_);
  or (_14416_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  or (_14417_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  and (_14418_, _14417_, _14416_);
  and (_14419_, _14418_, _05549_);
  or (_14420_, _14419_, _14415_);
  or (_14421_, _14420_, _09791_);
  or (_14422_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  or (_14423_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  and (_14424_, _14423_, _14422_);
  and (_14425_, _14424_, _09792_);
  or (_14426_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  or (_14427_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  and (_14428_, _14427_, _14426_);
  and (_14429_, _14428_, _05549_);
  or (_14430_, _14429_, _14425_);
  or (_14431_, _14430_, _05535_);
  and (_14432_, _14431_, _05542_);
  and (_14433_, _14432_, _14421_);
  or (_14434_, _14433_, _14411_);
  and (_14435_, _14434_, _05518_);
  and (_14436_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  and (_14437_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  or (_14438_, _14437_, _14436_);
  and (_14439_, _14438_, _09792_);
  and (_14440_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_14441_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  or (_14442_, _14441_, _14440_);
  and (_14443_, _14442_, _05549_);
  or (_14444_, _14443_, _14439_);
  or (_14445_, _14444_, _09791_);
  and (_14446_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  and (_14447_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  or (_14448_, _14447_, _14446_);
  and (_14449_, _14448_, _09792_);
  and (_14450_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_14451_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  or (_14452_, _14451_, _14450_);
  and (_14453_, _14452_, _05549_);
  or (_14454_, _14453_, _14449_);
  or (_14455_, _14454_, _05535_);
  and (_14456_, _14455_, _09805_);
  and (_14457_, _14456_, _14445_);
  or (_14458_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  or (_14459_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_14460_, _14459_, _05549_);
  and (_14461_, _14460_, _14458_);
  or (_14462_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  or (_14463_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  and (_14464_, _14463_, _09792_);
  and (_14465_, _14464_, _14462_);
  or (_14466_, _14465_, _14461_);
  or (_14467_, _14466_, _09791_);
  or (_14468_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  or (_14469_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  and (_14470_, _14469_, _05549_);
  and (_14471_, _14470_, _14468_);
  or (_14472_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  or (_14473_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_14474_, _14473_, _09792_);
  and (_14475_, _14474_, _14472_);
  or (_14476_, _14475_, _14471_);
  or (_14477_, _14476_, _05535_);
  and (_14478_, _14477_, _05542_);
  and (_14479_, _14478_, _14467_);
  or (_14480_, _14479_, _14457_);
  and (_14481_, _14480_, _09850_);
  or (_14482_, _14481_, _14435_);
  and (_14483_, _14482_, _09790_);
  and (_14484_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  and (_14485_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or (_14486_, _14485_, _14484_);
  and (_14487_, _14486_, _09792_);
  and (_14488_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  and (_14489_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or (_14490_, _14489_, _14488_);
  and (_14491_, _14490_, _05549_);
  or (_14492_, _14491_, _14487_);
  and (_14493_, _14492_, _05535_);
  and (_14494_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  and (_14495_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or (_14496_, _14495_, _14494_);
  and (_14497_, _14496_, _09792_);
  and (_14498_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  and (_14499_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  or (_14500_, _14499_, _14498_);
  and (_14501_, _14500_, _05549_);
  or (_14502_, _14501_, _14497_);
  and (_14503_, _14502_, _09791_);
  or (_14504_, _14503_, _14493_);
  and (_14505_, _14504_, _09805_);
  or (_14506_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or (_14507_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  and (_14508_, _14507_, _05549_);
  and (_14509_, _14508_, _14506_);
  or (_14510_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or (_14511_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  and (_14512_, _14511_, _09792_);
  and (_14513_, _14512_, _14510_);
  or (_14514_, _14513_, _14509_);
  and (_14515_, _14514_, _05535_);
  or (_14516_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or (_14517_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  and (_14518_, _14517_, _05549_);
  and (_14519_, _14518_, _14516_);
  or (_14520_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or (_14521_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  and (_14522_, _14521_, _09792_);
  and (_14523_, _14522_, _14520_);
  or (_14524_, _14523_, _14519_);
  and (_14525_, _14524_, _09791_);
  or (_14526_, _14525_, _14515_);
  and (_14527_, _14526_, _05542_);
  or (_14528_, _14527_, _14505_);
  and (_14529_, _14528_, _09850_);
  and (_14530_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  and (_14531_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or (_14532_, _14531_, _14530_);
  and (_14533_, _14532_, _09792_);
  and (_14534_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  and (_14535_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or (_14536_, _14535_, _14534_);
  and (_14537_, _14536_, _05549_);
  or (_14538_, _14537_, _14533_);
  and (_14539_, _14538_, _05535_);
  and (_14540_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  and (_14541_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or (_14542_, _14541_, _14540_);
  and (_14543_, _14542_, _09792_);
  and (_14544_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  and (_14545_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or (_14546_, _14545_, _14544_);
  and (_14547_, _14546_, _05549_);
  or (_14548_, _14547_, _14543_);
  and (_14549_, _14548_, _09791_);
  or (_14550_, _14549_, _14539_);
  and (_14551_, _14550_, _09805_);
  or (_14552_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or (_14553_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  and (_14554_, _14553_, _14552_);
  and (_14555_, _14554_, _09792_);
  or (_14556_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  or (_14557_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  and (_14558_, _14557_, _14556_);
  and (_14559_, _14558_, _05549_);
  or (_14560_, _14559_, _14555_);
  and (_14561_, _14560_, _05535_);
  or (_14562_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  or (_14563_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  and (_14564_, _14563_, _14562_);
  and (_14565_, _14564_, _09792_);
  or (_14566_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or (_14567_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  and (_14568_, _14567_, _14566_);
  and (_14569_, _14568_, _05549_);
  or (_14570_, _14569_, _14565_);
  and (_14571_, _14570_, _09791_);
  or (_14572_, _14571_, _14561_);
  and (_14573_, _14572_, _05542_);
  or (_14574_, _14573_, _14551_);
  and (_14575_, _14574_, _05518_);
  or (_14576_, _14575_, _14529_);
  and (_14577_, _14576_, _05520_);
  or (_14578_, _14577_, _14483_);
  or (_14579_, _14578_, _05526_);
  and (_14580_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  and (_14581_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  or (_14582_, _14581_, _14580_);
  and (_14583_, _14582_, _09792_);
  and (_14584_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  and (_14585_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_14586_, _14585_, _14584_);
  and (_14587_, _14586_, _05549_);
  or (_14588_, _14587_, _14583_);
  or (_14589_, _14588_, _09791_);
  and (_14590_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  and (_14591_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  or (_14592_, _14591_, _14590_);
  and (_14593_, _14592_, _09792_);
  and (_14594_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  and (_14595_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  or (_14596_, _14595_, _14594_);
  and (_14597_, _14596_, _05549_);
  or (_14598_, _14597_, _14593_);
  or (_14599_, _14598_, _05535_);
  and (_14600_, _14599_, _09805_);
  and (_14601_, _14600_, _14589_);
  or (_14602_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  or (_14603_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  and (_14604_, _14603_, _05549_);
  and (_14605_, _14604_, _14602_);
  or (_14606_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  or (_14607_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  and (_14608_, _14607_, _09792_);
  and (_14609_, _14608_, _14606_);
  or (_14610_, _14609_, _14605_);
  or (_14611_, _14610_, _09791_);
  or (_14612_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  or (_14613_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  and (_14614_, _14613_, _05549_);
  and (_14615_, _14614_, _14612_);
  or (_14616_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  or (_14617_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  and (_14618_, _14617_, _09792_);
  and (_14619_, _14618_, _14616_);
  or (_14620_, _14619_, _14615_);
  or (_14621_, _14620_, _05535_);
  and (_14622_, _14621_, _05542_);
  and (_14623_, _14622_, _14611_);
  or (_14624_, _14623_, _14601_);
  and (_14625_, _14624_, _09850_);
  and (_14626_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  and (_14627_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  or (_14628_, _14627_, _14626_);
  and (_14629_, _14628_, _09792_);
  and (_14630_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  and (_14631_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or (_14632_, _14631_, _14630_);
  and (_14633_, _14632_, _05549_);
  or (_14634_, _14633_, _14629_);
  or (_14635_, _14634_, _09791_);
  and (_14636_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  and (_14637_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_14638_, _14637_, _14636_);
  and (_14639_, _14638_, _09792_);
  and (_14640_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  and (_14641_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  or (_14642_, _14641_, _14640_);
  and (_14643_, _14642_, _05549_);
  or (_14644_, _14643_, _14639_);
  or (_14645_, _14644_, _05535_);
  and (_14646_, _14645_, _09805_);
  and (_14647_, _14646_, _14635_);
  or (_14648_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_14649_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  and (_14650_, _14649_, _14648_);
  and (_14651_, _14650_, _09792_);
  or (_14652_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_14653_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  and (_14654_, _14653_, _14652_);
  and (_14655_, _14654_, _05549_);
  or (_14656_, _14655_, _14651_);
  or (_14657_, _14656_, _09791_);
  or (_14658_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or (_14659_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  and (_14660_, _14659_, _14658_);
  and (_14661_, _14660_, _09792_);
  or (_14662_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  or (_14663_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  and (_14664_, _14663_, _14662_);
  and (_14665_, _14664_, _05549_);
  or (_14666_, _14665_, _14661_);
  or (_14667_, _14666_, _05535_);
  and (_14668_, _14667_, _05542_);
  and (_14669_, _14668_, _14657_);
  or (_14670_, _14669_, _14647_);
  and (_14671_, _14670_, _05518_);
  or (_14672_, _14671_, _14625_);
  and (_14673_, _14672_, _09790_);
  or (_14674_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  or (_14675_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  and (_14676_, _14675_, _14674_);
  and (_14677_, _14676_, _09792_);
  or (_14678_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  or (_14679_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  and (_14680_, _14679_, _14678_);
  and (_14681_, _14680_, _05549_);
  or (_14682_, _14681_, _14677_);
  and (_14683_, _14682_, _09791_);
  or (_14684_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  or (_14685_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  and (_14686_, _14685_, _14684_);
  and (_14687_, _14686_, _09792_);
  or (_14688_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  or (_14689_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  and (_14690_, _14689_, _14688_);
  and (_14691_, _14690_, _05549_);
  or (_14692_, _14691_, _14687_);
  and (_14693_, _14692_, _05535_);
  or (_14694_, _14693_, _14683_);
  and (_14695_, _14694_, _05542_);
  and (_14696_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  and (_14697_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  or (_14698_, _14697_, _14696_);
  and (_14699_, _14698_, _09792_);
  and (_14700_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  and (_14701_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  or (_14702_, _14701_, _14700_);
  and (_14703_, _14702_, _05549_);
  or (_14704_, _14703_, _14699_);
  and (_14705_, _14704_, _09791_);
  and (_14706_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  and (_14707_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  or (_14708_, _14707_, _14706_);
  and (_14709_, _14708_, _09792_);
  and (_14710_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  and (_14711_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  or (_14712_, _14711_, _14710_);
  and (_14713_, _14712_, _05549_);
  or (_14714_, _14713_, _14709_);
  and (_14715_, _14714_, _05535_);
  or (_14716_, _14715_, _14705_);
  and (_14717_, _14716_, _09805_);
  or (_14718_, _14717_, _14695_);
  and (_14719_, _14718_, _05518_);
  or (_14720_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_14721_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  and (_14722_, _14721_, _05549_);
  and (_14723_, _14722_, _14720_);
  or (_14724_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_14725_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  and (_14726_, _14725_, _09792_);
  and (_14727_, _14726_, _14724_);
  or (_14728_, _14727_, _14723_);
  and (_14729_, _14728_, _09791_);
  or (_14730_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  or (_14731_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  and (_14732_, _14731_, _05549_);
  and (_14733_, _14732_, _14730_);
  or (_14734_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  or (_14735_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  and (_14736_, _14735_, _09792_);
  and (_14737_, _14736_, _14734_);
  or (_14738_, _14737_, _14733_);
  and (_14739_, _14738_, _05535_);
  or (_14740_, _14739_, _14729_);
  and (_14741_, _14740_, _05542_);
  and (_14742_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  and (_14743_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  or (_14744_, _14743_, _14742_);
  and (_14745_, _14744_, _09792_);
  and (_14746_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  and (_14747_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_14748_, _14747_, _14746_);
  and (_14749_, _14748_, _05549_);
  or (_14750_, _14749_, _14745_);
  and (_14751_, _14750_, _09791_);
  and (_14752_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  and (_14753_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  or (_14754_, _14753_, _14752_);
  and (_14755_, _14754_, _09792_);
  and (_14756_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  and (_14757_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  or (_14758_, _14757_, _14756_);
  and (_14759_, _14758_, _05549_);
  or (_14760_, _14759_, _14755_);
  and (_14761_, _14760_, _05535_);
  or (_14762_, _14761_, _14751_);
  and (_14763_, _14762_, _09805_);
  or (_14764_, _14763_, _14741_);
  and (_14765_, _14764_, _09850_);
  or (_14766_, _14765_, _14719_);
  and (_14767_, _14766_, _05520_);
  or (_14768_, _14767_, _14673_);
  or (_14769_, _14768_, _10033_);
  and (_14770_, _14769_, _14579_);
  or (_14771_, _14770_, _04413_);
  and (_14772_, _14771_, _14389_);
  or (_14773_, _14772_, _05563_);
  or (_14774_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_14775_, _14774_, _22731_);
  and (_04746_, _14775_, _14773_);
  and (_14776_, _12442_, _24134_);
  and (_14777_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  or (_04765_, _14777_, _14776_);
  and (_14778_, _24476_, _24016_);
  and (_14779_, _14778_, _24089_);
  not (_14780_, _14778_);
  and (_14781_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  or (_27188_, _14781_, _14779_);
  and (_14782_, _14778_, _23583_);
  and (_14783_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  or (_04771_, _14783_, _14782_);
  and (_14784_, _08435_, _24134_);
  and (_14785_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  or (_04776_, _14785_, _14784_);
  and (_14786_, _14778_, _23887_);
  and (_14787_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  or (_04784_, _14787_, _14786_);
  and (_14788_, _14778_, _23548_);
  and (_14789_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  or (_04788_, _14789_, _14788_);
  and (_14790_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  and (_14791_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_14792_, _14791_, _14790_);
  and (_14793_, _14792_, _09792_);
  and (_14794_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  and (_14795_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_14796_, _14795_, _14794_);
  and (_14797_, _14796_, _05549_);
  or (_14798_, _14797_, _14793_);
  or (_14799_, _14798_, _09791_);
  and (_14800_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  and (_14801_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_14802_, _14801_, _14800_);
  and (_14803_, _14802_, _09792_);
  and (_14804_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  and (_14805_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_14806_, _14805_, _14804_);
  and (_14807_, _14806_, _05549_);
  or (_14808_, _14807_, _14803_);
  or (_14809_, _14808_, _05535_);
  and (_14810_, _14809_, _09805_);
  and (_14811_, _14810_, _14799_);
  or (_14812_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_14813_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  and (_14814_, _14813_, _14812_);
  and (_14815_, _14814_, _09792_);
  or (_14816_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  or (_14817_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  and (_14818_, _14817_, _14816_);
  and (_14819_, _14818_, _05549_);
  or (_14820_, _14819_, _14815_);
  or (_14821_, _14820_, _09791_);
  or (_14822_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  or (_14823_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  and (_14824_, _14823_, _14822_);
  and (_14825_, _14824_, _09792_);
  or (_14826_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  or (_14827_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  and (_14828_, _14827_, _14826_);
  and (_14829_, _14828_, _05549_);
  or (_14830_, _14829_, _14825_);
  or (_14831_, _14830_, _05535_);
  and (_14832_, _14831_, _05542_);
  and (_14833_, _14832_, _14821_);
  or (_14834_, _14833_, _14811_);
  or (_14835_, _14834_, _09850_);
  and (_14836_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  and (_14837_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_14838_, _14837_, _14836_);
  and (_14839_, _14838_, _09792_);
  and (_14840_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  and (_14841_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_14842_, _14841_, _14840_);
  and (_14843_, _14842_, _05549_);
  or (_14844_, _14843_, _14839_);
  or (_14845_, _14844_, _09791_);
  and (_14846_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  and (_14847_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_14848_, _14847_, _14846_);
  and (_14849_, _14848_, _09792_);
  and (_14850_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  and (_14851_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_14852_, _14851_, _14850_);
  and (_14853_, _14852_, _05549_);
  or (_14854_, _14853_, _14849_);
  or (_14855_, _14854_, _05535_);
  and (_14856_, _14855_, _09805_);
  and (_14857_, _14856_, _14845_);
  or (_14858_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_14859_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  and (_14860_, _14859_, _05549_);
  and (_14861_, _14860_, _14858_);
  or (_14862_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  or (_14863_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  and (_14864_, _14863_, _09792_);
  and (_14865_, _14864_, _14862_);
  or (_14866_, _14865_, _14861_);
  or (_14867_, _14866_, _09791_);
  or (_14868_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  or (_14869_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  and (_14870_, _14869_, _05549_);
  and (_14871_, _14870_, _14868_);
  or (_14872_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_14873_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  and (_14874_, _14873_, _09792_);
  and (_14875_, _14874_, _14872_);
  or (_14876_, _14875_, _14871_);
  or (_14877_, _14876_, _05535_);
  and (_14878_, _14877_, _05542_);
  and (_14879_, _14878_, _14867_);
  or (_14880_, _14879_, _14857_);
  or (_14881_, _14880_, _05518_);
  and (_14882_, _14881_, _09790_);
  and (_14883_, _14882_, _14835_);
  and (_14884_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_14885_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_14886_, _14885_, _14884_);
  and (_14887_, _14886_, _09792_);
  and (_14888_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_14889_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_14890_, _14889_, _14888_);
  and (_14891_, _14890_, _05549_);
  or (_14892_, _14891_, _14887_);
  and (_14893_, _14892_, _05535_);
  and (_14894_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_14895_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_14896_, _14895_, _14894_);
  and (_14897_, _14896_, _09792_);
  and (_14898_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_14899_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_14900_, _14899_, _14898_);
  and (_14901_, _14900_, _05549_);
  or (_14902_, _14901_, _14897_);
  and (_14903_, _14902_, _09791_);
  or (_14904_, _14903_, _05542_);
  or (_14905_, _14904_, _14893_);
  or (_14906_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_14907_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_14908_, _14907_, _05549_);
  and (_14909_, _14908_, _14906_);
  or (_14910_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_14911_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_14912_, _14911_, _09792_);
  and (_14913_, _14912_, _14910_);
  or (_14914_, _14913_, _14909_);
  and (_14915_, _14914_, _05535_);
  or (_14916_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_14917_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_14918_, _14917_, _05549_);
  and (_14919_, _14918_, _14916_);
  or (_14920_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_14921_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_14922_, _14921_, _09792_);
  and (_14923_, _14922_, _14920_);
  or (_14924_, _14923_, _14919_);
  and (_14925_, _14924_, _09791_);
  or (_14926_, _14925_, _09805_);
  or (_14927_, _14926_, _14915_);
  and (_14928_, _14927_, _14905_);
  or (_14929_, _14928_, _05518_);
  and (_14930_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  and (_14931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  or (_14932_, _14931_, _14930_);
  and (_14933_, _14932_, _09792_);
  and (_14934_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  and (_14935_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_14936_, _14935_, _14934_);
  and (_14937_, _14936_, _05549_);
  or (_14938_, _14937_, _14933_);
  and (_14939_, _14938_, _05535_);
  and (_14940_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  and (_14941_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  or (_14942_, _14941_, _14940_);
  and (_14943_, _14942_, _09792_);
  and (_14944_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  and (_14945_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_14946_, _14945_, _14944_);
  and (_14947_, _14946_, _05549_);
  or (_14948_, _14947_, _14943_);
  and (_14949_, _14948_, _09791_);
  or (_14950_, _14949_, _05542_);
  or (_14951_, _14950_, _14939_);
  or (_14952_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  or (_14953_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  and (_14954_, _14953_, _14952_);
  and (_14955_, _14954_, _09792_);
  or (_14956_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_14957_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  and (_14958_, _14957_, _14956_);
  and (_14959_, _14958_, _05549_);
  or (_14960_, _14959_, _14955_);
  and (_14961_, _14960_, _05535_);
  or (_14962_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  or (_14963_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  and (_14964_, _14963_, _14962_);
  and (_14965_, _14964_, _09792_);
  or (_14966_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_14967_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  and (_14968_, _14967_, _14966_);
  and (_14969_, _14968_, _05549_);
  or (_14970_, _14969_, _14965_);
  and (_14971_, _14970_, _09791_);
  or (_14972_, _14971_, _09805_);
  or (_14973_, _14972_, _14961_);
  and (_14974_, _14973_, _14951_);
  or (_14975_, _14974_, _09850_);
  and (_14976_, _14975_, _05520_);
  and (_14977_, _14976_, _14929_);
  or (_14978_, _14977_, _14883_);
  or (_14979_, _14978_, _05526_);
  and (_14980_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  and (_14981_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or (_14982_, _14981_, _14980_);
  and (_14983_, _14982_, _09792_);
  and (_14984_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  and (_14985_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or (_14986_, _14985_, _14984_);
  and (_14987_, _14986_, _05549_);
  or (_14988_, _14987_, _14983_);
  and (_14989_, _14988_, _05535_);
  and (_14990_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  and (_14991_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  or (_14992_, _14991_, _14990_);
  and (_14993_, _14992_, _09792_);
  and (_14994_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  and (_14995_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or (_14996_, _14995_, _14994_);
  and (_14997_, _14996_, _05549_);
  or (_14998_, _14997_, _14993_);
  and (_14999_, _14998_, _09791_);
  or (_15000_, _14999_, _05542_);
  or (_15001_, _15000_, _14989_);
  or (_15002_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  or (_15003_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  and (_15004_, _15003_, _15002_);
  and (_15005_, _15004_, _09792_);
  or (_15006_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or (_15007_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  and (_15008_, _15007_, _15006_);
  and (_15009_, _15008_, _05549_);
  or (_15010_, _15009_, _15005_);
  and (_15011_, _15010_, _05535_);
  or (_15012_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or (_15013_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  and (_15014_, _15013_, _15012_);
  and (_15015_, _15014_, _09792_);
  or (_15016_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or (_15017_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  and (_15018_, _15017_, _15016_);
  and (_15019_, _15018_, _05549_);
  or (_15020_, _15019_, _15015_);
  and (_15021_, _15020_, _09791_);
  or (_15022_, _15021_, _09805_);
  or (_15023_, _15022_, _15011_);
  and (_15024_, _15023_, _15001_);
  or (_15025_, _15024_, _05518_);
  and (_15026_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  and (_15027_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  or (_15028_, _15027_, _15026_);
  and (_15029_, _15028_, _09792_);
  and (_15030_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  and (_15031_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  or (_15032_, _15031_, _15030_);
  and (_15033_, _15032_, _05549_);
  or (_15034_, _15033_, _15029_);
  and (_15035_, _15034_, _05535_);
  and (_15036_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  and (_15037_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  or (_15038_, _15037_, _15036_);
  and (_15039_, _15038_, _09792_);
  and (_15040_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  and (_15041_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  or (_15042_, _15041_, _15040_);
  and (_15043_, _15042_, _05549_);
  or (_15044_, _15043_, _15039_);
  and (_15045_, _15044_, _09791_);
  or (_15046_, _15045_, _05542_);
  or (_15047_, _15046_, _15035_);
  or (_15048_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_15049_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  and (_15050_, _15049_, _15048_);
  and (_15051_, _15050_, _09792_);
  or (_15052_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_15053_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  and (_15054_, _15053_, _15052_);
  and (_15055_, _15054_, _05549_);
  or (_15056_, _15055_, _15051_);
  and (_15057_, _15056_, _05535_);
  or (_15058_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_15059_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  and (_15060_, _15059_, _15058_);
  and (_15061_, _15060_, _09792_);
  or (_15062_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_15063_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  and (_15064_, _15063_, _15062_);
  and (_15065_, _15064_, _05549_);
  or (_15066_, _15065_, _15061_);
  and (_15067_, _15066_, _09791_);
  or (_15068_, _15067_, _09805_);
  or (_15069_, _15068_, _15057_);
  and (_15070_, _15069_, _15047_);
  or (_15071_, _15070_, _09850_);
  and (_15072_, _15071_, _05520_);
  and (_15073_, _15072_, _15025_);
  and (_15074_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  and (_15075_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_15076_, _15075_, _15074_);
  and (_15077_, _15076_, _05549_);
  and (_15078_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  and (_15079_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_15080_, _15079_, _15078_);
  and (_15081_, _15080_, _09792_);
  or (_15082_, _15081_, _15077_);
  or (_15083_, _15082_, _09791_);
  and (_15084_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  and (_15085_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_15086_, _15085_, _15084_);
  and (_15087_, _15086_, _05549_);
  and (_15088_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  and (_15089_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_15090_, _15089_, _15088_);
  and (_15091_, _15090_, _09792_);
  or (_15092_, _15091_, _15087_);
  or (_15093_, _15092_, _05535_);
  and (_15094_, _15093_, _09805_);
  and (_15095_, _15094_, _15083_);
  or (_15096_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_15097_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  and (_15098_, _15097_, _09792_);
  and (_15099_, _15098_, _15096_);
  or (_15100_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_15101_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  and (_15102_, _15101_, _05549_);
  and (_15103_, _15102_, _15100_);
  or (_15104_, _15103_, _15099_);
  or (_15105_, _15104_, _09791_);
  or (_15106_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_15107_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  and (_15108_, _15107_, _09792_);
  and (_15109_, _15108_, _15106_);
  or (_15110_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_15111_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  and (_15112_, _15111_, _05549_);
  and (_15113_, _15112_, _15110_);
  or (_15114_, _15113_, _15109_);
  or (_15115_, _15114_, _05535_);
  and (_15116_, _15115_, _05542_);
  and (_15117_, _15116_, _15105_);
  or (_15118_, _15117_, _15095_);
  and (_15119_, _15118_, _09850_);
  and (_15120_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  and (_15121_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_15122_, _15121_, _09792_);
  or (_15123_, _15122_, _15120_);
  and (_15124_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  and (_15125_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_15126_, _15125_, _05549_);
  or (_15127_, _15126_, _15124_);
  and (_15128_, _15127_, _15123_);
  or (_15129_, _15128_, _09791_);
  and (_15130_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  and (_15131_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_15132_, _15131_, _09792_);
  or (_15133_, _15132_, _15130_);
  and (_15134_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  and (_15135_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_15136_, _15135_, _05549_);
  or (_15137_, _15136_, _15134_);
  and (_15138_, _15137_, _15133_);
  or (_15139_, _15138_, _05535_);
  and (_15140_, _15139_, _09805_);
  and (_15141_, _15140_, _15129_);
  or (_15142_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_15143_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  and (_15144_, _15143_, _15142_);
  or (_15145_, _15144_, _05549_);
  or (_15146_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_15147_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  and (_15148_, _15147_, _15146_);
  or (_15149_, _15148_, _09792_);
  and (_15150_, _15149_, _15145_);
  or (_15151_, _15150_, _09791_);
  or (_15152_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_15153_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  and (_15154_, _15153_, _15152_);
  or (_15155_, _15154_, _05549_);
  or (_15156_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_15157_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  and (_15158_, _15157_, _15156_);
  or (_15159_, _15158_, _09792_);
  and (_15160_, _15159_, _15155_);
  or (_15161_, _15160_, _05535_);
  and (_15163_, _15161_, _05542_);
  and (_15164_, _15163_, _15151_);
  or (_15165_, _15164_, _15141_);
  and (_15166_, _15165_, _05518_);
  or (_15167_, _15166_, _15119_);
  and (_15168_, _15167_, _09790_);
  or (_15169_, _15168_, _15073_);
  or (_15170_, _15169_, _10033_);
  and (_15171_, _15170_, _14979_);
  or (_15172_, _15171_, _00143_);
  and (_15173_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  and (_15174_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  or (_15175_, _15174_, _15173_);
  and (_15176_, _15175_, _09792_);
  and (_15177_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  and (_15178_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  or (_15179_, _15178_, _15177_);
  and (_15180_, _15179_, _05549_);
  or (_15181_, _15180_, _15176_);
  or (_15182_, _15181_, _09791_);
  and (_15183_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  and (_15184_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  or (_15185_, _15184_, _15183_);
  and (_15186_, _15185_, _09792_);
  and (_15187_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  and (_15188_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  or (_15189_, _15188_, _15187_);
  and (_15190_, _15189_, _05549_);
  or (_15191_, _15190_, _15186_);
  or (_15192_, _15191_, _05535_);
  and (_15193_, _15192_, _09805_);
  and (_15194_, _15193_, _15182_);
  or (_15195_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  or (_15196_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  and (_15197_, _15196_, _15195_);
  and (_15198_, _15197_, _09792_);
  or (_15199_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  or (_15200_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  and (_15201_, _15200_, _15199_);
  and (_15202_, _15201_, _05549_);
  or (_15203_, _15202_, _15198_);
  or (_15204_, _15203_, _09791_);
  or (_15205_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  or (_15206_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  and (_15207_, _15206_, _15205_);
  and (_15208_, _15207_, _09792_);
  or (_15209_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  or (_15210_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  and (_15211_, _15210_, _15209_);
  and (_15212_, _15211_, _05549_);
  or (_15214_, _15212_, _15208_);
  or (_15215_, _15214_, _05535_);
  and (_15216_, _15215_, _05542_);
  and (_15217_, _15216_, _15204_);
  or (_15218_, _15217_, _15194_);
  and (_15219_, _15218_, _05518_);
  and (_15220_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  and (_15221_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  or (_15222_, _15221_, _15220_);
  and (_15223_, _15222_, _09792_);
  and (_15224_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  and (_15225_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  or (_15226_, _15225_, _15224_);
  and (_15227_, _15226_, _05549_);
  or (_15228_, _15227_, _15223_);
  or (_15229_, _15228_, _09791_);
  and (_15230_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_15231_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  or (_15232_, _15231_, _15230_);
  and (_15233_, _15232_, _09792_);
  and (_15235_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  and (_15236_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  or (_15237_, _15236_, _15235_);
  and (_15238_, _15237_, _05549_);
  or (_15239_, _15238_, _15233_);
  or (_15240_, _15239_, _05535_);
  and (_15241_, _15240_, _09805_);
  and (_15242_, _15241_, _15229_);
  or (_15243_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  or (_15244_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_15245_, _15244_, _05549_);
  and (_15246_, _15245_, _15243_);
  or (_15247_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  or (_15248_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  and (_15249_, _15248_, _09792_);
  and (_15250_, _15249_, _15247_);
  or (_15251_, _15250_, _15246_);
  or (_15252_, _15251_, _09791_);
  or (_15253_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  or (_15254_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  and (_15255_, _15254_, _05549_);
  and (_15256_, _15255_, _15253_);
  or (_15257_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  or (_15258_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  and (_15259_, _15258_, _09792_);
  and (_15260_, _15259_, _15257_);
  or (_15261_, _15260_, _15256_);
  or (_15262_, _15261_, _05535_);
  and (_15263_, _15262_, _05542_);
  and (_15264_, _15263_, _15252_);
  or (_15265_, _15264_, _15242_);
  and (_15266_, _15265_, _09850_);
  or (_15267_, _15266_, _15219_);
  and (_15268_, _15267_, _09790_);
  and (_15269_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  and (_15270_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or (_15271_, _15270_, _15269_);
  and (_15272_, _15271_, _09792_);
  and (_15273_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  and (_15274_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or (_15275_, _15274_, _15273_);
  and (_15276_, _15275_, _05549_);
  or (_15277_, _15276_, _15272_);
  and (_15278_, _15277_, _05535_);
  and (_15279_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  and (_15280_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or (_15281_, _15280_, _15279_);
  and (_15282_, _15281_, _09792_);
  and (_15283_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  and (_15284_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or (_15285_, _15284_, _15283_);
  and (_15286_, _15285_, _05549_);
  or (_15287_, _15286_, _15282_);
  and (_15288_, _15287_, _09791_);
  or (_15289_, _15288_, _15278_);
  and (_15290_, _15289_, _09805_);
  or (_15291_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or (_15292_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  and (_15293_, _15292_, _05549_);
  and (_15294_, _15293_, _15291_);
  or (_15295_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or (_15296_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  and (_15297_, _15296_, _09792_);
  and (_15298_, _15297_, _15295_);
  or (_15299_, _15298_, _15294_);
  and (_15300_, _15299_, _05535_);
  or (_15301_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or (_15302_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  and (_15303_, _15302_, _05549_);
  and (_15304_, _15303_, _15301_);
  or (_15305_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or (_15306_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  and (_15307_, _15306_, _09792_);
  and (_15308_, _15307_, _15305_);
  or (_15309_, _15308_, _15304_);
  and (_15310_, _15309_, _09791_);
  or (_15311_, _15310_, _15300_);
  and (_15312_, _15311_, _05542_);
  or (_15313_, _15312_, _15290_);
  and (_15314_, _15313_, _09850_);
  and (_15315_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  and (_15316_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or (_15317_, _15316_, _15315_);
  and (_15318_, _15317_, _09792_);
  and (_15319_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  and (_15320_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or (_15321_, _15320_, _15319_);
  and (_15322_, _15321_, _05549_);
  or (_15323_, _15322_, _15318_);
  and (_15324_, _15323_, _05535_);
  and (_15325_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  and (_15326_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or (_15327_, _15326_, _15325_);
  and (_15328_, _15327_, _09792_);
  and (_15329_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  and (_15330_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or (_15331_, _15330_, _15329_);
  and (_15332_, _15331_, _05549_);
  or (_15333_, _15332_, _15328_);
  and (_15334_, _15333_, _09791_);
  or (_15335_, _15334_, _15324_);
  and (_15336_, _15335_, _09805_);
  or (_15337_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or (_15338_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  and (_15339_, _15338_, _15337_);
  and (_15340_, _15339_, _09792_);
  or (_15341_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  or (_15342_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  and (_15343_, _15342_, _15341_);
  and (_15344_, _15343_, _05549_);
  or (_15345_, _15344_, _15340_);
  and (_15346_, _15345_, _05535_);
  or (_15347_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  or (_15348_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  and (_15349_, _15348_, _15347_);
  and (_15350_, _15349_, _09792_);
  or (_15351_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  or (_15352_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  and (_15353_, _15352_, _15351_);
  and (_15354_, _15353_, _05549_);
  or (_15355_, _15354_, _15350_);
  and (_15356_, _15355_, _09791_);
  or (_15357_, _15356_, _15346_);
  and (_15358_, _15357_, _05542_);
  or (_15359_, _15358_, _15336_);
  and (_15360_, _15359_, _05518_);
  or (_15361_, _15360_, _15314_);
  and (_15362_, _15361_, _05520_);
  or (_15363_, _15362_, _15268_);
  or (_15364_, _15363_, _05526_);
  and (_15365_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  and (_15366_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  or (_15367_, _15366_, _15365_);
  and (_15368_, _15367_, _09792_);
  and (_15369_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  and (_15370_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_15371_, _15370_, _15369_);
  and (_15372_, _15371_, _05549_);
  or (_15373_, _15372_, _15368_);
  or (_15374_, _15373_, _09791_);
  and (_15375_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  and (_15376_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_15377_, _15376_, _15375_);
  and (_15378_, _15377_, _09792_);
  and (_15379_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  and (_15380_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  or (_15381_, _15380_, _15379_);
  and (_15382_, _15381_, _05549_);
  or (_15383_, _15382_, _15378_);
  or (_15384_, _15383_, _05535_);
  and (_15385_, _15384_, _09805_);
  and (_15386_, _15385_, _15374_);
  or (_15387_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  or (_15388_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  and (_15389_, _15388_, _05549_);
  and (_15390_, _15389_, _15387_);
  or (_15391_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_15392_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  and (_15393_, _15392_, _09792_);
  and (_15394_, _15393_, _15391_);
  or (_15395_, _15394_, _15390_);
  or (_15396_, _15395_, _09791_);
  or (_15397_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  or (_15398_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  and (_15399_, _15398_, _05549_);
  and (_15400_, _15399_, _15397_);
  or (_15401_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  or (_15402_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  and (_15403_, _15402_, _09792_);
  and (_15404_, _15403_, _15401_);
  or (_15405_, _15404_, _15400_);
  or (_15406_, _15405_, _05535_);
  and (_15407_, _15406_, _05542_);
  and (_15408_, _15407_, _15396_);
  or (_15409_, _15408_, _15386_);
  and (_15410_, _15409_, _09850_);
  and (_15411_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  and (_15412_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_15413_, _15412_, _15411_);
  and (_15414_, _15413_, _09792_);
  and (_15415_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  and (_15416_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  or (_15417_, _15416_, _15415_);
  and (_15418_, _15417_, _05549_);
  or (_15419_, _15418_, _15414_);
  or (_15420_, _15419_, _09791_);
  and (_15421_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  and (_15422_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or (_15423_, _15422_, _15421_);
  and (_15424_, _15423_, _09792_);
  and (_15425_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  and (_15426_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_15427_, _15426_, _15425_);
  and (_15428_, _15427_, _05549_);
  or (_15429_, _15428_, _15424_);
  or (_15430_, _15429_, _05535_);
  and (_15431_, _15430_, _09805_);
  and (_15432_, _15431_, _15420_);
  or (_15433_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  or (_15434_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  and (_15435_, _15434_, _15433_);
  and (_15436_, _15435_, _09792_);
  or (_15437_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  or (_15438_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  and (_15439_, _15438_, _15437_);
  and (_15440_, _15439_, _05549_);
  or (_15441_, _15440_, _15436_);
  or (_15442_, _15441_, _09791_);
  or (_15443_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  or (_15444_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  and (_15445_, _15444_, _15443_);
  and (_15446_, _15445_, _09792_);
  or (_15447_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_15448_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  and (_15449_, _15448_, _15447_);
  and (_15450_, _15449_, _05549_);
  or (_15451_, _15450_, _15446_);
  or (_15452_, _15451_, _05535_);
  and (_15453_, _15452_, _05542_);
  and (_15454_, _15453_, _15442_);
  or (_15455_, _15454_, _15432_);
  and (_15456_, _15455_, _05518_);
  or (_15457_, _15456_, _15410_);
  and (_15458_, _15457_, _09790_);
  or (_15459_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  or (_15460_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  and (_15461_, _15460_, _15459_);
  and (_15462_, _15461_, _09792_);
  or (_15463_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  or (_15464_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  and (_15465_, _15464_, _15463_);
  and (_15466_, _15465_, _05549_);
  or (_15467_, _15466_, _15462_);
  and (_15468_, _15467_, _09791_);
  or (_15469_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  or (_15470_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  and (_15471_, _15470_, _15469_);
  and (_15472_, _15471_, _09792_);
  or (_15473_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  or (_15474_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  and (_15475_, _15474_, _15473_);
  and (_15476_, _15475_, _05549_);
  or (_15477_, _15476_, _15472_);
  and (_15478_, _15477_, _05535_);
  or (_15479_, _15478_, _15468_);
  and (_15480_, _15479_, _05542_);
  and (_15481_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  and (_15482_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  or (_15483_, _15482_, _15481_);
  and (_15484_, _15483_, _09792_);
  and (_15485_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  and (_15486_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  or (_15487_, _15486_, _15485_);
  and (_15488_, _15487_, _05549_);
  or (_15489_, _15488_, _15484_);
  and (_15490_, _15489_, _09791_);
  and (_15491_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  and (_15492_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  or (_15493_, _15492_, _15491_);
  and (_15494_, _15493_, _09792_);
  and (_15495_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  and (_15496_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  or (_15497_, _15496_, _15495_);
  and (_15498_, _15497_, _05549_);
  or (_15499_, _15498_, _15494_);
  and (_15500_, _15499_, _05535_);
  or (_15501_, _15500_, _15490_);
  and (_15502_, _15501_, _09805_);
  or (_15503_, _15502_, _15480_);
  and (_15504_, _15503_, _05518_);
  or (_15505_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_15506_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  and (_15507_, _15506_, _05549_);
  and (_15508_, _15507_, _15505_);
  or (_15509_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_15510_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  and (_15511_, _15510_, _09792_);
  and (_15512_, _15511_, _15509_);
  or (_15513_, _15512_, _15508_);
  and (_15514_, _15513_, _09791_);
  or (_15515_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  or (_15516_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  and (_15517_, _15516_, _05549_);
  and (_15518_, _15517_, _15515_);
  or (_15519_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  or (_15520_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  and (_15521_, _15520_, _09792_);
  and (_15522_, _15521_, _15519_);
  or (_15523_, _15522_, _15518_);
  and (_15524_, _15523_, _05535_);
  or (_15525_, _15524_, _15514_);
  and (_15526_, _15525_, _05542_);
  and (_15527_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  and (_15528_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  or (_15529_, _15528_, _15527_);
  and (_15530_, _15529_, _09792_);
  and (_15531_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  and (_15532_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  or (_15533_, _15532_, _15531_);
  and (_15534_, _15533_, _05549_);
  or (_15535_, _15534_, _15530_);
  and (_15536_, _15535_, _09791_);
  and (_15537_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  and (_15538_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  or (_15539_, _15538_, _15537_);
  and (_15540_, _15539_, _09792_);
  and (_15541_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  and (_15542_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  or (_15543_, _15542_, _15541_);
  and (_15544_, _15543_, _05549_);
  or (_15545_, _15544_, _15540_);
  and (_15546_, _15545_, _05535_);
  or (_15547_, _15546_, _15536_);
  and (_15548_, _15547_, _09805_);
  or (_15549_, _15548_, _15526_);
  and (_15550_, _15549_, _09850_);
  or (_15551_, _15550_, _15504_);
  and (_15552_, _15551_, _05520_);
  or (_15553_, _15552_, _15458_);
  or (_15554_, _15553_, _10033_);
  and (_15555_, _15554_, _15364_);
  or (_15556_, _15555_, _04413_);
  and (_15557_, _15556_, _15172_);
  or (_15558_, _15557_, _05563_);
  or (_15559_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_15560_, _15559_, _22731_);
  and (_04805_, _15560_, _15558_);
  and (_15561_, _24496_, _22974_);
  and (_15562_, _15561_, _23996_);
  not (_15563_, _15561_);
  and (_15564_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_04811_, _15564_, _15562_);
  and (_15565_, _24451_, _24089_);
  and (_15566_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  or (_04814_, _15566_, _15565_);
  and (_15567_, _09779_, _24474_);
  and (_15568_, _15567_, _23583_);
  not (_15569_, _15567_);
  and (_15570_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  or (_04817_, _15570_, _15568_);
  and (_15571_, _14778_, _23996_);
  and (_15572_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  or (_04822_, _15572_, _15571_);
  and (_15573_, _15567_, _24051_);
  and (_15574_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  or (_26992_, _15574_, _15573_);
  and (_15575_, _14778_, _24134_);
  and (_15576_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  or (_04834_, _15576_, _15575_);
  and (_15577_, _14778_, _24051_);
  and (_15578_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  or (_04836_, _15578_, _15577_);
  and (_15579_, _15561_, _24134_);
  and (_15580_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  or (_04839_, _15580_, _15579_);
  and (_15581_, _24365_, _24159_);
  and (_15582_, _15581_, _24051_);
  not (_15583_, _15581_);
  and (_15584_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  or (_04842_, _15584_, _15582_);
  and (_15585_, _15567_, _24089_);
  and (_15586_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  or (_04845_, _15586_, _15585_);
  and (_15587_, _08435_, _24051_);
  and (_15588_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  or (_04850_, _15588_, _15587_);
  and (_15589_, _14778_, _24219_);
  and (_15590_, _14780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  or (_04857_, _15590_, _15589_);
  and (_15591_, _03236_, _24051_);
  and (_15592_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  or (_04863_, _15592_, _15591_);
  and (_15593_, _08523_, _23583_);
  and (_15594_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  or (_04870_, _15594_, _15593_);
  and (_15595_, _10746_, _24134_);
  and (_15596_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  or (_04873_, _15596_, _15595_);
  and (_15597_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  and (_15598_, _03221_, _24219_);
  or (_04883_, _15598_, _15597_);
  and (_15599_, _15561_, _24051_);
  and (_15600_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  or (_04889_, _15600_, _15599_);
  and (_15601_, _03320_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  and (_15602_, _03319_, _24051_);
  or (_04906_, _15602_, _15601_);
  and (_15603_, _03222_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  and (_15604_, _03221_, _23996_);
  or (_27093_, _15604_, _15603_);
  and (_15605_, _24899_, _24476_);
  and (_15606_, _15605_, _24089_);
  not (_15607_, _15605_);
  and (_15608_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  or (_04911_, _15608_, _15606_);
  and (_15609_, _10746_, _23996_);
  and (_15610_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  or (_04914_, _15610_, _15609_);
  and (_15611_, _15567_, _23996_);
  and (_15612_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_04917_, _15612_, _15611_);
  and (_15613_, _15605_, _23583_);
  and (_15614_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  or (_04919_, _15614_, _15613_);
  and (_15615_, _15605_, _23887_);
  and (_15616_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  or (_04922_, _15616_, _15615_);
  and (_15617_, _15567_, _24134_);
  and (_15618_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  or (_04927_, _15618_, _15617_);
  and (_15620_, _02432_, _23583_);
  and (_15621_, _02434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  or (_04929_, _15621_, _15620_);
  and (_15622_, _03370_, _23548_);
  and (_15623_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  or (_04931_, _15623_, _15622_);
  and (_15624_, _03370_, _23583_);
  and (_15625_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  or (_04934_, _15625_, _15624_);
  and (_15626_, _04865_, _23548_);
  and (_15627_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  or (_26963_, _15627_, _15626_);
  and (_15628_, _15605_, _23996_);
  and (_15629_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  or (_27181_, _15629_, _15628_);
  and (_15630_, _03236_, _23583_);
  and (_15631_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  or (_04954_, _15631_, _15630_);
  and (_15632_, _03236_, _24219_);
  and (_15633_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_04958_, _15633_, _15632_);
  and (_15634_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  and (_15635_, _04614_, _23548_);
  or (_04960_, _15635_, _15634_);
  and (_15636_, _03236_, _23548_);
  and (_15637_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  or (_04962_, _15637_, _15636_);
  and (_15638_, _15605_, _24134_);
  and (_15639_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  or (_04963_, _15639_, _15638_);
  and (_15640_, _09779_, _24056_);
  and (_15641_, _15640_, _23996_);
  not (_15642_, _15640_);
  and (_15643_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  or (_04966_, _15643_, _15641_);
  and (_15644_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_15645_, _03662_, _24219_);
  or (_04968_, _15645_, _15644_);
  and (_15646_, _15605_, _24051_);
  and (_15647_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  or (_27180_, _15647_, _15646_);
  and (_15648_, _04615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  and (_15649_, _04614_, _24051_);
  or (_04972_, _15649_, _15648_);
  and (_15650_, _15640_, _24134_);
  and (_15651_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  or (_26988_, _15651_, _15650_);
  and (_15652_, _03663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and (_15653_, _03662_, _23996_);
  or (_27096_, _15653_, _15652_);
  and (_15654_, _03236_, _23887_);
  and (_15655_, _03238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  or (_05005_, _15655_, _15654_);
  and (_15656_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  not (_15657_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_15658_, _02248_, _02237_);
  and (_15659_, _15658_, _02264_);
  not (_15660_, _02237_);
  and (_15661_, _02248_, _02236_);
  and (_15662_, _15661_, _15660_);
  and (_15663_, _15662_, _02272_);
  nor (_15664_, _15663_, _15659_);
  nand (_15665_, _15664_, _15657_);
  or (_15666_, _15664_, _15657_);
  nand (_15667_, _15666_, _15665_);
  nor (_15668_, _15667_, _02292_);
  and (_15669_, _02292_, _23880_);
  or (_15670_, _15669_, _15668_);
  and (_15671_, _15670_, _02295_);
  or (_05019_, _15671_, _15656_);
  and (_15672_, _24478_, _24134_);
  and (_15673_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  or (_05024_, _15673_, _15672_);
  and (_15674_, _08435_, _24089_);
  and (_15675_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  or (_05027_, _15675_, _15674_);
  and (_15676_, _24478_, _24051_);
  and (_15677_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  or (_05029_, _15677_, _15676_);
  and (_15678_, _03370_, _23996_);
  and (_15679_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_05052_, _15679_, _15678_);
  and (_15680_, _15567_, _23548_);
  and (_15681_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  or (_26990_, _15681_, _15680_);
  and (_15682_, _15567_, _24219_);
  and (_15683_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or (_26989_, _15683_, _15682_);
  and (_15684_, _15605_, _24219_);
  and (_15685_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  or (_05064_, _15685_, _15684_);
  and (_15686_, _10746_, _24051_);
  and (_15687_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  or (_05089_, _15687_, _15686_);
  and (_15688_, _24320_, _23548_);
  and (_15689_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  or (_05091_, _15689_, _15688_);
  and (_15690_, _24478_, _23996_);
  and (_15691_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_05093_, _15691_, _15690_);
  and (_15692_, _10746_, _23583_);
  and (_15693_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  or (_05113_, _15693_, _15692_);
  and (_15694_, _24142_, _23583_);
  and (_15695_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  or (_05116_, _15695_, _15694_);
  and (_15696_, _07038_, _24051_);
  and (_15697_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  or (_05135_, _15697_, _15696_);
  and (_15698_, _12429_, _23583_);
  and (_15699_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  or (_05143_, _15699_, _15698_);
  and (_15700_, _10746_, _24089_);
  and (_15701_, _10749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  or (_27116_, _15701_, _15700_);
  and (_15702_, _12429_, _23887_);
  and (_15703_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  or (_27184_, _15703_, _15702_);
  and (_15704_, _12429_, _23548_);
  and (_15705_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  or (_27183_, _15705_, _15704_);
  and (_15706_, _04654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  and (_15707_, _04653_, _23548_);
  or (_05154_, _15707_, _15706_);
  and (_15708_, _24319_, _24141_);
  and (_15709_, _15708_, _24051_);
  not (_15710_, _15708_);
  and (_15711_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  or (_05163_, _15711_, _15709_);
  and (_15712_, _15640_, _24219_);
  and (_15713_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  or (_05166_, _15713_, _15712_);
  and (_15714_, _03370_, _24089_);
  and (_15715_, _03372_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  or (_05168_, _15715_, _15714_);
  and (_15716_, _09779_, _24223_);
  and (_15717_, _15716_, _23996_);
  not (_15718_, _15716_);
  and (_15719_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or (_05172_, _15719_, _15717_);
  and (_15720_, _15708_, _23887_);
  and (_15721_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  or (_05175_, _15721_, _15720_);
  and (_15722_, _12429_, _24051_);
  and (_15723_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  or (_05187_, _15723_, _15722_);
  and (_15724_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  and (_15725_, _09705_, _24051_);
  or (_05189_, _15725_, _15724_);
  and (_15726_, _12429_, _24089_);
  and (_15727_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  or (_05206_, _15727_, _15726_);
  and (_15728_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  and (_15729_, _09705_, _23548_);
  or (_27023_, _15729_, _15728_);
  and (_15730_, _08523_, _23887_);
  and (_15731_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  or (_05217_, _15731_, _15730_);
  and (_15732_, _15640_, _23583_);
  and (_15733_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  or (_05220_, _15733_, _15732_);
  and (_15734_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  and (_15735_, _09676_, _24134_);
  or (_05222_, _15735_, _15734_);
  and (_15736_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_15737_, _09676_, _24219_);
  or (_05238_, _15737_, _15736_);
  and (_15738_, _15640_, _23887_);
  and (_15739_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  or (_05241_, _15739_, _15738_);
  and (_15740_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  and (_15741_, _09645_, _24051_);
  or (_05245_, _15741_, _15740_);
  and (_15742_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  and (_15743_, _09645_, _23548_);
  or (_05252_, _15743_, _15742_);
  and (_15744_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  and (_15745_, _08591_, _24134_);
  or (_05272_, _15745_, _15744_);
  and (_15746_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  and (_15747_, _08591_, _23583_);
  or (_27017_, _15747_, _15746_);
  and (_15748_, _15708_, _23583_);
  and (_15749_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  or (_26926_, _15749_, _15748_);
  and (_15750_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  and (_15751_, _06339_, _24089_);
  or (_05283_, _15751_, _15750_);
  and (_15752_, _24889_, _23548_);
  and (_15753_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  or (_05290_, _15753_, _15752_);
  and (_15754_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  and (_15755_, _06339_, _23548_);
  or (_27014_, _15755_, _15754_);
  and (_15756_, _15716_, _23887_);
  and (_15757_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  or (_05320_, _15757_, _15756_);
  and (_15758_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  and (_15759_, _05596_, _24134_);
  or (_05325_, _15759_, _15758_);
  and (_15760_, _07779_, _24089_);
  and (_15761_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  or (_05330_, _15761_, _15760_);
  and (_15762_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  and (_15763_, _05596_, _23548_);
  or (_05336_, _15763_, _15762_);
  and (_15764_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_15765_, _05580_, _23996_);
  or (_05346_, _15765_, _15764_);
  and (_15766_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  and (_15767_, _05580_, _23887_);
  or (_05354_, _15767_, _15766_);
  and (_15768_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  and (_15769_, _05567_, _23996_);
  or (_05357_, _15769_, _15768_);
  and (_15770_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  and (_15771_, _05567_, _23887_);
  or (_05369_, _15771_, _15770_);
  and (_15772_, _15708_, _23996_);
  and (_15773_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_05379_, _15773_, _15772_);
  and (_15774_, _09774_, _23548_);
  and (_15775_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  or (_05383_, _15775_, _15774_);
  and (_15776_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  and (_15777_, _04937_, _23583_);
  or (_05390_, _15777_, _15776_);
  and (_15778_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  and (_15779_, _04905_, _24089_);
  or (_05423_, _15779_, _15778_);
  and (_15780_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_15781_, _04905_, _24219_);
  or (_05433_, _15781_, _15780_);
  and (_15782_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  and (_15783_, _04897_, _24051_);
  or (_05445_, _15783_, _15782_);
  and (_15784_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  and (_15785_, _04879_, _24134_);
  or (_05447_, _15785_, _15784_);
  and (_15786_, _09774_, _24219_);
  and (_15787_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  or (_05450_, _15787_, _15786_);
  and (_15788_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  and (_15789_, _04879_, _23583_);
  or (_05452_, _15789_, _15788_);
  and (_15790_, _09670_, _23548_);
  and (_15791_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  or (_27203_, _15791_, _15790_);
  and (_15792_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_15793_, _05580_, _24219_);
  or (_27013_, _15793_, _15792_);
  nand (_15794_, _25025_, _24004_);
  or (_15795_, _15794_, _00883_);
  nand (_15796_, _15794_, _04308_);
  and (_15797_, _15796_, _24179_);
  and (_15798_, _15797_, _15795_);
  nor (_15799_, _24178_, _04308_);
  and (_15800_, _00327_, _25017_);
  and (_15801_, _15800_, _25481_);
  nand (_15802_, _15801_, _23504_);
  or (_15803_, _15801_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_15804_, _15803_, _24539_);
  and (_15805_, _15804_, _15802_);
  or (_15806_, _15805_, _15799_);
  or (_15807_, _15806_, _15798_);
  and (_05463_, _15807_, _22731_);
  and (_15808_, _02837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  and (_15809_, _02836_, _24219_);
  or (_05466_, _15809_, _15808_);
  and (_15810_, _07038_, _24089_);
  and (_15811_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  or (_05470_, _15811_, _15810_);
  and (_15812_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  and (_15813_, _09676_, _23887_);
  or (_05474_, _15813_, _15812_);
  and (_15814_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  not (_15815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_15816_, _11153_, _15815_);
  and (_15817_, _11153_, _15815_);
  nor (_15818_, _15817_, _15816_);
  nor (_15819_, _15818_, _02292_);
  and (_15820_, _02292_, _02728_);
  or (_15821_, _15820_, _15819_);
  and (_15822_, _15821_, _02295_);
  or (_05476_, _15822_, _15814_);
  or (_15823_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_15824_, _15823_, _22731_);
  or (_15825_, _11256_, _23577_);
  and (_05477_, _15825_, _15824_);
  and (_15826_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  and (_15827_, _09645_, _23996_);
  or (_05483_, _15827_, _15826_);
  and (_15828_, _09646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  and (_15829_, _09645_, _23583_);
  or (_05503_, _15829_, _15828_);
  and (_15830_, _24223_, _24141_);
  and (_15831_, _15830_, _24219_);
  not (_15832_, _15830_);
  and (_15833_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_26928_, _15833_, _15831_);
  and (_15834_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  and (_15835_, _08591_, _24219_);
  or (_27016_, _15835_, _15834_);
  and (_15836_, _05597_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  and (_15837_, _05596_, _23583_);
  or (_05557_, _15837_, _15836_);
  and (_15838_, _05582_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  and (_15839_, _05580_, _24089_);
  or (_05564_, _15839_, _15838_);
  and (_15840_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  and (_15841_, _05567_, _24089_);
  or (_05575_, _15841_, _15840_);
  and (_15842_, _05568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  and (_15843_, _05567_, _24219_);
  or (_05581_, _15843_, _15842_);
  and (_15844_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  and (_15845_, _04937_, _24051_);
  or (_05586_, _15845_, _15844_);
  and (_15846_, _04938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  and (_15847_, _04937_, _23548_);
  or (_05588_, _15847_, _15846_);
  and (_15848_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  and (_15849_, _04905_, _24134_);
  or (_05590_, _15849_, _15848_);
  and (_15850_, _04907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  and (_15851_, _04905_, _23887_);
  or (_27011_, _15851_, _15850_);
  and (_15852_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_15853_, _04897_, _23996_);
  or (_27009_, _15853_, _15852_);
  or (_15854_, _11099_, _23880_);
  and (_15855_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_15856_, _02256_, _02248_);
  or (_15857_, _15856_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_15858_, _11102_, _02281_);
  and (_15859_, _15858_, _15857_);
  and (_15860_, _02623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_15861_, _15860_, _15859_);
  nor (_15862_, _15861_, _02616_);
  nor (_15863_, _15862_, _15855_);
  nand (_15864_, _15863_, _11099_);
  and (_15865_, _15864_, _22731_);
  and (_05602_, _15865_, _15854_);
  and (_15866_, _09706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  and (_15867_, _09705_, _23887_);
  or (_05607_, _15867_, _15866_);
  and (_15868_, _08592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  and (_15869_, _08591_, _24089_);
  or (_05644_, _15869_, _15868_);
  and (_15870_, _08435_, _23996_);
  and (_15871_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  or (_05648_, _15871_, _15870_);
  and (_15872_, _06341_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  and (_15873_, _06339_, _24051_);
  or (_05650_, _15873_, _15872_);
  and (_15874_, _06154_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_15875_, _11134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_15876_, _15856_, _02281_);
  and (_15877_, _15876_, _15875_);
  and (_15878_, _02623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_15879_, _15878_, _15877_);
  nor (_15880_, _15879_, _02616_);
  or (_15881_, _15880_, _15874_);
  and (_15882_, _15881_, _02295_);
  and (_15883_, _02440_, _02728_);
  or (_05666_, _15883_, _15882_);
  and (_15884_, _03355_, _24051_);
  and (_15885_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  or (_05676_, _15885_, _15884_);
  and (_15886_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_15887_, _04879_, _23996_);
  or (_05695_, _15887_, _15886_);
  and (_15888_, _24496_, _24095_);
  and (_15889_, _15888_, _23996_);
  not (_15890_, _15888_);
  and (_15891_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_05703_, _15891_, _15889_);
  and (_15892_, _09677_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  and (_15893_, _09676_, _23583_);
  or (_05714_, _15893_, _15892_);
  and (_15894_, _15716_, _23548_);
  and (_15895_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  or (_05718_, _15895_, _15894_);
  and (_15896_, _15830_, _23548_);
  and (_15897_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  or (_26929_, _15897_, _15896_);
  and (_15898_, _04880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_15899_, _04879_, _24219_);
  or (_05729_, _15899_, _15898_);
  and (_15900_, _15716_, _24219_);
  and (_15901_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or (_05740_, _15901_, _15900_);
  and (_15902_, _09780_, _24051_);
  and (_15903_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  or (_05778_, _15903_, _15902_);
  and (_15904_, _10797_, _23548_);
  and (_15905_, _10799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  or (_05781_, _15905_, _15904_);
  and (_15906_, _15888_, _24134_);
  and (_15907_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  or (_05783_, _15907_, _15906_);
  and (_15908_, _10906_, _23583_);
  and (_15909_, _10908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  or (_05786_, _15909_, _15908_);
  and (_15910_, _15716_, _24051_);
  and (_15911_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  or (_05788_, _15911_, _15910_);
  and (_15912_, _25319_, _24533_);
  nand (_15913_, _15912_, _23504_);
  or (_15914_, _15912_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_15915_, _15914_, _24539_);
  and (_15916_, _15915_, _15913_);
  or (_15917_, _25328_, _23577_);
  or (_15918_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_15919_, _15918_, _24179_);
  and (_15920_, _15919_, _15917_);
  nor (_15921_, _24178_, _03939_);
  or (_15922_, _15921_, rst);
  or (_15923_, _15922_, _15920_);
  or (_05791_, _15923_, _15916_);
  and (_15924_, _15716_, _24089_);
  and (_15925_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  or (_05794_, _15925_, _15924_);
  and (_15926_, _12372_, _24134_);
  and (_15927_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  or (_26997_, _15927_, _15926_);
  and (_15928_, _12372_, _24219_);
  and (_15929_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  or (_26995_, _15929_, _15928_);
  and (_15930_, _25220_, _24636_);
  nand (_15931_, _15930_, _23504_);
  or (_15932_, _15930_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_15933_, _15932_, _24539_);
  and (_15934_, _15933_, _15931_);
  nand (_15935_, _25228_, _24082_);
  or (_15936_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_15937_, _15936_, _24179_);
  and (_15938_, _15937_, _15935_);
  nor (_15939_, _24178_, _03985_);
  or (_15940_, _15939_, rst);
  or (_15941_, _15940_, _15938_);
  or (_05805_, _15941_, _15934_);
  and (_15942_, _15640_, _24089_);
  and (_15943_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  or (_05812_, _15943_, _15942_);
  and (_15944_, _25124_, _24594_);
  nand (_15945_, _15944_, _23504_);
  or (_15946_, _15944_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_15947_, _15946_, _24539_);
  and (_15948_, _15947_, _15945_);
  nand (_15949_, _25130_, _24126_);
  or (_15950_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_15951_, _15950_, _24179_);
  and (_15952_, _15951_, _15949_);
  nor (_15953_, _24178_, _04230_);
  or (_15954_, _15953_, rst);
  or (_15955_, _15954_, _15952_);
  or (_05816_, _15955_, _15948_);
  and (_15956_, _09779_, _24319_);
  and (_15957_, _15956_, _23887_);
  not (_15958_, _15956_);
  and (_15959_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  or (_05820_, _15959_, _15957_);
  and (_15960_, _09779_, _22974_);
  and (_15961_, _15960_, _24089_);
  not (_15962_, _15960_);
  and (_15963_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  or (_05825_, _15963_, _15961_);
  and (_15964_, _15956_, _24089_);
  and (_15965_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  or (_05833_, _15965_, _15964_);
  and (_15966_, _15956_, _23583_);
  and (_15967_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  or (_05840_, _15967_, _15966_);
  and (_15968_, _25018_, _24636_);
  nand (_15969_, _15968_, _23504_);
  or (_15970_, _15968_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_15971_, _15970_, _24539_);
  and (_15972_, _15971_, _15969_);
  nand (_15973_, _25026_, _24082_);
  or (_15974_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_15975_, _15974_, _24179_);
  and (_15976_, _15975_, _15973_);
  nor (_15977_, _24178_, _04134_);
  or (_15978_, _15977_, rst);
  or (_15979_, _15978_, _15976_);
  or (_05843_, _15979_, _15972_);
  and (_15980_, _03308_, _24159_);
  and (_15981_, _15980_, _23583_);
  not (_15982_, _15980_);
  and (_15983_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  or (_26976_, _15983_, _15981_);
  and (_15984_, _03308_, _24297_);
  and (_15985_, _15984_, _24051_);
  not (_15986_, _15984_);
  and (_15987_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  or (_26975_, _15987_, _15985_);
  and (_15988_, _03308_, _24016_);
  and (_15989_, _15988_, _23996_);
  not (_15990_, _15988_);
  and (_15991_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or (_05859_, _15991_, _15989_);
  and (_15992_, _03308_, _24236_);
  and (_15993_, _15992_, _23887_);
  not (_15994_, _15992_);
  and (_15995_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  or (_05866_, _15995_, _15993_);
  and (_15996_, _24141_, _24016_);
  and (_15997_, _15996_, _24219_);
  not (_15998_, _15996_);
  and (_15999_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  or (_05892_, _15999_, _15997_);
  and (_16000_, _03308_, _23941_);
  and (_16001_, _16000_, _23887_);
  not (_16002_, _16000_);
  and (_16003_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  or (_05909_, _16003_, _16001_);
  and (_16004_, _03308_, _24474_);
  and (_16005_, _16004_, _23996_);
  not (_16006_, _16004_);
  and (_16007_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  or (_05913_, _16007_, _16005_);
  and (_16008_, _03308_, _24319_);
  and (_16009_, _16008_, _24051_);
  not (_16010_, _16008_);
  and (_16011_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  or (_05917_, _16011_, _16009_);
  and (_16012_, _15956_, _24134_);
  and (_16013_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  or (_05928_, _16013_, _16012_);
  and (_16014_, _03308_, _24095_);
  and (_16015_, _16014_, _23583_);
  not (_16016_, _16014_);
  and (_16017_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  or (_05932_, _16017_, _16015_);
  and (_16018_, _11441_, _23996_);
  and (_16019_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or (_05935_, _16019_, _16018_);
  and (_16020_, _03308_, _24146_);
  and (_16021_, _16020_, _24134_);
  not (_16022_, _16020_);
  and (_16023_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  or (_26950_, _16023_, _16021_);
  and (_16024_, _16020_, _23887_);
  and (_16025_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  or (_05945_, _16025_, _16024_);
  and (_16026_, _03308_, _24140_);
  and (_16027_, _16026_, _23887_);
  not (_16028_, _16026_);
  and (_16029_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  or (_05951_, _16029_, _16027_);
  and (_16030_, _03355_, _24134_);
  and (_16031_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  or (_05954_, _16031_, _16030_);
  and (_16032_, _03355_, _23887_);
  and (_16033_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  or (_05960_, _16033_, _16032_);
  and (_16034_, _24297_, _24141_);
  and (_16035_, _16034_, _24051_);
  not (_16036_, _16034_);
  and (_16037_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  or (_05974_, _16037_, _16035_);
  and (_16038_, _15830_, _23583_);
  and (_16039_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  or (_05978_, _16039_, _16038_);
  and (_16040_, _15996_, _23887_);
  and (_16041_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  or (_05981_, _16041_, _16040_);
  and (_16042_, _15960_, _23996_);
  and (_16043_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  or (_05998_, _16043_, _16042_);
  and (_16044_, _15960_, _24134_);
  and (_16045_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  or (_06021_, _16045_, _16044_);
  and (_16046_, _11046_, _24051_);
  and (_16047_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  or (_27000_, _16047_, _16046_);
  and (_16048_, _24372_, _24141_);
  and (_16049_, _16048_, _24219_);
  not (_16050_, _16048_);
  and (_16051_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_06045_, _16051_, _16049_);
  and (_16052_, _12442_, _23548_);
  and (_16053_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  or (_26993_, _16053_, _16052_);
  and (_16054_, _16048_, _23887_);
  and (_16055_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  or (_06054_, _16055_, _16054_);
  and (_16056_, _15956_, _23548_);
  and (_16057_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  or (_06059_, _16057_, _16056_);
  and (_16058_, _16048_, _23583_);
  and (_16059_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  or (_06065_, _16059_, _16058_);
  and (_16060_, _09779_, _24146_);
  and (_16061_, _16060_, _23548_);
  not (_16062_, _16060_);
  and (_16063_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  or (_06068_, _16063_, _16061_);
  and (_16064_, _25658_, _23996_);
  and (_16065_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_06071_, _16065_, _16064_);
  and (_16066_, _03308_, _22974_);
  and (_16067_, _16066_, _23887_);
  not (_16068_, _16066_);
  and (_16069_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  or (_06086_, _16069_, _16067_);
  and (_16070_, _06208_, _24219_);
  and (_16071_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_06088_, _16071_, _16070_);
  and (_16072_, _03308_, _24372_);
  and (_16073_, _16072_, _23996_);
  not (_16074_, _16072_);
  and (_16075_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  or (_26956_, _16075_, _16073_);
  and (_16076_, _16026_, _23996_);
  and (_16077_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or (_06095_, _16077_, _16076_);
  and (_16078_, _15960_, _23548_);
  and (_16079_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  or (_06107_, _16079_, _16078_);
  and (_16080_, _15996_, _24134_);
  and (_16081_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  or (_26947_, _16081_, _16080_);
  and (_16082_, _04865_, _24089_);
  and (_16083_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  or (_26965_, _16083_, _16082_);
  and (_16084_, _03309_, _24051_);
  and (_16085_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  or (_06120_, _16085_, _16084_);
  and (_16086_, _15960_, _24219_);
  and (_16087_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  or (_06123_, _16087_, _16086_);
  and (_16088_, _12372_, _23996_);
  and (_16089_, _12374_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  or (_06147_, _16089_, _16088_);
  and (_16090_, _15640_, _24051_);
  and (_16091_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  or (_06149_, _16091_, _16090_);
  and (_16092_, _15960_, _24051_);
  and (_16093_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  or (_06151_, _16093_, _16092_);
  and (_16094_, _02438_, _24607_);
  nand (_16095_, _16094_, _24043_);
  not (_16096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_16097_, _15658_, _02265_);
  and (_16098_, _15662_, _02273_);
  or (_16099_, _16098_, _16097_);
  and (_16100_, _16099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_16101_, _16100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_16102_, _16101_, _16096_);
  and (_16103_, _16101_, _16096_);
  or (_16104_, _16103_, _16102_);
  or (_16105_, _16104_, _02616_);
  and (_16106_, _16105_, _02295_);
  and (_16107_, _16106_, _16095_);
  and (_16108_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_06161_, _16108_, _16107_);
  and (_16109_, _25414_, _23583_);
  and (_16110_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  or (_27159_, _16110_, _16109_);
  and (_16111_, _03308_, _24349_);
  and (_16112_, _16111_, _24219_);
  not (_16113_, _16111_);
  and (_16114_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  or (_06169_, _16114_, _16112_);
  and (_16115_, _16008_, _24134_);
  and (_16116_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  or (_06179_, _16116_, _16115_);
  and (_16117_, _15960_, _23583_);
  and (_16118_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  or (_26985_, _16118_, _16117_);
  and (_16119_, _15960_, _23887_);
  and (_16120_, _15962_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  or (_26984_, _16120_, _16119_);
  and (_16121_, _24319_, _24301_);
  and (_16122_, _16121_, _23996_);
  not (_16123_, _16121_);
  and (_16124_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_06207_, _16124_, _16122_);
  and (_16125_, _16004_, _23548_);
  and (_16126_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  or (_06214_, _16126_, _16125_);
  and (_16127_, _16004_, _24219_);
  and (_16128_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  or (_06225_, _16128_, _16127_);
  and (_16129_, _03309_, _23548_);
  and (_16130_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  or (_06229_, _16130_, _16129_);
  and (_16131_, _03309_, _24089_);
  and (_16132_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  or (_06232_, _16132_, _16131_);
  and (_16133_, _24134_, _24017_);
  and (_16134_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  or (_06239_, _16134_, _16133_);
  and (_16135_, _03309_, _24134_);
  and (_16136_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  or (_06243_, _16136_, _16135_);
  and (_16137_, _09779_, _24095_);
  and (_16138_, _16137_, _23583_);
  not (_16139_, _16137_);
  and (_16140_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  or (_26983_, _16140_, _16138_);
  and (_16141_, _16137_, _23887_);
  and (_16142_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  or (_06248_, _16142_, _16141_);
  and (_16143_, _04865_, _23583_);
  and (_16144_, _04867_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  or (_26964_, _16144_, _16143_);
  and (_16145_, _16137_, _23548_);
  and (_16146_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  or (_06266_, _16146_, _16145_);
  and (_16147_, _06208_, _23548_);
  and (_16148_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  or (_06268_, _16148_, _16147_);
  and (_16149_, _15996_, _23548_);
  and (_16150_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  or (_06275_, _16150_, _16149_);
  and (_16151_, _15996_, _24051_);
  and (_16152_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  or (_06277_, _16152_, _16151_);
  and (_16153_, _16137_, _24219_);
  and (_16154_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  or (_06280_, _16154_, _16153_);
  and (_16155_, _15996_, _24089_);
  and (_16156_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  or (_06282_, _16156_, _16155_);
  and (_16157_, _16034_, _23548_);
  and (_16158_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  or (_06285_, _16158_, _16157_);
  and (_16159_, _16034_, _23583_);
  and (_16160_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  or (_06288_, _16160_, _16159_);
  and (_16161_, _16026_, _24134_);
  and (_16162_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  or (_06297_, _16162_, _16161_);
  and (_16163_, _16020_, _24089_);
  and (_16164_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  or (_06309_, _16164_, _16163_);
  and (_16165_, _16072_, _23887_);
  and (_16166_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  or (_26955_, _16166_, _16165_);
  and (_16167_, _16137_, _24134_);
  and (_16168_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  or (_06314_, _16168_, _16167_);
  and (_16169_, _16137_, _24051_);
  and (_16170_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  or (_06327_, _16170_, _16169_);
  and (_16171_, _16137_, _24089_);
  and (_16172_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  or (_06333_, _16172_, _16171_);
  and (_16173_, _16014_, _23548_);
  and (_16174_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  or (_06336_, _16174_, _16173_);
  and (_16175_, _24302_, _23887_);
  and (_16176_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  or (_06338_, _16176_, _16175_);
  and (_16177_, _16066_, _23548_);
  and (_16178_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  or (_06340_, _16178_, _16177_);
  and (_16179_, _16066_, _24051_);
  and (_16180_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  or (_06346_, _16180_, _16179_);
  and (_16181_, _24219_, _24017_);
  and (_16182_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  or (_06349_, _16182_, _16181_);
  and (_16183_, _16008_, _23887_);
  and (_16184_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  or (_06350_, _16184_, _16183_);
  and (_16185_, _03308_, _24899_);
  and (_16186_, _16185_, _24051_);
  not (_16187_, _16185_);
  and (_16188_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  or (_06355_, _16188_, _16186_);
  and (_16189_, _16000_, _23996_);
  and (_16190_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or (_06373_, _16190_, _16189_);
  and (_16191_, _09779_, _24372_);
  and (_16192_, _16191_, _23548_);
  not (_16193_, _16191_);
  and (_16194_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  or (_06380_, _16194_, _16192_);
  and (_16195_, _16111_, _24051_);
  and (_16196_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  or (_06390_, _16196_, _16195_);
  and (_16197_, _16111_, _23887_);
  and (_16198_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  or (_26969_, _16198_, _16197_);
  and (_16199_, _16191_, _23583_);
  and (_16200_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  or (_06396_, _16200_, _16199_);
  and (_16201_, _15988_, _24219_);
  and (_16202_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or (_06401_, _16202_, _16201_);
  and (_16203_, _15992_, _24134_);
  and (_16204_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  or (_06403_, _16204_, _16203_);
  and (_16205_, _16191_, _23887_);
  and (_16206_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  or (_06408_, _16206_, _16205_);
  and (_16207_, _16048_, _24089_);
  and (_16208_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  or (_06414_, _16208_, _16207_);
  and (_16209_, _16048_, _23996_);
  and (_16210_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_06416_, _16210_, _16209_);
  and (_16211_, _09779_, _24140_);
  and (_16212_, _16211_, _23887_);
  not (_16213_, _16211_);
  and (_16214_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  or (_06420_, _16214_, _16212_);
  and (_16215_, _15980_, _23996_);
  and (_16216_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  or (_26978_, _16216_, _16215_);
  and (_16217_, _16060_, _24219_);
  and (_16218_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or (_06428_, _16218_, _16217_);
  and (_16219_, _16191_, _24219_);
  and (_16220_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or (_06434_, _16220_, _16219_);
  and (_16221_, _16060_, _24051_);
  and (_16222_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  or (_06436_, _16222_, _16221_);
  and (_16223_, _16191_, _23996_);
  and (_16224_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_06439_, _16224_, _16223_);
  and (_16225_, _16191_, _24089_);
  and (_16226_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  or (_06444_, _16226_, _16225_);
  and (_16227_, _16137_, _23996_);
  and (_16228_, _16139_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  or (_06445_, _16228_, _16227_);
  and (_16229_, _15956_, _24219_);
  and (_16230_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or (_06457_, _16230_, _16229_);
  and (_16231_, _15956_, _23996_);
  and (_16232_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_06459_, _16232_, _16231_);
  and (_16233_, _15956_, _24051_);
  and (_16234_, _15958_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  or (_06462_, _16234_, _16233_);
  and (_16235_, _16191_, _24134_);
  and (_16236_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  or (_06465_, _16236_, _16235_);
  and (_16237_, _15716_, _24134_);
  and (_16238_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  or (_06467_, _16238_, _16237_);
  and (_16239_, _15716_, _23583_);
  and (_16240_, _15718_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  or (_26987_, _16240_, _16239_);
  and (_16241_, _15640_, _23548_);
  and (_16242_, _15642_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  or (_06477_, _16242_, _16241_);
  and (_16243_, _15567_, _23887_);
  and (_16244_, _15569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  or (_26991_, _16244_, _16243_);
  and (_16245_, _16191_, _24051_);
  and (_16246_, _16193_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  or (_26982_, _16246_, _16245_);
  and (_16247_, _12442_, _24219_);
  and (_16248_, _12444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  or (_06485_, _16248_, _16247_);
  or (_16249_, _15794_, _26570_);
  not (_16250_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_16251_, _15794_, _16250_);
  and (_16252_, _16251_, _24179_);
  and (_16253_, _16252_, _16249_);
  nor (_16254_, _24178_, _16250_);
  or (_16255_, _15794_, _24531_);
  and (_16256_, _16251_, _24539_);
  and (_16257_, _16256_, _16255_);
  or (_16258_, _16257_, _16254_);
  or (_16259_, _16258_, _16253_);
  and (_06501_, _16259_, _22731_);
  or (_16260_, _15794_, _00473_);
  not (_16261_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_16262_, _15794_, _16261_);
  and (_16263_, _16262_, _24179_);
  and (_16264_, _16263_, _16260_);
  nor (_16265_, _24178_, _16261_);
  and (_16266_, _15800_, _24562_);
  nand (_16267_, _16266_, _23504_);
  or (_16268_, _16266_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_16269_, _16268_, _24539_);
  and (_16270_, _16269_, _16267_);
  or (_16271_, _16270_, _16265_);
  or (_16272_, _16271_, _16264_);
  and (_06504_, _16272_, _22731_);
  or (_16273_, _15794_, _00393_);
  not (_16274_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_16275_, _15794_, _16274_);
  and (_16276_, _16275_, _24179_);
  and (_16277_, _16276_, _16273_);
  nor (_16278_, _24178_, _16274_);
  and (_16279_, _15800_, _24177_);
  nand (_16280_, _16279_, _23504_);
  or (_16281_, _16279_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_16282_, _16281_, _24539_);
  and (_16283_, _16282_, _16280_);
  or (_16284_, _16283_, _16278_);
  or (_16285_, _16284_, _16277_);
  and (_06506_, _16285_, _22731_);
  or (_16286_, _15794_, _00569_);
  not (_16287_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_16288_, _15794_, _16287_);
  and (_16289_, _16288_, _24179_);
  and (_16290_, _16289_, _16286_);
  nor (_16291_, _24178_, _16287_);
  and (_16292_, _15800_, _24533_);
  nand (_16293_, _16292_, _23504_);
  or (_16294_, _16292_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_16295_, _16294_, _24539_);
  and (_16296_, _16295_, _16293_);
  or (_16297_, _16296_, _16291_);
  or (_16298_, _16297_, _16290_);
  and (_06511_, _16298_, _22731_);
  or (_16299_, _15794_, _00747_);
  nand (_16300_, _15794_, _04315_);
  and (_16301_, _16300_, _24179_);
  and (_16302_, _16301_, _16299_);
  nor (_16303_, _24178_, _04315_);
  and (_16304_, _15800_, _24607_);
  nand (_16305_, _16304_, _23504_);
  or (_16306_, _16304_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_16307_, _16306_, _24539_);
  and (_16308_, _16307_, _16305_);
  or (_16309_, _16308_, _16303_);
  or (_16310_, _16309_, _16302_);
  and (_06514_, _16310_, _22731_);
  or (_16311_, _15794_, _00654_);
  nand (_16312_, _15794_, _04325_);
  and (_16313_, _16312_, _24179_);
  and (_16314_, _16313_, _16311_);
  nor (_16315_, _24178_, _04325_);
  and (_16316_, _15800_, _24636_);
  nand (_16317_, _16316_, _23504_);
  or (_16318_, _16316_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_16319_, _16318_, _24539_);
  and (_16320_, _16319_, _16317_);
  or (_16321_, _16320_, _16315_);
  or (_16322_, _16321_, _16314_);
  and (_06517_, _16322_, _22731_);
  and (_16323_, _11264_, _24051_);
  and (_16324_, _11266_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  or (_06519_, _16324_, _16323_);
  or (_16325_, _15794_, _00814_);
  nand (_16326_, _15794_, _04329_);
  and (_16327_, _16326_, _24179_);
  and (_16328_, _16327_, _16325_);
  nor (_16329_, _24178_, _04329_);
  and (_16330_, _15800_, _24594_);
  nand (_16331_, _16330_, _23504_);
  or (_16332_, _16330_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_16333_, _16332_, _24539_);
  and (_16334_, _16333_, _16331_);
  or (_16335_, _16334_, _16329_);
  or (_16336_, _16335_, _16328_);
  and (_06526_, _16336_, _22731_);
  and (_16337_, _11046_, _24089_);
  and (_16338_, _11049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  or (_06530_, _16338_, _16337_);
  and (_16339_, _16060_, _23887_);
  and (_16340_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  or (_26980_, _16340_, _16339_);
  and (_16341_, _16060_, _24089_);
  and (_16342_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  or (_06541_, _16342_, _16341_);
  and (_16343_, _16060_, _23583_);
  and (_16344_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  or (_06547_, _16344_, _16343_);
  and (_16345_, _11311_, _23548_);
  and (_16346_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  or (_06555_, _16346_, _16345_);
  and (_16347_, _09780_, _23887_);
  and (_16348_, _09782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  or (_06558_, _16348_, _16347_);
  and (_16349_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  and (_16350_, _04853_, _23996_);
  or (_06564_, _16350_, _16349_);
  and (_16351_, _04854_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  and (_16352_, _04853_, _24089_);
  or (_06569_, _16352_, _16351_);
  and (_16353_, _02478_, _23548_);
  and (_16354_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  or (_06574_, _16354_, _16353_);
  and (_16355_, _11311_, _23583_);
  and (_16356_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  or (_06604_, _16356_, _16355_);
  and (_16357_, _16060_, _24134_);
  and (_16358_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  or (_26981_, _16358_, _16357_);
  and (_16359_, _09670_, _24051_);
  and (_16360_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  or (_06614_, _16360_, _16359_);
  and (_16361_, _02996_, _24134_);
  and (_16362_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  or (_27211_, _16362_, _16361_);
  and (_16363_, _16060_, _23996_);
  and (_16364_, _16062_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or (_06627_, _16364_, _16363_);
  and (_16365_, _16211_, _23583_);
  and (_16366_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  or (_06667_, _16366_, _16365_);
  and (_26864_, _00143_, _22731_);
  and (_16367_, _26687_, _22731_);
  and (_26889_, _16367_, _26716_);
  and (_06681_, _26889_, _26811_);
  nor (_06701_, _00104_, rst);
  and (_16368_, _16211_, _24089_);
  and (_16369_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  or (_06707_, _16369_, _16368_);
  nor (_26865_[4], _25834_, rst);
  and (_26866_[7], _00124_, _22731_);
  and (_16370_, _16211_, _24051_);
  and (_16371_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  or (_06744_, _16371_, _16370_);
  and (_26887_, _02050_, _22731_);
  and (_26880_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _22731_);
  and (_16372_, _26880_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_26886_, _16372_, _26887_);
  and (_16373_, _16211_, _23996_);
  and (_16374_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  or (_26979_, _16374_, _16373_);
  nor (_16375_, _26605_, rst);
  and (_26868_, _16375_, _00339_);
  and (_26869_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _22731_);
  and (_16376_, _16211_, _24134_);
  and (_16377_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  or (_06760_, _16377_, _16376_);
  and (_16378_, _15561_, _24219_);
  and (_16379_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or (_06787_, _16379_, _16378_);
  and (_16380_, _02996_, _24051_);
  and (_16381_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  or (_06806_, _16381_, _16380_);
  and (_16382_, _00883_, _26605_);
  and (_16383_, _03853_, _26574_);
  and (_16384_, _26613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_16385_, _26606_, _00885_);
  or (_16386_, _16385_, _16384_);
  or (_16387_, _16386_, _16383_);
  or (_16388_, _16387_, _16382_);
  or (_16389_, _01362_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_16390_, _01364_, _23057_);
  or (_16391_, _16390_, _00892_);
  and (_16392_, _16391_, _16389_);
  nand (_16393_, _16392_, _23003_);
  or (_16394_, _16392_, _23003_);
  and (_16395_, _16394_, _16393_);
  and (_16396_, _16395_, _26662_);
  or (_16397_, _16396_, _16388_);
  nand (_16398_, _01306_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_16399_, _01306_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_16400_, _16399_, _26665_);
  nand (_16401_, _16400_, _16398_);
  nand (_16402_, _16401_, _00339_);
  or (_16403_, _16402_, _16397_);
  and (_16404_, _01377_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_16405_, _01377_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_16406_, _16405_, _16404_);
  or (_16407_, _16406_, _00339_);
  and (_16408_, _16407_, _22731_);
  and (_26870_[15], _16408_, _16403_);
  and (_16409_, _01382_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_16410_, _01751_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_16411_, _01751_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_16412_, _16411_, _16410_);
  not (_16413_, _16412_);
  nor (_16414_, _16413_, _01754_);
  and (_16415_, _16413_, _01754_);
  or (_16416_, _16415_, _16414_);
  or (_16417_, _16416_, _24471_);
  or (_16418_, _24470_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_16419_, _16418_, _01554_);
  and (_16420_, _16419_, _16417_);
  or (_26871_[15], _16420_, _16409_);
  nor (_16421_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_26872_, _16421_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_16422_, _15980_, _24089_);
  and (_16423_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  or (_26977_, _16423_, _16422_);
  and (_16424_, _15980_, _24134_);
  and (_16425_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  or (_06817_, _16425_, _16424_);
  and (_16426_, _15980_, _24051_);
  and (_16427_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  or (_06823_, _16427_, _16426_);
  and (_16428_, _25672_, _24089_);
  and (_16429_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  or (_06869_, _16429_, _16428_);
  and (_16430_, _16211_, _23548_);
  and (_16431_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  or (_06881_, _16431_, _16430_);
  and (_16432_, _16211_, _24219_);
  and (_16433_, _16213_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  or (_06886_, _16433_, _16432_);
  and (_16434_, _06356_, _24134_);
  and (_16435_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  or (_06897_, _16435_, _16434_);
  and (_16436_, _07779_, _24219_);
  and (_16437_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  or (_06923_, _16437_, _16436_);
  and (_16438_, _06356_, _24051_);
  and (_16439_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  or (_06928_, _16439_, _16438_);
  and (_16440_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_16441_, _04897_, _24219_);
  or (_06948_, _16441_, _16440_);
  and (_16442_, _04898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  and (_16443_, _04897_, _23548_);
  or (_06955_, _16443_, _16442_);
  and (_16444_, _16034_, _23887_);
  and (_16445_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  or (_26948_, _16445_, _16444_);
  and (_16446_, _15984_, _23996_);
  and (_16447_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or (_06960_, _16447_, _16446_);
  and (_16448_, _15984_, _24134_);
  and (_16449_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  or (_06964_, _16449_, _16448_);
  and (_26873_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _22731_);
  nand (_16450_, _22737_, _01621_);
  nand (_16451_, _16450_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_16452_, _16451_, _01773_);
  and (_26874_, _16452_, _22731_);
  and (_16453_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _22731_);
  and (_16454_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _22731_);
  and (_16455_, _16454_, _01773_);
  or (_26875_[7], _16455_, _16453_);
  nand (_06974_, _00166_, _22731_);
  nor (_16456_, _25694_, _25454_);
  nand (_16457_, _01797_, _01794_);
  and (_16458_, _16457_, _22737_);
  and (_16459_, _16458_, _23588_);
  nor (_16460_, _16458_, _23588_);
  nor (_16461_, _16460_, _16459_);
  nor (_16462_, _16461_, _16456_);
  and (_16463_, _23600_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_16464_, _16463_, _16456_);
  and (_16465_, _16464_, _01544_);
  or (_16466_, _16465_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_16467_, _16466_, _16462_);
  and (_26876_[2], _16467_, _22731_);
  and (_16468_, _24236_, _24141_);
  and (_16469_, _16468_, _24089_);
  not (_16470_, _16468_);
  and (_16471_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  or (_06978_, _16471_, _16469_);
  nand (_06980_, _00187_, _22731_);
  and (_16472_, _16468_, _23887_);
  and (_16473_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  or (_06983_, _16473_, _16472_);
  nor (_06988_, _26804_, rst);
  nor (_06990_, _00014_, rst);
  nand (_06992_, _00204_, _22731_);
  and (_16474_, _03313_, _24089_);
  and (_16475_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  or (_06994_, _16475_, _16474_);
  nor (_06997_, _00084_, rst);
  nor (_06999_, _00046_, rst);
  and (_16476_, _24349_, _24141_);
  and (_16477_, _16476_, _23583_);
  not (_16478_, _16476_);
  and (_16479_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  or (_07003_, _16479_, _16477_);
  and (_16480_, _23890_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  or (_16481_, _24244_, _23930_);
  or (_16482_, _16481_, _24275_);
  or (_16483_, _23842_, _23815_);
  or (_16484_, _23904_, _23897_);
  or (_16485_, _16484_, _16483_);
  or (_16486_, _16485_, _16482_);
  or (_16487_, _16486_, _23795_);
  or (_16488_, _01980_, _23913_);
  or (_16489_, _16488_, _09759_);
  or (_16490_, _16489_, _23835_);
  or (_16491_, _16490_, _11472_);
  or (_16492_, _16491_, _16487_);
  and (_16493_, _16492_, _24295_);
  or (_26851_[1], _16493_, _16480_);
  and (_16494_, _24141_, _23941_);
  and (_16495_, _16494_, _23996_);
  not (_16496_, _16494_);
  and (_16497_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  or (_26937_, _16497_, _16495_);
  and (_16498_, _15980_, _24219_);
  and (_16499_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  or (_07010_, _16499_, _16498_);
  and (_16500_, _23720_, _23635_);
  and (_16501_, _16500_, _23761_);
  and (_16502_, _23699_, _23675_);
  and (_16503_, _16502_, _23740_);
  and (_16504_, _22738_, _22731_);
  and (_16505_, _16504_, _23656_);
  and (_16506_, _16505_, _23612_);
  and (_16507_, _16506_, _16503_);
  and (_26878_, _16507_, _16501_);
  and (_16508_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _01836_);
  and (_16509_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_16510_, _16509_, _16508_);
  and (_26879_[7], _16510_, _22731_);
  and (_16511_, _16494_, _23887_);
  and (_16512_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  or (_07033_, _16512_, _16511_);
  and (_16513_, _24899_, _24141_);
  and (_16514_, _16513_, _23996_);
  not (_16515_, _16513_);
  and (_16516_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  or (_07037_, _16516_, _16514_);
  and (_16517_, _15980_, _23887_);
  and (_16518_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  or (_07039_, _16518_, _16517_);
  and (_16519_, _16513_, _23887_);
  and (_16520_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  or (_07043_, _16520_, _16519_);
  and (_16521_, _15980_, _23548_);
  and (_16522_, _15982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  or (_07049_, _16522_, _16521_);
  and (_16523_, _24141_, _24095_);
  and (_16524_, _16523_, _23548_);
  not (_16525_, _16523_);
  and (_16526_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  or (_07051_, _16526_, _16524_);
  and (_16527_, _16523_, _23583_);
  and (_16528_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  or (_07054_, _16528_, _16527_);
  and (_16529_, _24474_, _24141_);
  and (_16530_, _16529_, _23583_);
  not (_16531_, _16529_);
  and (_16532_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  or (_07059_, _16532_, _16530_);
  and (_16533_, _16529_, _23548_);
  and (_16534_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  or (_07061_, _16534_, _16533_);
  and (_16535_, _24141_, _24056_);
  and (_16536_, _16535_, _23996_);
  not (_16537_, _16535_);
  and (_16538_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  or (_26931_, _16538_, _16536_);
  and (_16539_, _16535_, _23583_);
  and (_16540_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  or (_07075_, _16540_, _16539_);
  and (_16541_, _24301_, _23941_);
  and (_16542_, _16541_, _24051_);
  not (_16543_, _16541_);
  and (_16544_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  or (_27225_, _16544_, _16542_);
  and (_16545_, _15708_, _24219_);
  and (_16546_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_07081_, _16546_, _16545_);
  and (_16547_, _06356_, _23548_);
  and (_16548_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  or (_07083_, _16548_, _16547_);
  and (_16549_, _15984_, _23887_);
  and (_16550_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  or (_07089_, _16550_, _16549_);
  and (_16551_, _24141_, _22974_);
  and (_16552_, _16551_, _23996_);
  not (_16553_, _16551_);
  and (_16554_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  or (_07092_, _16554_, _16552_);
  and (_16555_, _16551_, _24051_);
  and (_16556_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  or (_07094_, _16556_, _16555_);
  and (_16557_, _11441_, _24134_);
  and (_16558_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  or (_07100_, _16558_, _16557_);
  and (_16559_, _15561_, _23548_);
  and (_16560_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  or (_07103_, _16560_, _16559_);
  and (_16561_, _16523_, _24134_);
  and (_16562_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  or (_07107_, _16562_, _16561_);
  nand (_16563_, _01816_, _24043_);
  and (_16564_, _08221_, _08217_);
  and (_16565_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_16566_, _16565_, _16564_);
  and (_16567_, _16566_, _02193_);
  and (_16568_, _08221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_16569_, _16568_, _16567_);
  or (_16570_, _16569_, _01816_);
  and (_16571_, _16570_, _22731_);
  and (_07109_, _16571_, _16563_);
  and (_16572_, _16523_, _23887_);
  and (_16573_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  or (_26924_, _16573_, _16572_);
  and (_16574_, _16523_, _24219_);
  and (_16575_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  or (_07113_, _16575_, _16574_);
  and (_16576_, _15984_, _23548_);
  and (_16577_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  or (_07115_, _16577_, _16576_);
  and (_16578_, _06356_, _24219_);
  and (_16579_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_07117_, _16579_, _16578_);
  and (_16580_, _08523_, _24134_);
  and (_16581_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  or (_07123_, _16581_, _16580_);
  and (_16582_, _15984_, _24219_);
  and (_16583_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_07125_, _16583_, _16582_);
  and (_16584_, _16048_, _24051_);
  and (_16585_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  or (_07130_, _16585_, _16584_);
  and (_16586_, _16048_, _23548_);
  and (_16587_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  or (_07141_, _16587_, _16586_);
  and (_16588_, _15830_, _23887_);
  and (_16589_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  or (_26930_, _16589_, _16588_);
  and (_16590_, _16523_, _24051_);
  and (_16591_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  or (_07145_, _16591_, _16590_);
  and (_16592_, _15708_, _24089_);
  and (_16593_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  or (_07164_, _16593_, _16592_);
  and (_16594_, _15708_, _24134_);
  and (_16595_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  or (_26927_, _16595_, _16594_);
  not (_16596_, _01862_);
  and (_16597_, _01865_, _16596_);
  or (_16598_, _01867_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_26882_[3], _16598_, _22731_);
  and (_16599_, _26882_[3], _01870_);
  and (_26881_, _16599_, _16597_);
  and (_16600_, _16523_, _23996_);
  and (_16601_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  or (_07177_, _16601_, _16600_);
  and (_16602_, _16541_, _24089_);
  and (_16603_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  or (_07180_, _16603_, _16602_);
  and (_16604_, _15984_, _24089_);
  and (_16605_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  or (_07185_, _16605_, _16604_);
  and (_16606_, _16476_, _24051_);
  and (_16607_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  or (_07188_, _16607_, _16606_);
  and (_16608_, _16494_, _24089_);
  and (_16609_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  or (_07194_, _16609_, _16608_);
  and (_16610_, _16513_, _24089_);
  and (_16611_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  or (_07197_, _16611_, _16610_);
  and (_16612_, _16513_, _24219_);
  and (_16613_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  or (_26934_, _16613_, _16612_);
  and (_16614_, _16529_, _24051_);
  and (_16615_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  or (_07201_, _16615_, _16614_);
  and (_16616_, _15984_, _23583_);
  and (_16617_, _15986_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  or (_07204_, _16617_, _16616_);
  and (_16618_, _06356_, _23583_);
  and (_16619_, _06358_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  or (_27178_, _16619_, _16618_);
  and (_16620_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_16621_, _01218_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or (_16622_, _16621_, _16620_);
  and (_26883_[31], _16622_, _22731_);
  and (_16623_, _07779_, _23887_);
  and (_16624_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  or (_07214_, _16624_, _16623_);
  and (_16625_, _16535_, _24219_);
  and (_16626_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  or (_07216_, _16626_, _16625_);
  and (_16627_, _16551_, _24219_);
  and (_16628_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  or (_07221_, _16628_, _16627_);
  and (_16629_, _24017_, _23887_);
  and (_16630_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  or (_07226_, _16630_, _16629_);
  and (_16631_, _16551_, _23887_);
  and (_16632_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  or (_07232_, _16632_, _16631_);
  and (_16633_, _16523_, _24089_);
  and (_16634_, _16525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  or (_26925_, _16634_, _16633_);
  and (_16635_, _15830_, _24089_);
  and (_16636_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  or (_07245_, _16636_, _16635_);
  and (_16637_, _08523_, _24051_);
  and (_16638_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  or (_27082_, _16638_, _16637_);
  and (_16639_, _15988_, _23583_);
  and (_16640_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  or (_07251_, _16640_, _16639_);
  and (_16641_, _15988_, _23887_);
  and (_16642_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  or (_07266_, _16642_, _16641_);
  and (_16643_, _15988_, _23548_);
  and (_16644_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  or (_07270_, _16644_, _16643_);
  or (_16645_, _25694_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand (_16646_, _25694_, _25457_);
  and (_16647_, _16646_, _22731_);
  and (_26884_[31], _16647_, _16645_);
  and (_16648_, _16551_, _23548_);
  and (_16649_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  or (_07293_, _16649_, _16648_);
  and (_16650_, _16535_, _24089_);
  and (_16651_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  or (_07297_, _16651_, _16650_);
  and (_16652_, _15708_, _23548_);
  and (_16653_, _15710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  or (_07300_, _16653_, _16652_);
  and (_16654_, _03241_, _23996_);
  and (_16655_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  or (_07306_, _16655_, _16654_);
  and (_16656_, _16048_, _24134_);
  and (_16657_, _16050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  or (_07309_, _16657_, _16656_);
  and (_16658_, _03241_, _24134_);
  and (_16659_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  or (_27173_, _16659_, _16658_);
  and (_16660_, _16494_, _24219_);
  and (_16661_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  or (_07317_, _16661_, _16660_);
  and (_16662_, _15830_, _24051_);
  and (_16663_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  or (_07324_, _16663_, _16662_);
  and (_16664_, _15988_, _24134_);
  and (_16665_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  or (_26974_, _16665_, _16664_);
  and (_16666_, _24394_, _23548_);
  and (_16667_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  or (_07338_, _16667_, _16666_);
  and (_16668_, _15988_, _24051_);
  and (_16669_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  or (_07341_, _16669_, _16668_);
  and (_16670_, _24496_, _24159_);
  and (_16671_, _16670_, _24134_);
  not (_16672_, _16670_);
  and (_16673_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  or (_07344_, _16673_, _16671_);
  and (_16674_, _16670_, _24219_);
  and (_16675_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  or (_07346_, _16675_, _16674_);
  and (_16676_, _15988_, _24089_);
  and (_16677_, _15990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  or (_07349_, _16677_, _16676_);
  and (_16678_, _24496_, _24297_);
  and (_16679_, _16678_, _23887_);
  not (_16680_, _16678_);
  and (_16681_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  or (_07353_, _16681_, _16679_);
  and (_16682_, _03043_, _24134_);
  and (_16683_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  or (_07355_, _16683_, _16682_);
  and (_16684_, _05478_, _24219_);
  and (_16685_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  or (_27249_, _16685_, _16684_);
  and (_16686_, _02502_, _23548_);
  and (_16687_, _02504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  or (_07360_, _16687_, _16686_);
  and (_16688_, _02478_, _23887_);
  and (_16689_, _02480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  or (_27246_, _16689_, _16688_);
  and (_16690_, _06129_, _24219_);
  and (_16691_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  or (_07370_, _16691_, _16690_);
  and (_16692_, _15561_, _23887_);
  and (_16693_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  or (_27241_, _16693_, _16692_);
  and (_16694_, _15888_, _24051_);
  and (_16695_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  or (_07391_, _16695_, _16694_);
  and (_16696_, _15992_, _24051_);
  and (_16697_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  or (_07394_, _16697_, _16696_);
  and (_16698_, _24496_, _24372_);
  and (_16699_, _16698_, _23583_);
  not (_16700_, _16698_);
  and (_16701_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  or (_07397_, _16701_, _16699_);
  and (_16702_, _02767_, _23887_);
  and (_16703_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  or (_07399_, _16703_, _16702_);
  nor (_26867_[0], _26630_, rst);
  and (_16704_, _24496_, _24140_);
  and (_16705_, _16704_, _24089_);
  not (_16706_, _16704_);
  and (_16707_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  or (_07403_, _16707_, _16705_);
  and (_16708_, _02767_, _23548_);
  and (_16709_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  or (_27174_, _16709_, _16708_);
  and (_16710_, _15992_, _24089_);
  and (_16711_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  or (_07407_, _16711_, _16710_);
  or (_16712_, _08401_, _23880_);
  and (_16713_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_16714_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_16715_, _16714_, _16713_);
  or (_16716_, _16715_, _25608_);
  and (_16717_, _16716_, _25617_);
  and (_16718_, _16717_, _16712_);
  and (_16719_, _25603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_16720_, _16719_, _16718_);
  and (_07409_, _16720_, _22731_);
  and (_16721_, _15992_, _23583_);
  and (_16722_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  or (_26973_, _16722_, _16721_);
  and (_16723_, _02045_, _24134_);
  and (_16724_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  or (_07414_, _16724_, _16723_);
  and (_16725_, _16551_, _23583_);
  and (_16726_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  or (_07418_, _16726_, _16725_);
  and (_16727_, _02767_, _24219_);
  and (_16728_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_07425_, _16728_, _16727_);
  and (_16729_, _11311_, _23887_);
  and (_16730_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  or (_07427_, _16730_, _16729_);
  and (_16731_, _24899_, _24301_);
  and (_16732_, _16731_, _24134_);
  not (_16733_, _16731_);
  and (_16734_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  or (_07433_, _16734_, _16732_);
  and (_16735_, _05485_, _23996_);
  and (_16736_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_07444_, _16736_, _16735_);
  and (_16737_, _11441_, _24051_);
  and (_16738_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  or (_07449_, _16738_, _16737_);
  and (_16739_, _16551_, _24089_);
  and (_16740_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  or (_07456_, _16740_, _16739_);
  and (_16741_, _24451_, _24051_);
  and (_16742_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  or (_07462_, _16742_, _16741_);
  and (_16743_, _16551_, _24134_);
  and (_16744_, _16553_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  or (_07469_, _16744_, _16743_);
  and (_16745_, _15992_, _23996_);
  and (_16746_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  or (_07471_, _16746_, _16745_);
  and (_16747_, _25672_, _23996_);
  and (_16748_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_27206_, _16748_, _16747_);
  and (_16749_, _25672_, _23583_);
  and (_16750_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  or (_07499_, _16750_, _16749_);
  and (_16751_, _03241_, _23548_);
  and (_16752_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  or (_07501_, _16752_, _16751_);
  and (_16753_, _09670_, _24134_);
  and (_16754_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  or (_07503_, _16754_, _16753_);
  and (_16755_, _06208_, _23583_);
  and (_16756_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  or (_07506_, _16756_, _16755_);
  and (_16757_, _03241_, _24219_);
  and (_16758_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  or (_07511_, _16758_, _16757_);
  and (_16759_, _16541_, _23996_);
  and (_16760_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  or (_07513_, _16760_, _16759_);
  and (_16761_, _25637_, _23548_);
  and (_16762_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  or (_07515_, _16762_, _16761_);
  and (_16763_, _16111_, _23996_);
  and (_16764_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  or (_07528_, _16764_, _16763_);
  and (_16765_, _15830_, _24134_);
  and (_16766_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  or (_07535_, _16766_, _16765_);
  and (_16767_, _25658_, _24051_);
  and (_16768_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  or (_07540_, _16768_, _16767_);
  and (_16769_, _16111_, _24134_);
  and (_16770_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  or (_07542_, _16770_, _16769_);
  and (_16771_, _15888_, _24219_);
  and (_16772_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or (_07544_, _16772_, _16771_);
  and (_16773_, _24496_, _24146_);
  and (_16774_, _16773_, _23583_);
  not (_16775_, _16773_);
  and (_16776_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  or (_07546_, _16776_, _16774_);
  and (_16777_, _03241_, _23887_);
  and (_16778_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  or (_07550_, _16778_, _16777_);
  and (_16779_, _03241_, _24089_);
  and (_16780_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  or (_07554_, _16780_, _16779_);
  and (_16781_, _25479_, _24636_);
  and (_16782_, _16781_, _23504_);
  nor (_16783_, _16781_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_16784_, _16783_, _16782_);
  nand (_16785_, _16784_, _08541_);
  nand (_16786_, _25489_, _24082_);
  and (_16787_, _16786_, _22731_);
  and (_07558_, _16787_, _16785_);
  and (_16788_, _25479_, _24533_);
  nand (_16789_, _16788_, _23504_);
  or (_16790_, _16788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_16791_, _16790_, _08541_);
  and (_16792_, _16791_, _16789_);
  and (_16793_, _25489_, _23577_);
  or (_16794_, _16793_, _16792_);
  and (_07562_, _16794_, _22731_);
  and (_16795_, _03001_, _24089_);
  and (_16796_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  or (_07565_, _16796_, _16795_);
  and (_16797_, _03241_, _23583_);
  and (_16798_, _03243_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  or (_27172_, _16798_, _16797_);
  and (_16799_, _25479_, _24562_);
  nand (_16800_, _16799_, _23504_);
  or (_16801_, _16799_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_16802_, _16801_, _08541_);
  and (_16803_, _16802_, _16800_);
  and (_16804_, _25489_, _23880_);
  or (_16805_, _16804_, _16803_);
  and (_07577_, _16805_, _22731_);
  and (_16806_, _24451_, _23548_);
  and (_16807_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  or (_07580_, _16807_, _16806_);
  and (_16808_, _15992_, _23548_);
  and (_16809_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  or (_07586_, _16809_, _16808_);
  and (_16810_, _15581_, _23548_);
  and (_16811_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  or (_07588_, _16811_, _16810_);
  nand (_16812_, _03797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_16813_, _16812_, _25479_);
  or (_16814_, _16813_, _03798_);
  not (_16815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_16816_, _25528_, _16815_);
  or (_16817_, _16816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_16818_, _16817_, _25479_);
  and (_16819_, _16818_, _16814_);
  or (_16820_, _16819_, _25489_);
  nand (_16821_, _25489_, _24126_);
  and (_16822_, _16821_, _22731_);
  and (_07603_, _16822_, _16820_);
  and (_16823_, _15992_, _24219_);
  and (_16824_, _15994_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  or (_07607_, _16824_, _16823_);
  or (_16825_, _25550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_16826_, _25541_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_16827_, _25543_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_16828_, _25544_, _25531_);
  or (_16829_, _16828_, _25499_);
  and (_16830_, _16829_, _16827_);
  or (_16831_, _16830_, _16826_);
  and (_16832_, _16831_, _16825_);
  or (_16833_, _16832_, _25558_);
  nand (_16834_, _25558_, _24126_);
  and (_16835_, _16834_, _22731_);
  and (_07624_, _16835_, _16833_);
  and (_16836_, _24394_, _23887_);
  and (_16837_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  or (_07626_, _16837_, _16836_);
  and (_16838_, _25479_, _24577_);
  nand (_16839_, _16838_, _23504_);
  or (_16840_, _16838_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_16841_, _16840_, _08541_);
  and (_16842_, _16841_, _16839_);
  and (_16843_, _25489_, _24671_);
  or (_16844_, _16843_, _16842_);
  and (_07639_, _16844_, _22731_);
  and (_16845_, _05478_, _23548_);
  and (_16846_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  or (_27250_, _16846_, _16845_);
  and (_16847_, _03245_, _23583_);
  and (_16848_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  or (_07646_, _16848_, _16847_);
  and (_16849_, _16111_, _23548_);
  and (_16850_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  or (_07648_, _16850_, _16849_);
  and (_16851_, _03245_, _23887_);
  and (_16852_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  or (_07868_, _16852_, _16851_);
  and (_16853_, _15561_, _23583_);
  and (_16854_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  or (_07870_, _16854_, _16853_);
  and (_16855_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_16856_, _16855_, _25523_);
  and (_16857_, _25514_, _25507_);
  or (_16858_, _16857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_16859_, _16857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_16860_, _16859_, _16858_);
  or (_16861_, _16860_, _25531_);
  or (_16862_, _16861_, _16856_);
  or (_16863_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_16864_, _16863_, _25502_);
  and (_16865_, _16864_, _16862_);
  and (_16866_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_16867_, _25558_, _24671_);
  or (_16868_, _16867_, _16866_);
  or (_16869_, _16868_, _16865_);
  and (_07875_, _16869_, _22731_);
  and (_16870_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_16871_, _16870_, _25523_);
  nand (_16872_, _25518_, _25507_);
  and (_16873_, _16872_, _08420_);
  nor (_16874_, _16873_, _08458_);
  or (_16875_, _16874_, _25531_);
  or (_16876_, _16875_, _16871_);
  or (_16877_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_16878_, _16877_, _25502_);
  and (_16879_, _16878_, _16876_);
  and (_16880_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_16881_, _16880_, _16879_);
  and (_16882_, _08468_, _02700_);
  or (_16883_, _16882_, _16881_);
  and (_07877_, _16883_, _22731_);
  and (_16884_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_16885_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_16886_, _16885_, _25523_);
  and (_16887_, _25517_, _25507_);
  or (_16888_, _16887_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_16889_, _16888_, _16872_);
  or (_16890_, _16889_, _25531_);
  or (_16891_, _16890_, _16886_);
  or (_16892_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_16893_, _16892_, _25502_);
  and (_16894_, _16893_, _16891_);
  or (_16895_, _16894_, _16884_);
  and (_16896_, _08468_, _23577_);
  or (_16897_, _16896_, _16895_);
  and (_07879_, _16897_, _22731_);
  and (_16898_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_16899_, _16898_, _25523_);
  and (_16900_, _25516_, _25507_);
  nor (_16901_, _16900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_16902_, _16901_, _16887_);
  or (_16903_, _16902_, _25531_);
  or (_16904_, _16903_, _16899_);
  or (_16905_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_16906_, _16905_, _25502_);
  and (_16907_, _16906_, _16904_);
  and (_16908_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_16909_, _16908_, _16907_);
  and (_16910_, _08468_, _23880_);
  or (_16911_, _16910_, _16909_);
  and (_07881_, _16911_, _22731_);
  and (_16912_, _07038_, _24219_);
  and (_16913_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_27226_, _16913_, _16912_);
  and (_16914_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_16915_, _16914_, _25523_);
  and (_16916_, _25515_, _25507_);
  nor (_16917_, _16916_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_16918_, _16917_, _16900_);
  or (_16919_, _16918_, _25531_);
  or (_16920_, _16919_, _16915_);
  or (_16921_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_16922_, _16921_, _25502_);
  and (_16923_, _16922_, _16920_);
  and (_16924_, _25499_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_16925_, _25558_, _02728_);
  or (_16926_, _16925_, _16924_);
  or (_16927_, _16926_, _16923_);
  and (_07884_, _16927_, _22731_);
  and (_16928_, _25499_, _23880_);
  and (_16929_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_16930_, _16929_, _25523_);
  and (_16931_, _25508_, _25507_);
  or (_16932_, _16931_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_16933_, _16932_, _08442_);
  or (_16934_, _16933_, _25531_);
  or (_16935_, _16934_, _16930_);
  or (_16936_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_16937_, _16936_, _25502_);
  and (_16938_, _16937_, _16935_);
  and (_16939_, _25501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_16940_, _16939_, _16938_);
  or (_16941_, _16940_, _16928_);
  and (_07889_, _16941_, _22731_);
  and (_16942_, _25507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  not (_16943_, _16942_);
  nor (_16944_, _16943_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_16945_, _16943_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_16946_, _16945_, _25531_);
  or (_16947_, _16946_, _16944_);
  and (_16948_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_16949_, _16948_, _25523_);
  or (_16950_, _16949_, _16947_);
  or (_16951_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_16952_, _16951_, _25502_);
  and (_16953_, _16952_, _16950_);
  nor (_16954_, _25550_, _23542_);
  and (_16955_, _25558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_16956_, _16955_, _16954_);
  or (_16957_, _16956_, _16953_);
  and (_07891_, _16957_, _22731_);
  or (_16958_, _25507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_16959_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_16960_, _16959_, _25522_);
  or (_16961_, _16960_, _16943_);
  and (_16962_, _16961_, _16958_);
  or (_16963_, _16962_, _25531_);
  or (_16964_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_16965_, _16964_, _25502_);
  and (_16966_, _16965_, _16963_);
  and (_16967_, _25499_, _24671_);
  and (_16968_, _25558_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_16969_, _16968_, _16967_);
  or (_16970_, _16969_, _16966_);
  and (_07896_, _16970_, _22731_);
  and (_16971_, _02996_, _24219_);
  and (_16972_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  or (_07898_, _16972_, _16971_);
  and (_16973_, _16111_, _24089_);
  and (_16974_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  or (_07902_, _16974_, _16973_);
  and (_16975_, _03245_, _24134_);
  and (_16976_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  or (_07904_, _16976_, _16975_);
  nor (_16977_, _25550_, _24043_);
  and (_16978_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_16979_, _16978_, _25523_);
  nand (_16980_, _25511_, _25507_);
  nor (_16981_, _16980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_16982_, _16980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_16983_, _16982_, _25531_);
  or (_16984_, _16983_, _16981_);
  or (_16985_, _16984_, _16979_);
  or (_16986_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_16987_, _16986_, _25502_);
  and (_16988_, _16987_, _16985_);
  and (_16989_, _25501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_16990_, _16989_, _16988_);
  or (_16991_, _16990_, _16977_);
  and (_07905_, _16991_, _22731_);
  and (_16992_, _16111_, _23583_);
  and (_16993_, _16113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  or (_07908_, _16993_, _16992_);
  and (_16994_, _06208_, _24089_);
  and (_16995_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  or (_07910_, _16995_, _16994_);
  and (_16996_, _25637_, _23996_);
  and (_16997_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_07912_, _16997_, _16996_);
  nor (_16998_, _25550_, _24126_);
  and (_16999_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_17000_, _16999_, _25523_);
  and (_17001_, _25512_, _25507_);
  nor (_17002_, _17001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_17003_, _17002_, _25582_);
  or (_17004_, _17003_, _25531_);
  or (_17005_, _17004_, _17000_);
  or (_17006_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_17007_, _17006_, _25502_);
  and (_17008_, _17007_, _17005_);
  and (_17009_, _25501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_17010_, _17009_, _17008_);
  or (_17011_, _17010_, _16998_);
  and (_07914_, _17011_, _22731_);
  nor (_17012_, _25550_, _24082_);
  and (_17013_, _25539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_17014_, _17013_, _25523_);
  and (_17015_, _25510_, _25507_);
  or (_17016_, _17015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_17017_, _17016_, _16980_);
  or (_17018_, _17017_, _25531_);
  or (_17019_, _17018_, _17014_);
  or (_17020_, _08448_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_17021_, _17020_, _25502_);
  and (_17022_, _17021_, _17019_);
  and (_17023_, _25501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_17024_, _17023_, _17022_);
  or (_17025_, _17024_, _17012_);
  and (_07917_, _17025_, _22731_);
  and (_17026_, _15830_, _23996_);
  and (_17027_, _15832_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_07952_, _17027_, _17026_);
  and (_17028_, _16535_, _23548_);
  and (_17029_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  or (_07959_, _17029_, _17028_);
  and (_17030_, _15561_, _24089_);
  and (_17031_, _15563_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  or (_07961_, _17031_, _17030_);
  and (_17032_, _24372_, _24098_);
  and (_17033_, _17032_, _24219_);
  not (_17034_, _17032_);
  and (_17035_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  or (_07965_, _17035_, _17033_);
  and (_17036_, _24146_, _24098_);
  and (_17037_, _17036_, _23996_);
  not (_17038_, _17036_);
  and (_17039_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  or (_07968_, _17039_, _17037_);
  and (_17040_, _17036_, _23548_);
  and (_17041_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  or (_07972_, _17041_, _17040_);
  and (_17042_, _24140_, _24098_);
  and (_17043_, _17042_, _24089_);
  not (_17044_, _17042_);
  and (_17045_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  or (_07975_, _17045_, _17043_);
  and (_17046_, _24159_, _22982_);
  and (_17047_, _17046_, _24089_);
  not (_17048_, _17046_);
  and (_17049_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  or (_07981_, _17049_, _17047_);
  and (_17050_, _17046_, _23887_);
  and (_17051_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  or (_07983_, _17051_, _17050_);
  and (_17052_, _24297_, _22982_);
  and (_17053_, _17052_, _24089_);
  not (_17054_, _17052_);
  and (_17055_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  or (_07988_, _17055_, _17053_);
  and (_17056_, _17052_, _23887_);
  and (_17057_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  or (_07990_, _17057_, _17056_);
  and (_17058_, _24016_, _22982_);
  and (_17059_, _17058_, _24051_);
  not (_17060_, _17058_);
  and (_17061_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  or (_07993_, _17061_, _17059_);
  and (_17062_, _17058_, _23583_);
  and (_17063_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  or (_07995_, _17063_, _17062_);
  and (_17064_, _17058_, _24219_);
  and (_17065_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  or (_07997_, _17065_, _17064_);
  and (_17066_, _24236_, _22982_);
  and (_17067_, _17066_, _24134_);
  not (_17068_, _17066_);
  and (_17069_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  or (_08002_, _17069_, _17067_);
  and (_17070_, _17066_, _23887_);
  and (_17071_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  or (_08005_, _17071_, _17070_);
  and (_17072_, _24899_, _22982_);
  and (_17073_, _17072_, _24134_);
  not (_17074_, _17072_);
  and (_17075_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  or (_08012_, _17075_, _17073_);
  and (_17076_, _11360_, _24051_);
  and (_17077_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  or (_27079_, _17077_, _17076_);
  and (_17078_, _24474_, _22982_);
  and (_17079_, _17078_, _24134_);
  not (_17080_, _17078_);
  and (_17081_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  or (_08020_, _17081_, _17079_);
  and (_17082_, _17078_, _24089_);
  and (_17083_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  or (_27285_, _17083_, _17082_);
  and (_17084_, _17078_, _24219_);
  and (_17085_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_08023_, _17085_, _17084_);
  nand (_17086_, _25603_, _24126_);
  and (_17087_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_17088_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_17089_, _17088_, _17087_);
  or (_17090_, _17089_, _25603_);
  and (_17091_, _17090_, _22731_);
  and (_08237_, _17091_, _17086_);
  and (_17092_, _24057_, _23996_);
  and (_17093_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  or (_08238_, _17093_, _17092_);
  and (_17094_, _03245_, _24051_);
  and (_17095_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  or (_08240_, _17095_, _17094_);
  nand (_17096_, _25603_, _24043_);
  and (_17097_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_17098_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_17099_, _17098_, _17097_);
  or (_17100_, _17099_, _25603_);
  and (_17101_, _17100_, _22731_);
  and (_08242_, _17101_, _17096_);
  and (_17102_, _24349_, _22982_);
  and (_17103_, _17102_, _24089_);
  not (_17104_, _17102_);
  and (_17105_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  or (_08247_, _17105_, _17103_);
  and (_17106_, _16000_, _24089_);
  and (_17107_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  or (_08249_, _17107_, _17106_);
  and (_17108_, _16000_, _23583_);
  and (_17109_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  or (_08253_, _17109_, _17108_);
  and (_17110_, _23941_, _22982_);
  and (_17111_, _17110_, _24051_);
  not (_17112_, _17110_);
  and (_17113_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  or (_27291_, _17113_, _17111_);
  and (_17114_, _03255_, _24134_);
  and (_17115_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  or (_08256_, _17115_, _17114_);
  and (_17116_, _16535_, _23887_);
  and (_17117_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  or (_08259_, _17117_, _17116_);
  and (_17118_, _03255_, _24051_);
  and (_17119_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  or (_08261_, _17119_, _17118_);
  or (_17120_, _25617_, _23577_);
  and (_17121_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_17122_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_17123_, _17122_, _17121_);
  or (_17124_, _17123_, _25603_);
  and (_17125_, _17124_, _22731_);
  and (_08266_, _17125_, _17120_);
  or (_17126_, _25617_, _23880_);
  and (_17127_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_17128_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_17129_, _17128_, _17127_);
  or (_17130_, _17129_, _25603_);
  and (_17131_, _17130_, _22731_);
  and (_08268_, _17131_, _17126_);
  and (_17132_, _25610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_17133_, _25609_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_17134_, _17133_, _17132_);
  or (_17135_, _17134_, _25603_);
  nand (_17136_, _25603_, _23542_);
  and (_17137_, _17136_, _22731_);
  and (_08270_, _17137_, _17135_);
  and (_17138_, _03255_, _24089_);
  and (_17139_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  or (_08272_, _17139_, _17138_);
  and (_17140_, _17036_, _23583_);
  and (_17141_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  or (_08275_, _17141_, _17140_);
  and (_17142_, _16000_, _24134_);
  and (_17143_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  or (_08278_, _17143_, _17142_);
  and (_17144_, _16000_, _24051_);
  and (_17145_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  or (_08280_, _17145_, _17144_);
  and (_17146_, _16535_, _24051_);
  and (_17147_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  or (_08284_, _17147_, _17146_);
  and (_17148_, _17042_, _23548_);
  and (_17149_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  or (_27301_, _17149_, _17148_);
  nor (_17150_, _08401_, _24043_);
  and (_17151_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_17152_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_17153_, _17152_, _17151_);
  nor (_17154_, _17153_, _25608_);
  or (_17155_, _17154_, _08404_);
  or (_17156_, _17155_, _17150_);
  or (_17157_, _08413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_17158_, _17157_, _22731_);
  and (_08288_, _17158_, _17156_);
  and (_17159_, _17046_, _24134_);
  and (_17160_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  or (_08290_, _17160_, _17159_);
  and (_17161_, _02364_, _24219_);
  and (_17162_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_08369_, _17162_, _17161_);
  and (_17163_, _02364_, _23548_);
  and (_17164_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  or (_08381_, _17164_, _17163_);
  not (_17165_, _23855_);
  or (_26842_[1], _02006_, _17165_);
  and (_17166_, _24142_, _24051_);
  and (_17167_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  or (_08393_, _17167_, _17166_);
  and (_17168_, _22734_, _22735_);
  and (_17169_, _17168_, _26571_);
  and (_17170_, _01432_, _01411_);
  or (_17171_, _17170_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_17172_, _01391_, _01402_);
  and (_17173_, _01475_, _17172_);
  and (_17174_, _01432_, _01526_);
  and (_17175_, _01502_, _01420_);
  or (_17176_, _17175_, _17174_);
  or (_17177_, _17176_, _17173_);
  or (_17178_, _17177_, _17171_);
  and (_17179_, _17178_, _17169_);
  nor (_17180_, _17168_, _26571_);
  or (_17181_, _17180_, rst);
  or (_26843_[0], _17181_, _17179_);
  or (_17182_, _01985_, _24253_);
  or (_17183_, _02385_, _24275_);
  or (_17184_, _17183_, _17182_);
  and (_17185_, _17184_, _22737_);
  and (_17186_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_17187_, _17186_, _02359_);
  or (_17188_, _17187_, _17185_);
  and (_26846_[1], _17188_, _22731_);
  and (_17189_, _23890_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or (_17190_, _26576_, _00287_);
  or (_17191_, _17190_, _01979_);
  or (_17192_, _00240_, _04800_);
  or (_17193_, _26584_, _23894_);
  or (_17194_, _26742_, _23923_);
  or (_17195_, _17194_, _17193_);
  or (_17196_, _17195_, _17192_);
  or (_17197_, _17196_, _17191_);
  and (_17198_, _17197_, _23855_);
  or (_26845_, _17198_, _17189_);
  and (_17199_, _05478_, _23887_);
  and (_17200_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  or (_08400_, _17200_, _17199_);
  and (_17201_, _05478_, _23583_);
  and (_17202_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  or (_08408_, _17202_, _17201_);
  and (_17203_, _24409_, _24051_);
  and (_17204_, _24411_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  or (_08410_, _17204_, _17203_);
  and (_17205_, _09717_, _24134_);
  and (_17206_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  or (_08597_, _17206_, _17205_);
  or (_17207_, _04786_, _01978_);
  or (_17208_, _24267_, _23917_);
  or (_17209_, _17208_, _17207_);
  or (_17210_, _23815_, _23790_);
  or (_17211_, _26694_, _23919_);
  or (_17212_, _17211_, _17210_);
  nand (_17213_, _23838_, _01990_);
  nand (_17214_, _17213_, _26699_);
  or (_17215_, _17214_, _03906_);
  or (_17216_, _23836_, _23833_);
  or (_17217_, _17216_, _17215_);
  or (_17218_, _17217_, _17212_);
  or (_17219_, _26754_, _26731_);
  and (_17220_, _23927_, _23687_);
  or (_17221_, _17220_, _01979_);
  or (_17222_, _17221_, _17219_);
  or (_17223_, _17222_, _09756_);
  or (_17224_, _17223_, _17218_);
  or (_17225_, _17224_, _17209_);
  and (_17226_, _17225_, _22737_);
  and (_17227_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_17228_, _17227_, _02010_);
  or (_17229_, _17228_, _17226_);
  and (_26846_[0], _17229_, _22731_);
  and (_17230_, _09717_, _23996_);
  and (_17231_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_08602_, _17231_, _17230_);
  or (_17232_, _23703_, _26679_);
  or (_17233_, _22736_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_17234_, _17233_, _22731_);
  and (_26844_[4], _17234_, _17232_);
  and (_17235_, _09717_, _24051_);
  and (_17236_, _09719_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  or (_27072_, _17236_, _17235_);
  and (_26841_[0], _26713_, _22731_);
  or (_17237_, _23765_, _26679_);
  or (_17238_, _22736_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_17239_, _17238_, _22731_);
  and (_26844_[5], _17239_, _17237_);
  and (_17240_, _24350_, _23548_);
  and (_17241_, _24352_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  or (_27057_, _17241_, _17240_);
  or (_17242_, _23660_, _26679_);
  or (_17243_, _22736_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_17244_, _17243_, _22731_);
  and (_26844_[1], _17244_, _17242_);
  and (_17245_, _02364_, _24051_);
  and (_17246_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  or (_08629_, _17246_, _17245_);
  or (_17247_, _23639_, _26679_);
  or (_17248_, _22736_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_17249_, _17248_, _22731_);
  and (_26844_[2], _17249_, _17247_);
  and (_17250_, _02364_, _24134_);
  and (_17251_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  or (_08634_, _17251_, _17250_);
  and (_17252_, _05460_, _24134_);
  and (_17253_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  or (_08650_, _17253_, _17252_);
  and (_17254_, _05460_, _23996_);
  and (_17255_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or (_08655_, _17255_, _17254_);
  and (_17256_, _03001_, _24051_);
  and (_17257_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  or (_27216_, _17257_, _17256_);
  nand (_17258_, _16094_, _24082_);
  nor (_17259_, _16100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_17260_, _17259_, _16101_);
  or (_17261_, _17260_, _02616_);
  and (_17262_, _17261_, _02295_);
  and (_17263_, _17262_, _17258_);
  and (_17264_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_08662_, _17264_, _17263_);
  and (_17265_, _24442_, _24219_);
  and (_17266_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  or (_08667_, _17266_, _17265_);
  and (_17267_, _17052_, _24134_);
  and (_17268_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  or (_08694_, _17268_, _17267_);
  and (_17269_, _17058_, _23996_);
  and (_17270_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  or (_27297_, _17270_, _17269_);
  nor (_17271_, _08401_, _24082_);
  and (_17272_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_17273_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor (_17274_, _17273_, _17272_);
  nor (_17275_, _17274_, _25608_);
  or (_17276_, _17275_, _08404_);
  or (_17277_, _17276_, _17271_);
  or (_17278_, _08413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_17279_, _17278_, _22731_);
  and (_08701_, _17279_, _17277_);
  or (_17280_, _08401_, _23577_);
  and (_17281_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_17282_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_17283_, _17282_, _17281_);
  or (_17284_, _17283_, _25608_);
  and (_17285_, _17284_, _25617_);
  and (_17286_, _17285_, _17280_);
  and (_17287_, _25603_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_17288_, _17287_, _17286_);
  and (_08711_, _17288_, _22731_);
  and (_17289_, _24142_, _23887_);
  and (_17290_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  or (_08728_, _17290_, _17289_);
  or (_17291_, _23681_, _26679_);
  or (_17292_, _22736_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_17293_, _17292_, _22731_);
  and (_26844_[0], _17293_, _17291_);
  and (_17294_, _05460_, _24089_);
  and (_17295_, _05462_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  or (_08738_, _17295_, _17294_);
  nand (_17296_, _23615_, _22736_);
  or (_17297_, _22736_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_17298_, _17297_, _22731_);
  and (_26844_[3], _17298_, _17296_);
  or (_17299_, _23745_, _26679_);
  or (_17300_, _22736_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_17301_, _17300_, _22731_);
  and (_26844_[6], _17301_, _17299_);
  and (_17302_, _03355_, _24219_);
  and (_17303_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_08780_, _17303_, _17302_);
  and (_17304_, _11360_, _24089_);
  and (_17305_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  or (_08782_, _17305_, _17304_);
  and (_17306_, _17110_, _23548_);
  and (_17307_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  or (_08799_, _17307_, _17306_);
  and (_17308_, _17072_, _23583_);
  and (_17309_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  or (_08802_, _17309_, _17308_);
  and (_17310_, _17102_, _24134_);
  and (_17311_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  or (_08809_, _17311_, _17310_);
  and (_17312_, _17032_, _23548_);
  and (_17313_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  or (_08812_, _17313_, _17312_);
  and (_17314_, _17042_, _24051_);
  and (_17315_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  or (_08814_, _17315_, _17314_);
  and (_17316_, _24237_, _23548_);
  and (_17317_, _24239_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  or (_08817_, _17317_, _17316_);
  and (_17318_, _03245_, _24219_);
  and (_17319_, _03247_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  or (_27169_, _17319_, _17318_);
  and (_17320_, _16731_, _23996_);
  and (_17321_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  or (_08825_, _17321_, _17320_);
  nor (_26867_[7], _00139_, rst);
  and (_17322_, _17072_, _24219_);
  and (_17323_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  or (_08847_, _17323_, _17322_);
  and (_17324_, _17102_, _24219_);
  and (_17325_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_08851_, _17325_, _17324_);
  and (_17326_, _17052_, _23996_);
  and (_17327_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  or (_08855_, _17327_, _17326_);
  and (_17328_, _16185_, _23996_);
  and (_17329_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or (_08862_, _17329_, _17328_);
  and (_17330_, _08523_, _24219_);
  and (_17331_, _08525_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  or (_08865_, _17331_, _17330_);
  and (_17332_, _11360_, _23996_);
  and (_17333_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or (_08873_, _17333_, _17332_);
  and (_17334_, _24297_, _24098_);
  and (_17335_, _17334_, _24089_);
  not (_17336_, _17334_);
  and (_17337_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  or (_08887_, _17337_, _17335_);
  and (_17338_, _24098_, _24016_);
  and (_17339_, _17338_, _24134_);
  not (_17340_, _17338_);
  and (_17341_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  or (_08892_, _17341_, _17339_);
  and (_17342_, _17338_, _23548_);
  and (_17343_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  or (_08896_, _17343_, _17342_);
  and (_17344_, _24236_, _24098_);
  and (_17345_, _17344_, _23996_);
  not (_17346_, _17344_);
  and (_17347_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  or (_26910_, _17347_, _17345_);
  and (_17348_, _03255_, _23996_);
  and (_17349_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_08903_, _17349_, _17348_);
  and (_17350_, _16185_, _24134_);
  and (_17351_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  or (_08905_, _17351_, _17350_);
  nand (_17352_, _25608_, _24210_);
  or (_17353_, _25605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_17354_, _25606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_17355_, _17354_, _17353_);
  or (_17356_, _17355_, _25608_);
  and (_17357_, _17356_, _17352_);
  or (_17358_, _17357_, _08404_);
  or (_17359_, _08413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_17360_, _17359_, _22731_);
  and (_08907_, _17360_, _17358_);
  and (_17361_, _16535_, _24134_);
  and (_17362_, _16537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  or (_08912_, _17362_, _17361_);
  and (_17363_, _24349_, _24098_);
  and (_17364_, _17363_, _24134_);
  not (_17365_, _17363_);
  and (_17366_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  or (_08923_, _17366_, _17364_);
  and (_17367_, _17363_, _23583_);
  and (_17368_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  or (_08925_, _17368_, _17367_);
  and (_17369_, _24098_, _23941_);
  and (_17370_, _17369_, _24089_);
  not (_17371_, _17369_);
  and (_17372_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  or (_08932_, _17372_, _17370_);
  and (_17373_, _15581_, _23887_);
  and (_17374_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  or (_08947_, _17374_, _17373_);
  and (_17375_, _05478_, _24089_);
  and (_17376_, _05480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  or (_08949_, _17376_, _17375_);
  and (_17377_, _24518_, _24134_);
  and (_17378_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  or (_27220_, _17378_, _17377_);
  and (_26840_[7], _23724_, _22731_);
  and (_17379_, _24899_, _24098_);
  and (_17380_, _17379_, _24051_);
  not (_17381_, _17379_);
  and (_17382_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  or (_26903_, _17382_, _17380_);
  and (_17383_, _17379_, _24219_);
  and (_17384_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_08986_, _17384_, _17383_);
  and (_17385_, _24474_, _24098_);
  and (_17386_, _17385_, _24134_);
  not (_17387_, _17385_);
  and (_17388_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  or (_08989_, _17388_, _17386_);
  and (_17389_, _17385_, _23548_);
  and (_17390_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  or (_08992_, _17390_, _17389_);
  and (_17391_, _24223_, _24098_);
  and (_17392_, _17391_, _24089_);
  not (_17393_, _17391_);
  and (_17394_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  or (_08995_, _17394_, _17392_);
  and (_17395_, _24319_, _24098_);
  and (_17396_, _17395_, _23996_);
  not (_17397_, _17395_);
  and (_17398_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  or (_08999_, _17398_, _17396_);
  and (_17399_, _16000_, _23548_);
  and (_17400_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  or (_09002_, _17400_, _17399_);
  and (_17401_, _03269_, _23996_);
  and (_17402_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  or (_09004_, _17402_, _17401_);
  and (_17403_, _17395_, _24089_);
  and (_17404_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  or (_09009_, _17404_, _17403_);
  and (_17405_, _16541_, _23887_);
  and (_17406_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  or (_09014_, _17406_, _17405_);
  and (_17407_, _16541_, _23548_);
  and (_17408_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  or (_09017_, _17408_, _17407_);
  and (_17409_, _17395_, _23548_);
  and (_17410_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  or (_09034_, _17410_, _17409_);
  and (_17411_, _24098_, _22974_);
  and (_17412_, _17411_, _24134_);
  not (_17413_, _17411_);
  and (_17414_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  or (_09038_, _17414_, _17412_);
  and (_17415_, _17411_, _23583_);
  and (_17416_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  or (_09042_, _17416_, _17415_);
  and (_17417_, _24098_, _24056_);
  and (_17418_, _17417_, _24051_);
  not (_17419_, _17417_);
  and (_17420_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  or (_26900_, _17420_, _17418_);
  and (_17421_, _17417_, _23583_);
  and (_17422_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  or (_09048_, _17422_, _17421_);
  and (_17423_, _16000_, _24219_);
  and (_17424_, _16002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_09056_, _17424_, _17423_);
  and (_17425_, _17334_, _23548_);
  and (_17426_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  or (_09057_, _17426_, _17425_);
  and (_17427_, _03269_, _24134_);
  and (_17428_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  or (_09059_, _17428_, _17427_);
  and (_17429_, _03269_, _24051_);
  and (_17430_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  or (_09061_, _17430_, _17429_);
  and (_17431_, _16121_, _23583_);
  and (_17432_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  or (_09063_, _17432_, _17431_);
  and (_17433_, _16185_, _23548_);
  and (_17434_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  or (_09069_, _17434_, _17433_);
  and (_17435_, _17338_, _23583_);
  and (_17436_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  or (_26913_, _17436_, _17435_);
  nand (_17437_, _16094_, _23989_);
  or (_17438_, _02267_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_17439_, _02268_, _15660_);
  and (_17440_, _17439_, _17438_);
  and (_17441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_17442_, _02277_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  not (_17443_, _02271_);
  nor (_17444_, _02278_, _17443_);
  and (_17445_, _17444_, _17442_);
  or (_17446_, _17445_, _17441_);
  or (_17447_, _17446_, _17440_);
  or (_17448_, _17447_, _02616_);
  and (_17449_, _17448_, _02295_);
  and (_17450_, _17449_, _17437_);
  and (_17451_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_09079_, _17451_, _17450_);
  and (_17452_, _11360_, _24219_);
  and (_17453_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or (_09096_, _17453_, _17452_);
  and (_17454_, _08435_, _23887_);
  and (_17455_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  or (_09103_, _17455_, _17454_);
  and (_17456_, _17344_, _23887_);
  and (_17457_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  or (_26907_, _17457_, _17456_);
  and (_17458_, _17363_, _24219_);
  and (_17459_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  or (_09108_, _17459_, _17458_);
  and (_17460_, _17369_, _23548_);
  and (_17461_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  or (_26904_, _17461_, _17460_);
  and (_17462_, _17379_, _23887_);
  and (_17463_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  or (_09112_, _17463_, _17462_);
  and (_17464_, _17385_, _23583_);
  and (_17465_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  or (_09113_, _17465_, _17464_);
  and (_17466_, _16529_, _24219_);
  and (_17467_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_09119_, _17467_, _17466_);
  and (_17468_, _16185_, _24219_);
  and (_17469_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or (_09122_, _17469_, _17468_);
  and (_17470_, _17417_, _23996_);
  and (_17471_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_09130_, _17471_, _17470_);
  and (_17472_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_17473_, _17472_, _26165_);
  and (_17474_, _17472_, _26165_);
  or (_17475_, _17474_, _17473_);
  and (_09133_, _17475_, _22731_);
  or (_17476_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_17477_, _17476_, _22731_);
  nand (_17478_, _24189_, _24043_);
  and (_09136_, _17478_, _17477_);
  and (_17479_, _17334_, _24051_);
  and (_17480_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  or (_09139_, _17480_, _17479_);
  and (_09141_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _22731_);
  and (_09145_, _00855_, _22731_);
  and (_09148_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _22731_);
  or (_17481_, _23528_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_17482_, _17472_, rst);
  and (_09152_, _17482_, _17481_);
  and (_17483_, _16529_, _23887_);
  and (_17484_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  or (_09157_, _17484_, _17483_);
  and (_17485_, _03255_, _23887_);
  and (_17486_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  or (_09159_, _17486_, _17485_);
  and (_17487_, _17363_, _24089_);
  and (_17488_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  or (_09177_, _17488_, _17487_);
  and (_17489_, _17369_, _24051_);
  and (_17490_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  or (_09180_, _17490_, _17489_);
  and (_17491_, _17385_, _23996_);
  and (_17492_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  or (_09183_, _17492_, _17491_);
  and (_17493_, _17395_, _23887_);
  and (_17494_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  or (_09188_, _17494_, _17493_);
  and (_17495_, _17417_, _24219_);
  and (_17496_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_09191_, _17496_, _17495_);
  and (_17497_, _16529_, _24089_);
  and (_17498_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  or (_09196_, _17498_, _17497_);
  and (_17499_, _17379_, _24134_);
  and (_17500_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  or (_09198_, _17500_, _17499_);
  and (_17501_, _16529_, _24134_);
  and (_17502_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  or (_09201_, _17502_, _17501_);
  and (_17503_, _25637_, _24134_);
  and (_17504_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  or (_09207_, _17504_, _17503_);
  and (_17505_, _17391_, _23996_);
  and (_17506_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  or (_09209_, _17506_, _17505_);
  and (_17507_, _17110_, _23996_);
  and (_17508_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  or (_09211_, _17508_, _17507_);
  and (_17509_, _25637_, _24089_);
  and (_17510_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  or (_09214_, _17510_, _17509_);
  and (_17511_, _17391_, _24051_);
  and (_17512_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  or (_09216_, _17512_, _17511_);
  and (_17513_, _16121_, _24134_);
  and (_17514_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  or (_09218_, _17514_, _17513_);
  and (_17515_, _03255_, _23548_);
  and (_17516_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  or (_09220_, _17516_, _17515_);
  and (_17517_, _03255_, _24219_);
  and (_17518_, _03257_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or (_09224_, _17518_, _17517_);
  and (_17519_, _17110_, _24089_);
  and (_17520_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  or (_09226_, _17520_, _17519_);
  and (_17521_, _16185_, _24089_);
  and (_17522_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  or (_09228_, _17522_, _17521_);
  and (_17523_, _25672_, _24134_);
  and (_17524_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  or (_09230_, _17524_, _17523_);
  and (_17525_, _16185_, _23583_);
  and (_17526_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  or (_09232_, _17526_, _17525_);
  and (_17527_, _16731_, _23887_);
  and (_17528_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  or (_09256_, _17528_, _17527_);
  and (_17529_, _16731_, _23548_);
  and (_17530_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  or (_09268_, _17530_, _17529_);
  and (_17531_, _08559_, _23996_);
  and (_17532_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  or (_09270_, _17532_, _17531_);
  and (_17533_, _16731_, _24051_);
  and (_17534_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  or (_09276_, _17534_, _17533_);
  and (_17535_, _16731_, _24089_);
  and (_17536_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  or (_27223_, _17536_, _17535_);
  and (_17537_, _24155_, _23996_);
  and (_17538_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  or (_09287_, _17538_, _17537_);
  and (_17539_, _11360_, _23887_);
  and (_17540_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  or (_27078_, _17540_, _17539_);
  and (_17541_, _11360_, _23548_);
  and (_17542_, _11362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  or (_09317_, _17542_, _17541_);
  and (_17543_, _04812_, _24219_);
  and (_17544_, _04815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_09328_, _17544_, _17543_);
  and (_17545_, _24496_, _24016_);
  and (_17546_, _17545_, _23548_);
  not (_17547_, _17545_);
  and (_17548_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  or (_09331_, _17548_, _17546_);
  and (_17549_, _02514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  and (_17550_, _02513_, _24051_);
  or (_09347_, _17550_, _17549_);
  and (_17551_, _06208_, _24134_);
  and (_17552_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  or (_09357_, _17552_, _17551_);
  and (_17553_, _06208_, _24051_);
  and (_17554_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  or (_09367_, _17554_, _17553_);
  and (_17555_, _08559_, _23887_);
  and (_17556_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  or (_09391_, _17556_, _17555_);
  and (_17557_, _08559_, _23548_);
  and (_17558_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  or (_09402_, _17558_, _17557_);
  and (_17559_, _02996_, _23996_);
  and (_17560_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  or (_09412_, _17560_, _17559_);
  and (_17561_, _08559_, _24219_);
  and (_17562_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  or (_09416_, _17562_, _17561_);
  and (_17563_, _17545_, _23887_);
  and (_17564_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  or (_09427_, _17564_, _17563_);
  not (_17565_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_17566_, _02205_, _17565_);
  or (_17567_, _02321_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_17568_, _17567_, _08225_);
  nor (_17569_, _17568_, _02219_);
  nor (_17570_, _17569_, _02323_);
  nor (_17571_, _17570_, _17566_);
  nor (_17572_, _17571_, _01816_);
  and (_09462_, _17572_, _01815_);
  and (_17573_, _06208_, _23996_);
  and (_17574_, _06210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_27221_, _17574_, _17573_);
  and (_17575_, _12429_, _24134_);
  and (_17576_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  or (_09513_, _17576_, _17575_);
  and (_17577_, _08559_, _24051_);
  and (_17578_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  or (_09544_, _17578_, _17577_);
  nor (_26867_[6], _00069_, rst);
  and (_17579_, _11311_, _24134_);
  and (_17580_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  or (_09613_, _17580_, _17579_);
  and (_17581_, _24301_, _22974_);
  and (_17582_, _17581_, _23996_);
  not (_17583_, _17581_);
  and (_17584_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  or (_09630_, _17584_, _17582_);
  and (_17585_, _03043_, _23887_);
  and (_17586_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  or (_09649_, _17586_, _17585_);
  and (_17587_, _03043_, _23548_);
  and (_17588_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  or (_09662_, _17588_, _17587_);
  and (_17589_, _17581_, _24134_);
  and (_17590_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  or (_09664_, _17590_, _17589_);
  and (_17591_, _03043_, _24219_);
  and (_17592_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  or (_09666_, _17592_, _17591_);
  and (_17593_, _08435_, _23548_);
  and (_17594_, _08437_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  or (_09686_, _17594_, _17593_);
  and (_17595_, _15888_, _23887_);
  and (_17596_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  or (_09688_, _17596_, _17595_);
  and (_17597_, _15888_, _23548_);
  and (_17598_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  or (_09691_, _17598_, _17597_);
  and (_17599_, _15888_, _24089_);
  and (_17600_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  or (_09721_, _17600_, _17599_);
  and (_17601_, _16121_, _24089_);
  and (_17602_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  or (_09735_, _17602_, _17601_);
  and (_17603_, _24179_, _22867_);
  and (_17604_, _17603_, _24174_);
  nand (_17605_, _17604_, _24533_);
  and (_17606_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_17607_, _15912_, _24178_);
  and (_17608_, _17607_, _22869_);
  and (_17609_, _17608_, _00747_);
  or (_17610_, _17609_, _17606_);
  or (_17611_, _17610_, _04433_);
  nand (_17612_, _04433_, _01281_);
  and (_17613_, _17612_, _22731_);
  and (_09741_, _17613_, _17611_);
  and (_17614_, _08559_, _24089_);
  and (_17615_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  or (_09743_, _17615_, _17614_);
  and (_17616_, _17391_, _24134_);
  and (_17617_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  or (_26898_, _17617_, _17616_);
  and (_17619_, _17110_, _24134_);
  and (_17620_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  or (_09748_, _17620_, _17619_);
  and (_17621_, _16529_, _23996_);
  and (_17622_, _16531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_09755_, _17622_, _17621_);
  and (_17623_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_17624_, _17608_, _00883_);
  or (_17625_, _17624_, _17623_);
  or (_17626_, _17625_, _04433_);
  not (_17627_, _04433_);
  or (_17628_, _17627_, _03853_);
  and (_17629_, _17628_, _22731_);
  and (_09766_, _17629_, _17626_);
  and (_17630_, _17417_, _23548_);
  and (_17631_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  or (_09768_, _17631_, _17630_);
  and (_17632_, _17102_, _23548_);
  and (_17633_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  or (_09770_, _17633_, _17632_);
  and (_17634_, _17604_, _24562_);
  nor (_17635_, _17634_, _04433_);
  or (_17636_, _17635_, _26570_);
  not (_17637_, _17635_);
  or (_17638_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_17639_, _17638_, _22731_);
  and (_09776_, _17639_, _17636_);
  not (_17640_, _01520_);
  or (_17641_, _17176_, _17640_);
  or (_17642_, _17641_, _17171_);
  and (_17643_, _01434_, _01384_);
  and (_17644_, _01475_, _01424_);
  or (_17645_, _01431_, _01387_);
  and (_17646_, _17645_, _01488_);
  or (_17647_, _17646_, _17644_);
  or (_17648_, _17647_, _17643_);
  or (_17649_, _01528_, _01492_);
  or (_17650_, _17173_, _01522_);
  or (_17651_, _17650_, _17649_);
  not (_17652_, _01448_);
  nor (_17653_, _01539_, _17652_);
  nand (_17654_, _17653_, _01414_);
  or (_17655_, _17654_, _17651_);
  or (_17656_, _17655_, _17648_);
  or (_17657_, _17656_, _17642_);
  and (_17658_, _17657_, _22738_);
  nor (_17659_, _17169_, _02002_);
  or (_17660_, _17659_, rst);
  or (_26843_[1], _17660_, _17658_);
  and (_17661_, _16185_, _23887_);
  and (_17662_, _16187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  or (_09788_, _17662_, _17661_);
  or (_17663_, _17635_, _00569_);
  or (_17664_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_17665_, _17664_, _22731_);
  and (_09800_, _17665_, _17663_);
  and (_17666_, _17102_, _23887_);
  and (_17667_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  or (_27292_, _17667_, _17666_);
  or (_17668_, _24246_, _17165_);
  or (_26842_[2], _17668_, _02008_);
  and (_17669_, _24518_, _24051_);
  and (_17670_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  or (_09807_, _17670_, _17669_);
  and (_17671_, _17417_, _23887_);
  and (_17672_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  or (_09810_, _17672_, _17671_);
  and (_17673_, _03269_, _23548_);
  and (_17674_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  or (_27166_, _17674_, _17673_);
  not (_17675_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_17676_, _25481_, _17675_);
  or (_17677_, _17676_, _25482_);
  and (_17678_, _17677_, _00308_);
  and (_17679_, _00312_, _23504_);
  and (_17680_, _00311_, _17675_);
  or (_17681_, _17680_, _00308_);
  or (_17682_, _17681_, _17679_);
  nand (_17683_, _17682_, _25684_);
  or (_17684_, _17683_, _17678_);
  nand (_17685_, _25683_, _23989_);
  and (_17686_, _17685_, _22731_);
  and (_09826_, _17686_, _17684_);
  and (_17687_, _17417_, _24089_);
  and (_17688_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  or (_26899_, _17688_, _17687_);
  nand (_17689_, _17637_, _00813_);
  or (_17690_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_17691_, _17690_, _22731_);
  and (_09835_, _17691_, _17689_);
  or (_17692_, _17635_, _00473_);
  or (_17693_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_17694_, _17693_, _22731_);
  and (_09837_, _17694_, _17692_);
  and (_17695_, _17102_, _23583_);
  and (_17696_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  or (_09844_, _17696_, _17695_);
  and (_17697_, _24518_, _23996_);
  and (_17698_, _24520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  or (_09846_, _17698_, _17697_);
  and (_17699_, _17417_, _24134_);
  and (_17700_, _17419_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  or (_09854_, _17700_, _17699_);
  and (_17701_, _17102_, _24051_);
  and (_17702_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  or (_27293_, _17702_, _17701_);
  and (_17703_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_17704_, _17608_, _00654_);
  or (_17705_, _17704_, _17703_);
  or (_17706_, _17705_, _04433_);
  nand (_17707_, _04433_, _01192_);
  and (_17708_, _17707_, _22731_);
  and (_09864_, _17708_, _17706_);
  and (_17709_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_17710_, _17608_, _00569_);
  or (_17711_, _17710_, _17709_);
  or (_17712_, _17711_, _04433_);
  nand (_17713_, _04433_, _01121_);
  and (_17714_, _17713_, _22731_);
  and (_09875_, _17714_, _17712_);
  and (_17715_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_17716_, _17608_, _00473_);
  or (_17717_, _17716_, _17715_);
  or (_17718_, _17717_, _04433_);
  nand (_17719_, _04433_, _01061_);
  and (_17720_, _17719_, _22731_);
  and (_09881_, _17720_, _17718_);
  and (_17721_, _24099_, _23996_);
  and (_17722_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_09884_, _17722_, _17721_);
  and (_17723_, _24057_, _24051_);
  and (_17724_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  or (_09886_, _17724_, _17723_);
  and (_17725_, _09670_, _23887_);
  and (_17726_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  or (_09891_, _17726_, _17725_);
  and (_17727_, _03269_, _23887_);
  and (_17728_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  or (_27167_, _17728_, _17727_);
  and (_17729_, _09670_, _24219_);
  and (_17730_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  or (_09896_, _17730_, _17729_);
  and (_17731_, _17411_, _24219_);
  and (_17732_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_26895_, _17732_, _17731_);
  and (_17733_, _24134_, _24057_);
  and (_17734_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  or (_09908_, _17734_, _17733_);
  or (_17735_, _17635_, _00393_);
  or (_17736_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_17737_, _17736_, _22731_);
  and (_09911_, _17737_, _17735_);
  or (_17738_, _17635_, _00747_);
  or (_17739_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_17740_, _17739_, _22731_);
  and (_09914_, _17740_, _17738_);
  or (_17741_, _17635_, _00654_);
  or (_17742_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_17743_, _17742_, _22731_);
  and (_09916_, _17743_, _17741_);
  and (_17744_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_17745_, _17608_, _00393_);
  or (_17746_, _17745_, _17744_);
  or (_17747_, _17746_, _04433_);
  nand (_17748_, _04433_, _01009_);
  and (_17749_, _17748_, _22731_);
  and (_09918_, _17749_, _17747_);
  and (_17750_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_17751_, _17608_, _26570_);
  or (_17753_, _17751_, _17750_);
  or (_17754_, _17753_, _04433_);
  or (_17755_, _17627_, _00939_);
  and (_17756_, _17755_, _22731_);
  and (_09920_, _17756_, _17754_);
  and (_17757_, _09670_, _24089_);
  and (_17758_, _09672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  or (_27204_, _17758_, _17757_);
  and (_17759_, _16004_, _23583_);
  and (_17760_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  or (_26967_, _17760_, _17759_);
  or (_17761_, _17635_, _00883_);
  or (_17762_, _17637_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_17763_, _17762_, _22731_);
  and (_09929_, _17763_, _17761_);
  and (_17764_, _17411_, _23548_);
  and (_17765_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  or (_09939_, _17765_, _17764_);
  and (_17766_, _16004_, _23887_);
  and (_17767_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  or (_26966_, _17767_, _17766_);
  and (_17769_, _25672_, _24219_);
  and (_17770_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_27205_, _17770_, _17769_);
  and (_17771_, _17078_, _23548_);
  and (_17772_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  or (_09950_, _17772_, _17771_);
  and (_17773_, _17411_, _23887_);
  and (_17774_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  or (_09953_, _17774_, _17773_);
  nand (_17775_, _16094_, _25951_);
  nor (_17776_, _16099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_17777_, _17776_, _16100_);
  or (_17778_, _17777_, _02616_);
  and (_17779_, _17778_, _02295_);
  and (_17780_, _17779_, _17775_);
  and (_17781_, _02440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_09955_, _17781_, _17780_);
  nor (_17782_, _17605_, _00813_);
  and (_17783_, _17605_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_17784_, _17783_, _04433_);
  or (_17785_, _17784_, _17782_);
  nand (_17786_, _04433_, _01353_);
  and (_17787_, _17786_, _22731_);
  and (_09959_, _17787_, _17785_);
  and (_17788_, _17411_, _24089_);
  and (_17789_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  or (_09961_, _17789_, _17788_);
  and (_17790_, _17078_, _23887_);
  and (_17791_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  or (_09966_, _17791_, _17790_);
  and (_17792_, _02364_, _23887_);
  and (_17793_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  or (_27207_, _17793_, _17792_);
  and (_17794_, _15581_, _24219_);
  and (_17795_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  or (_09970_, _17795_, _17794_);
  and (_17796_, _17411_, _24051_);
  and (_17797_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  or (_09972_, _17797_, _17796_);
  and (_17798_, _17078_, _23583_);
  and (_17799_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  or (_09974_, _17799_, _17798_);
  and (_17800_, _17581_, _24051_);
  and (_17801_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  or (_09977_, _17801_, _17800_);
  and (_17802_, _02364_, _23996_);
  and (_17803_, _02366_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_09980_, _17803_, _17802_);
  and (_17804_, _16121_, _24051_);
  and (_17805_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  or (_09996_, _17805_, _17804_);
  and (_17806_, _15581_, _24089_);
  and (_17807_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  or (_10001_, _17807_, _17806_);
  and (_17808_, _16004_, _24089_);
  and (_17809_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  or (_10003_, _17809_, _17808_);
  and (_17810_, _17411_, _23996_);
  and (_17811_, _17413_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_10006_, _17811_, _17810_);
  and (_17812_, _17078_, _24051_);
  and (_17813_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  or (_10008_, _17813_, _17812_);
  and (_17814_, _15581_, _23583_);
  and (_17815_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  or (_27209_, _17815_, _17814_);
  and (_17816_, _17078_, _23996_);
  and (_17817_, _17080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_27286_, _17817_, _17816_);
  and (_17819_, _17395_, _24219_);
  and (_17820_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  or (_10018_, _17820_, _17819_);
  and (_17821_, _16004_, _24134_);
  and (_17822_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  or (_26968_, _17822_, _17821_);
  and (_17823_, _17072_, _23548_);
  and (_17824_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  or (_10040_, _17824_, _17823_);
  and (_17825_, _02996_, _24089_);
  and (_17826_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  or (_10043_, _17826_, _17825_);
  and (_17827_, _17395_, _23583_);
  and (_17828_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  or (_10045_, _17828_, _17827_);
  and (_17829_, _08559_, _23583_);
  and (_17830_, _08561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  or (_10048_, _17830_, _17829_);
  and (_17831_, _16004_, _24051_);
  and (_17832_, _16006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  or (_10050_, _17832_, _17831_);
  and (_17833_, _17395_, _24051_);
  and (_17834_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  or (_10055_, _17834_, _17833_);
  and (_17835_, _24451_, _24219_);
  and (_17836_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_10059_, _17836_, _17835_);
  and (_17837_, _17072_, _23887_);
  and (_17838_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  or (_10061_, _17838_, _17837_);
  and (_17839_, _17072_, _24089_);
  and (_17840_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  or (_10070_, _17840_, _17839_);
  and (_17841_, _17395_, _24134_);
  and (_17842_, _17397_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  or (_26896_, _17842_, _17841_);
  and (_17843_, _24451_, _23583_);
  and (_17844_, _24453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  or (_27212_, _17844_, _17843_);
  and (_17845_, _03001_, _23583_);
  and (_17846_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  or (_27215_, _17846_, _17845_);
  and (_17847_, _17072_, _24051_);
  and (_17848_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  or (_27287_, _17848_, _17847_);
  and (_17849_, _03269_, _23583_);
  and (_17850_, _03271_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  or (_27168_, _17850_, _17849_);
  and (_17851_, _03001_, _24219_);
  and (_17852_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_27214_, _17852_, _17851_);
  and (_17854_, _01810_, _23548_);
  and (_17855_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  or (_10090_, _17855_, _17854_);
  and (_17856_, _17391_, _24219_);
  and (_17857_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  or (_10093_, _17857_, _17856_);
  and (_17858_, _17072_, _23996_);
  and (_17859_, _17074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  or (_27288_, _17859_, _17858_);
  and (_17860_, _03001_, _23996_);
  and (_17861_, _03003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_10097_, _17861_, _17860_);
  and (_17862_, _00308_, _24636_);
  nand (_17863_, _17862_, _23504_);
  or (_17864_, _17862_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_17865_, _17864_, _25684_);
  and (_17866_, _17865_, _17863_);
  or (_17867_, _17866_, _25833_);
  and (_10102_, _17867_, _22731_);
  and (_17868_, _01810_, _23996_);
  and (_17869_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  or (_10111_, _17869_, _17868_);
  and (_17870_, _17391_, _23548_);
  and (_17871_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  or (_10113_, _17871_, _17870_);
  and (_17872_, _17110_, _24219_);
  and (_17873_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  or (_10115_, _17873_, _17872_);
  and (_17874_, _00308_, _24533_);
  nand (_17875_, _17874_, _23504_);
  or (_17876_, _17874_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_17877_, _17876_, _25684_);
  and (_17878_, _17877_, _17875_);
  or (_17879_, _17878_, _25686_);
  and (_10118_, _17879_, _22731_);
  and (_17880_, _00308_, _24607_);
  nand (_17881_, _17880_, _23504_);
  or (_17882_, _17880_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_17883_, _17882_, _25684_);
  and (_17884_, _17883_, _17881_);
  nor (_17885_, _25684_, _24043_);
  or (_17886_, _17885_, _17884_);
  and (_10120_, _17886_, _22731_);
  and (_17887_, _17110_, _23887_);
  and (_17888_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  or (_10126_, _17888_, _17887_);
  or (_17889_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_17890_, _23382_, _23380_);
  not (_17891_, _23051_);
  nand (_17892_, _23380_, _17891_);
  and (_17893_, _17892_, _22995_);
  and (_17894_, _17893_, _17890_);
  nand (_17895_, _23427_, _23392_);
  or (_17896_, _23427_, _23053_);
  and (_17897_, _17896_, _23390_);
  and (_17898_, _17897_, _17895_);
  and (_17899_, _23528_, _23120_);
  and (_17900_, _17899_, _23323_);
  and (_17901_, _01104_, _26163_);
  and (_17902_, _17901_, _01258_);
  nand (_17903_, _17902_, _17900_);
  nand (_17904_, _17903_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_17905_, _17904_, _17898_);
  nor (_17906_, _17905_, _17894_);
  nand (_17907_, _17906_, _00788_);
  or (_17908_, _00364_, _26560_);
  or (_17909_, _17908_, _00449_);
  or (_17910_, _17909_, _00530_);
  or (_17911_, _00715_, _00627_);
  or (_17912_, _17911_, _17910_);
  and (_17913_, _17912_, _23531_);
  or (_17914_, _17913_, _17907_);
  or (_17915_, _17914_, _00862_);
  and (_17916_, _17915_, _17889_);
  or (_17917_, _17916_, _00308_);
  and (_17918_, _02578_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_17919_, _17918_, _02580_);
  or (_17920_, _17919_, _00309_);
  and (_17921_, _17920_, _17917_);
  or (_17923_, _17921_, _25683_);
  or (_17924_, _25684_, _23880_);
  and (_17925_, _17924_, _22731_);
  and (_10130_, _17925_, _17923_);
  and (_17926_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_17927_, _17926_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_17928_, _23376_, _22995_);
  and (_17929_, _23413_, _23390_);
  nand (_17930_, _23484_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_17931_, _17930_, _17926_);
  or (_17932_, _17931_, _17929_);
  or (_17933_, _17932_, _17928_);
  and (_17934_, _17933_, _17927_);
  or (_17935_, _17934_, _00308_);
  or (_17936_, _24594_, _00546_);
  nand (_17937_, _17936_, _00308_);
  or (_17938_, _17937_, _03798_);
  and (_17939_, _17938_, _17935_);
  or (_17940_, _17939_, _25683_);
  nand (_17941_, _25683_, _24126_);
  and (_17943_, _17941_, _22731_);
  and (_10132_, _17943_, _17940_);
  and (_17944_, _17391_, _23887_);
  and (_17945_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  or (_26897_, _17945_, _17944_);
  and (_17946_, _17110_, _23583_);
  and (_17947_, _17112_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  or (_10140_, _17947_, _17946_);
  and (_17948_, _17391_, _23583_);
  and (_17949_, _17393_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  or (_10144_, _17949_, _17948_);
  and (_10147_, _03857_, _22731_);
  and (_17950_, _16008_, _23548_);
  and (_17951_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  or (_10151_, _17951_, _17950_);
  and (_17952_, _11441_, _24219_);
  and (_17953_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or (_10154_, _17953_, _17952_);
  and (_17954_, _00308_, _24177_);
  nand (_17955_, _17954_, _23504_);
  or (_17957_, _17954_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_17958_, _17957_, _25684_);
  and (_17959_, _17958_, _17955_);
  nor (_17960_, _25684_, _23542_);
  or (_17961_, _17960_, _17959_);
  and (_10161_, _17961_, _22731_);
  and (_17962_, _16731_, _24219_);
  and (_17963_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  or (_27222_, _17963_, _17962_);
  and (_17964_, _17385_, _24219_);
  and (_17965_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  or (_10166_, _17965_, _17964_);
  and (_17966_, _16008_, _24219_);
  and (_17967_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  or (_26960_, _17967_, _17966_);
  and (_17968_, _17102_, _23996_);
  and (_17969_, _17104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_27294_, _17969_, _17968_);
  and (_17970_, _17385_, _23887_);
  and (_17971_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  or (_10170_, _17971_, _17970_);
  and (_17972_, _17066_, _24219_);
  and (_17973_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_10173_, _17973_, _17972_);
  and (_17974_, _03275_, _24051_);
  and (_17975_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  or (_10175_, _17975_, _17974_);
  and (_17976_, _16731_, _23583_);
  and (_17977_, _16733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  or (_10177_, _17977_, _17976_);
  and (_17978_, _17385_, _24089_);
  and (_17979_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  or (_10179_, _17979_, _17978_);
  and (_17980_, _16541_, _23583_);
  and (_17981_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  or (_10181_, _17981_, _17980_);
  and (_17982_, _17066_, _23548_);
  and (_17983_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  or (_27295_, _17983_, _17982_);
  and (_17984_, _16541_, _24219_);
  and (_17985_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  or (_27224_, _17985_, _17984_);
  and (_17986_, _17066_, _23583_);
  and (_17987_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  or (_10186_, _17987_, _17986_);
  and (_17988_, _17385_, _24051_);
  and (_17989_, _17387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  or (_26901_, _17989_, _17988_);
  and (_17990_, _16541_, _24134_);
  and (_17991_, _16543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  or (_10190_, _17991_, _17990_);
  and (_17992_, _16008_, _24089_);
  and (_17993_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  or (_10194_, _17993_, _17992_);
  and (_17994_, _17066_, _24089_);
  and (_17995_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  or (_10196_, _17995_, _17994_);
  and (_17996_, _07038_, _24134_);
  and (_17997_, _07041_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  or (_10198_, _17997_, _17996_);
  and (_17999_, _17379_, _23548_);
  and (_18000_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  or (_10201_, _18000_, _17999_);
  and (_18001_, _04920_, _24089_);
  and (_18002_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  or (_10214_, _18002_, _18001_);
  nor (_10220_, _03809_, rst);
  and (_18003_, _17066_, _24051_);
  and (_18004_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  or (_10242_, _18004_, _18003_);
  and (_18005_, _04920_, _23548_);
  and (_18006_, _04923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  or (_10244_, _18006_, _18005_);
  and (_18007_, _16008_, _23583_);
  and (_18008_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  or (_26961_, _18008_, _18007_);
  and (_18009_, _17379_, _23583_);
  and (_18010_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  or (_26902_, _18010_, _18009_);
  and (_18011_, _17066_, _23996_);
  and (_18012_, _17068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_10260_, _18012_, _18011_);
  and (_10266_, _03732_, _22731_);
  nor (_10304_, _03721_, rst);
  and (_10324_, _03792_, _22731_);
  and (_18013_, _17379_, _24089_);
  and (_18014_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  or (_10337_, _18014_, _18013_);
  and (_10358_, _03779_, _22731_);
  and (_18015_, _02970_, _24089_);
  and (_18016_, _02972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  or (_10366_, _18016_, _18015_);
  and (_18017_, _03275_, _23996_);
  and (_18018_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_27165_, _18018_, _18017_);
  and (_18019_, _17379_, _23996_);
  and (_18020_, _17381_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_10375_, _18020_, _18019_);
  and (_18021_, _17058_, _23548_);
  and (_18022_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  or (_10379_, _18022_, _18021_);
  and (_18023_, _16034_, _24089_);
  and (_18024_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  or (_10420_, _18024_, _18023_);
  and (_18025_, _17369_, _24219_);
  and (_18026_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_10428_, _18026_, _18025_);
  and (_18027_, _16066_, _23583_);
  and (_18028_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  or (_10431_, _18028_, _18027_);
  and (_18029_, _16066_, _24089_);
  and (_18030_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  or (_10434_, _18030_, _18029_);
  nor (_10442_, _03759_, rst);
  and (_18031_, _17058_, _23887_);
  and (_18032_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  or (_10446_, _18032_, _18031_);
  and (_10454_, _03746_, _22731_);
  and (_18033_, _17369_, _23887_);
  and (_18034_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  or (_10461_, _18034_, _18033_);
  and (_18035_, _17058_, _24089_);
  and (_18036_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  or (_27296_, _18036_, _18035_);
  and (_18037_, _16704_, _24219_);
  and (_18038_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or (_27234_, _18038_, _18037_);
  and (_18039_, _16513_, _23548_);
  and (_18040_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  or (_10506_, _18040_, _18039_);
  and (_18041_, _17058_, _24134_);
  and (_18042_, _17060_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  or (_10508_, _18042_, _18041_);
  and (_18043_, _16773_, _23887_);
  and (_18044_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  or (_10513_, _18044_, _18043_);
  and (_18045_, _17369_, _23583_);
  and (_18046_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  or (_10523_, _18046_, _18045_);
  and (_18047_, _17369_, _24134_);
  and (_18048_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  or (_10528_, _18048_, _18047_);
  and (_18049_, _17052_, _24219_);
  and (_18050_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  or (_10534_, _18050_, _18049_);
  and (_18051_, _16513_, _23583_);
  and (_18052_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  or (_10539_, _18052_, _18051_);
  and (_18053_, _16121_, _23887_);
  and (_18054_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  or (_10551_, _18054_, _18053_);
  and (_18055_, _17369_, _23996_);
  and (_18056_, _17371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_26905_, _18056_, _18055_);
  and (_18057_, _03360_, _23548_);
  and (_18058_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  or (_10560_, _18058_, _18057_);
  and (_18059_, _17052_, _23548_);
  and (_18060_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  or (_10562_, _18060_, _18059_);
  and (_18061_, _16513_, _24051_);
  and (_18062_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  or (_10569_, _18062_, _18061_);
  and (_18063_, _17363_, _23548_);
  and (_18064_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  or (_10572_, _18064_, _18063_);
  and (_18065_, _16698_, _24051_);
  and (_18066_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  or (_10574_, _18066_, _18065_);
  and (_18067_, _16121_, _23548_);
  and (_18068_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  or (_10577_, _18068_, _18067_);
  and (_18069_, _17052_, _23583_);
  and (_18070_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  or (_10583_, _18070_, _18069_);
  and (_18071_, _15888_, _23583_);
  and (_18072_, _15890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  or (_10589_, _18072_, _18071_);
  and (_18073_, _17052_, _24051_);
  and (_18074_, _17054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  or (_27298_, _18074_, _18073_);
  and (_18075_, _16513_, _24134_);
  and (_18076_, _16515_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  or (_26935_, _18076_, _18075_);
  and (_18077_, _16698_, _24089_);
  and (_18078_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  or (_10599_, _18078_, _18077_);
  and (_18079_, _17363_, _23887_);
  and (_18080_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  or (_10601_, _18080_, _18079_);
  and (_18081_, _17046_, _24219_);
  and (_18082_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_10607_, _18082_, _18081_);
  and (_18083_, _09774_, _23887_);
  and (_18084_, _09777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  or (_10609_, _18084_, _18083_);
  and (_18085_, _16121_, _24219_);
  and (_18086_, _16123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_10613_, _18086_, _18085_);
  and (_18087_, _17363_, _24051_);
  and (_18088_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  or (_10618_, _18088_, _18087_);
  and (_18089_, _02617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_18090_, _02260_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_18091_, _18090_, _02284_);
  and (_18092_, _02283_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_18093_, _18092_, _02263_);
  or (_18094_, _18093_, _18091_);
  nor (_18095_, _02248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_18096_, _18095_, _02615_);
  nand (_18097_, _18096_, _18094_);
  nor (_18098_, _18097_, _02616_);
  or (_18099_, _18098_, _18089_);
  and (_18100_, _18099_, _02295_);
  and (_18101_, _02440_, _02450_);
  or (_10620_, _18101_, _18100_);
  and (_18102_, _11441_, _23887_);
  and (_18103_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  or (_10622_, _18103_, _18102_);
  and (_18104_, _17363_, _23996_);
  and (_18106_, _17365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  or (_10624_, _18106_, _18104_);
  and (_18107_, _08578_, _24089_);
  and (_18108_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  or (_10630_, _18108_, _18107_);
  and (_18109_, _16494_, _23548_);
  and (_18110_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  or (_10639_, _18110_, _18109_);
  and (_18111_, _16494_, _23583_);
  and (_18112_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  or (_26936_, _18112_, _18111_);
  and (_18113_, _17046_, _23548_);
  and (_18114_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  or (_27299_, _18114_, _18113_);
  and (_18115_, _17344_, _24219_);
  and (_18116_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  or (_10645_, _18116_, _18115_);
  and (_18117_, _16494_, _24051_);
  and (_18118_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  or (_10648_, _18118_, _18117_);
  and (_18120_, _06129_, _24134_);
  and (_18121_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  or (_10650_, _18121_, _18120_);
  and (_18122_, _03309_, _23996_);
  and (_18123_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  or (_10653_, _18123_, _18122_);
  and (_18124_, _17046_, _23583_);
  and (_18125_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  or (_10656_, _18125_, _18124_);
  and (_18126_, _06129_, _23583_);
  and (_18127_, _06131_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  or (_10658_, _18127_, _18126_);
  and (_18128_, _11441_, _23583_);
  and (_18129_, _11444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  or (_10668_, _18129_, _18128_);
  and (_18130_, _17046_, _24051_);
  and (_18131_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  or (_10671_, _18131_, _18130_);
  and (_18132_, _25658_, _24089_);
  and (_18133_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  or (_10675_, _18133_, _18132_);
  and (_18135_, _17344_, _23548_);
  and (_18136_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  or (_26906_, _18136_, _18135_);
  and (_18137_, _25658_, _23548_);
  and (_18138_, _25660_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  or (_10681_, _18138_, _18137_);
  and (_18139_, _17344_, _23583_);
  and (_18140_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  or (_26908_, _18140_, _18139_);
  and (_18141_, _24497_, _24089_);
  and (_18142_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  or (_10686_, _18142_, _18141_);
  and (_18143_, _17046_, _23996_);
  and (_18144_, _17048_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_10688_, _18144_, _18143_);
  and (_18145_, _05485_, _23548_);
  and (_18146_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  or (_10690_, _18146_, _18145_);
  and (_18147_, _16494_, _24134_);
  and (_18148_, _16496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  or (_10692_, _18148_, _18147_);
  and (_18149_, _16034_, _23996_);
  and (_18150_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  or (_10694_, _18150_, _18149_);
  and (_18151_, _17344_, _24089_);
  and (_18152_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  or (_10696_, _18152_, _18151_);
  and (_18153_, _17042_, _24219_);
  and (_18154_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_27300_, _18154_, _18153_);
  and (_18156_, _03275_, _23548_);
  and (_18157_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  or (_10703_, _18157_, _18156_);
  and (_18158_, _03275_, _24219_);
  and (_18159_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_10705_, _18159_, _18158_);
  and (_18160_, _16698_, _23996_);
  and (_18161_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  or (_10711_, _18161_, _18160_);
  and (_18162_, _24497_, _23996_);
  and (_18163_, _24500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  or (_10713_, _18163_, _18162_);
  and (_18164_, _16698_, _24134_);
  and (_18165_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  or (_10716_, _18165_, _18164_);
  and (_18166_, _17344_, _24051_);
  and (_18167_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  or (_26909_, _18167_, _18166_);
  and (_18168_, _17042_, _23887_);
  and (_18169_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  or (_10720_, _18169_, _18168_);
  and (_18170_, _16476_, _24219_);
  and (_18171_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_10723_, _18171_, _18170_);
  and (_18172_, _16476_, _23548_);
  and (_18173_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  or (_10734_, _18173_, _18172_);
  and (_18174_, _08578_, _23583_);
  and (_18175_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  or (_10736_, _18175_, _18174_);
  and (_18177_, _16066_, _24134_);
  and (_18178_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  or (_10739_, _18178_, _18177_);
  and (_18179_, _17344_, _24134_);
  and (_18180_, _17346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  or (_10747_, _18180_, _18179_);
  and (_18181_, _17042_, _23583_);
  and (_18182_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  or (_27302_, _18182_, _18181_);
  and (_18183_, _25124_, _25481_);
  nand (_18184_, _18183_, _23504_);
  or (_18185_, _18183_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_18186_, _18185_, _24539_);
  and (_18187_, _18186_, _18184_);
  nand (_18188_, _25130_, _23989_);
  or (_18189_, _25130_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_18190_, _18189_, _24179_);
  and (_18191_, _18190_, _18188_);
  nor (_18192_, _24178_, _04206_);
  or (_18193_, _18192_, rst);
  or (_18194_, _18193_, _18191_);
  or (_10753_, _18194_, _18187_);
  and (_18195_, _17042_, _24134_);
  and (_18196_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  or (_27303_, _18196_, _18195_);
  and (_18197_, _16066_, _23996_);
  and (_18198_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or (_26959_, _18198_, _18197_);
  and (_18199_, _17338_, _24219_);
  and (_18200_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_26911_, _18200_, _18199_);
  and (_18201_, _16476_, _23887_);
  and (_18202_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  or (_26938_, _18202_, _18201_);
  and (_18203_, _16476_, _24089_);
  and (_18204_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  or (_26939_, _18204_, _18203_);
  and (_18205_, _17338_, _23887_);
  and (_18206_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  or (_26912_, _18206_, _18205_);
  and (_18207_, _11419_, _24089_);
  and (_18208_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  or (_27087_, _18208_, _18207_);
  and (_18209_, _16476_, _24134_);
  and (_18210_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  or (_26940_, _18210_, _18209_);
  and (_18211_, _17042_, _23996_);
  and (_18212_, _17044_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_27304_, _18212_, _18211_);
  and (_18213_, _03043_, _23583_);
  and (_18214_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  or (_27251_, _18214_, _18213_);
  and (_18215_, _17338_, _24089_);
  and (_18216_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  or (_26914_, _18216_, _18215_);
  and (_18217_, _17545_, _23583_);
  and (_18218_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  or (_27254_, _18218_, _18217_);
  and (_18219_, _17036_, _24219_);
  and (_18220_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  or (_27305_, _18220_, _18219_);
  and (_18221_, _17545_, _24219_);
  and (_18222_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or (_27253_, _18222_, _18221_);
  and (_18223_, _16476_, _23996_);
  and (_18224_, _16478_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_26941_, _18224_, _18223_);
  and (_18225_, _17036_, _23887_);
  and (_18226_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  or (_27306_, _18226_, _18225_);
  and (_18227_, _16468_, _24219_);
  and (_18228_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_26942_, _18228_, _18227_);
  and (_18229_, _17338_, _24051_);
  and (_18230_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  or (_26915_, _18230_, _18229_);
  and (_18231_, _16773_, _23996_);
  and (_18232_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  or (_27239_, _18232_, _18231_);
  and (_18233_, _11419_, _23583_);
  and (_18234_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  or (_27086_, _18234_, _18233_);
  and (_18235_, _17338_, _23996_);
  and (_18236_, _17340_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_26916_, _18236_, _18235_);
  and (_18237_, _17036_, _24089_);
  and (_18238_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  or (_27307_, _18238_, _18237_);
  and (_18239_, _16468_, _23548_);
  and (_18240_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  or (_26943_, _18240_, _18239_);
  and (_18241_, _16773_, _24134_);
  and (_18242_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  or (_27238_, _18242_, _18241_);
  and (_18243_, _17334_, _24219_);
  and (_18244_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_26918_, _18244_, _18243_);
  and (_18245_, _11419_, _23887_);
  and (_18246_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  or (_27085_, _18246_, _18245_);
  and (_18247_, _17036_, _24051_);
  and (_18248_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  or (_27308_, _18248_, _18247_);
  and (_18249_, _16468_, _23583_);
  and (_18250_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  or (_26944_, _18250_, _18249_);
  and (_18251_, _17334_, _23887_);
  and (_18252_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  or (_26919_, _18252_, _18251_);
  and (_18253_, _16773_, _24051_);
  and (_18254_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  or (_27237_, _18254_, _18253_);
  and (_18255_, _10867_, _23583_);
  and (_18256_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  or (_27261_, _18256_, _18255_);
  and (_18257_, _08578_, _23887_);
  and (_18258_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  or (_27077_, _18258_, _18257_);
  and (_18259_, _16468_, _24051_);
  and (_18260_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  or (_26945_, _18260_, _18259_);
  and (_18261_, _03275_, _23583_);
  and (_18262_, _03277_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  or (_10810_, _18262_, _18261_);
  and (_18263_, _17036_, _24134_);
  and (_18264_, _17038_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  or (_10812_, _18264_, _18263_);
  and (_18265_, _17334_, _23583_);
  and (_18266_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  or (_26920_, _18266_, _18265_);
  and (_18268_, _02996_, _23548_);
  and (_18269_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  or (_10818_, _18269_, _18268_);
  and (_18270_, _10867_, _24134_);
  and (_18271_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  or (_10820_, _18271_, _18270_);
  and (_18272_, _16468_, _24134_);
  and (_18273_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  or (_26946_, _18273_, _18272_);
  and (_18274_, _16468_, _23996_);
  and (_18275_, _16470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_10826_, _18275_, _18274_);
  and (_18276_, _16014_, _24089_);
  and (_18277_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  or (_10828_, _18277_, _18276_);
  and (_18278_, _16014_, _24134_);
  and (_18279_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  or (_10831_, _18279_, _18278_);
  and (_18280_, _16773_, _24089_);
  and (_18281_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  or (_10833_, _18281_, _18280_);
  and (_18282_, _24394_, _24219_);
  and (_18283_, _24396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_10838_, _18283_, _18282_);
  and (_18284_, _25018_, _25481_);
  nand (_18285_, _18284_, _23504_);
  or (_18286_, _18284_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_18287_, _18286_, _24539_);
  and (_18288_, _18287_, _18285_);
  nand (_18289_, _25026_, _23989_);
  or (_18290_, _25026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_18291_, _18290_, _24179_);
  and (_18292_, _18291_, _18289_);
  nor (_18293_, _24178_, _04146_);
  or (_18294_, _18293_, rst);
  or (_18295_, _18294_, _18292_);
  or (_10842_, _18295_, _18288_);
  and (_18296_, _11311_, _24051_);
  and (_18297_, _11313_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  or (_10844_, _18297_, _18296_);
  and (_18298_, _05465_, _23548_);
  and (_18299_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  or (_27067_, _18299_, _18298_);
  and (_18300_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_18301_, _26724_, _22737_);
  or (_18302_, _18301_, _18300_);
  or (_18303_, _18302_, _02359_);
  and (_26848_[2], _18303_, _22731_);
  and (_18304_, _23890_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_18305_, _23784_, _23824_);
  or (_18306_, _04793_, _04795_);
  or (_18307_, _18306_, _18305_);
  or (_18308_, _26703_, _23828_);
  or (_18309_, _18308_, _17182_);
  or (_18310_, _18309_, _18307_);
  or (_18311_, _18310_, _11472_);
  and (_18312_, _18311_, _23855_);
  or (_26847_[1], _18312_, _18304_);
  and (_18313_, _17581_, _23548_);
  and (_18314_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  or (_10853_, _18314_, _18313_);
  or (_18315_, _23724_, _26679_);
  or (_18316_, _22736_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_18317_, _18316_, _22731_);
  and (_26844_[7], _18317_, _18315_);
  and (_18318_, _25220_, _25481_);
  nand (_18319_, _18318_, _23504_);
  or (_18320_, _18318_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_18321_, _18320_, _24539_);
  and (_18322_, _18321_, _18319_);
  nand (_18323_, _25228_, _23989_);
  or (_18324_, _25228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_18325_, _18324_, _24179_);
  and (_18326_, _18325_, _18323_);
  nor (_18327_, _24178_, _04001_);
  or (_18328_, _18327_, rst);
  or (_18329_, _18328_, _18326_);
  or (_10857_, _18329_, _18322_);
  and (_18330_, _16014_, _24051_);
  and (_18331_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  or (_10864_, _18331_, _18330_);
  and (_18332_, _10867_, _23996_);
  and (_18333_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  or (_10866_, _18333_, _18332_);
  and (_18334_, _25319_, _25481_);
  nand (_18335_, _18334_, _23504_);
  or (_18336_, _18334_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_18337_, _18336_, _24539_);
  and (_18338_, _18337_, _18335_);
  nand (_18339_, _25327_, _23989_);
  or (_18340_, _25327_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_18341_, _18340_, _24179_);
  and (_18342_, _18341_, _18339_);
  nor (_18343_, _24178_, _03944_);
  or (_18344_, _18343_, rst);
  or (_18345_, _18344_, _18342_);
  or (_10870_, _18345_, _18338_);
  and (_18346_, _16698_, _24219_);
  and (_18347_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  or (_10881_, _18347_, _18346_);
  and (_18348_, _16698_, _23887_);
  and (_18349_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  or (_10883_, _18349_, _18348_);
  and (_18350_, _17581_, _24219_);
  and (_18351_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  or (_27218_, _18351_, _18350_);
  and (_18352_, _11419_, _24134_);
  and (_18353_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  or (_10886_, _18353_, _18352_);
  and (_18354_, _16698_, _23548_);
  and (_18355_, _16700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  or (_27240_, _18355_, _18354_);
  and (_18356_, _11419_, _23996_);
  and (_18357_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_10891_, _18357_, _18356_);
  and (_18358_, _03281_, _24051_);
  and (_18359_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  or (_10893_, _18359_, _18358_);
  and (_18360_, _16670_, _23996_);
  and (_18361_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  or (_10897_, _18361_, _18360_);
  and (_18362_, _03360_, _23887_);
  and (_18363_, _03362_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  or (_10899_, _18363_, _18362_);
  and (_18364_, _10867_, _24219_);
  and (_18365_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  or (_10901_, _18365_, _18364_);
  and (_18366_, _25414_, _23996_);
  and (_18367_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_10910_, _18367_, _18366_);
  and (_18368_, _03281_, _24089_);
  and (_18369_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  or (_10915_, _18369_, _18368_);
  and (_18370_, _08578_, _24051_);
  and (_18371_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  or (_10918_, _18371_, _18370_);
  and (_18372_, _16034_, _24134_);
  and (_18373_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  or (_10921_, _18373_, _18372_);
  and (_18374_, _16066_, _24219_);
  and (_18375_, _16068_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or (_10923_, _18375_, _18374_);
  and (_18376_, _08578_, _24134_);
  and (_18377_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  or (_10925_, _18377_, _18376_);
  and (_18378_, _02996_, _23887_);
  and (_18379_, _02998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  or (_10928_, _18379_, _18378_);
  and (_18380_, _24142_, _24089_);
  and (_18381_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  or (_10933_, _18381_, _18380_);
  and (_18382_, _25414_, _24134_);
  and (_18383_, _25416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  or (_10936_, _18383_, _18382_);
  and (_18384_, _24089_, _22983_);
  and (_18385_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  or (_10938_, _18385_, _18384_);
  and (_18386_, _16704_, _23996_);
  and (_18387_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or (_10941_, _18387_, _18386_);
  and (_18388_, _24099_, _23548_);
  and (_18389_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  or (_10942_, _18389_, _18388_);
  and (_18390_, _24160_, _24051_);
  and (_18391_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  or (_10944_, _18391_, _18390_);
  and (_18392_, _24160_, _23583_);
  and (_18393_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  or (_26922_, _18393_, _18392_);
  and (_18394_, _17032_, _23996_);
  and (_18395_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  or (_10946_, _18395_, _18394_);
  and (_18396_, _24219_, _22983_);
  and (_18397_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  or (_10948_, _18397_, _18396_);
  and (_18398_, _16014_, _23996_);
  and (_18399_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or (_26958_, _18399_, _18398_);
  and (_18400_, _24320_, _23887_);
  and (_18401_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  or (_10950_, _18401_, _18400_);
  and (_18402_, _24160_, _24089_);
  and (_18403_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  or (_10951_, _18403_, _18402_);
  and (_18404_, _24219_, _24099_);
  and (_18405_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_10953_, _18405_, _18404_);
  and (_18406_, _23996_, _22983_);
  and (_18407_, _23550_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  or (_10955_, _18407_, _18406_);
  and (_18408_, _16704_, _24134_);
  and (_18409_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  or (_10958_, _18409_, _18408_);
  and (_18410_, _24219_, _24147_);
  and (_18411_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_10964_, _18411_, _18410_);
  and (_18412_, _24142_, _23996_);
  and (_18413_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  or (_10967_, _18413_, _18412_);
  and (_18414_, _24057_, _23583_);
  and (_18415_, _24092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  or (_10968_, _18415_, _18414_);
  and (_18416_, _03309_, _23887_);
  and (_18417_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  or (_10970_, _18417_, _18416_);
  and (_18418_, _16704_, _24051_);
  and (_18419_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  or (_27235_, _18419_, _18418_);
  and (_18420_, _25637_, _23887_);
  and (_18421_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  or (_10974_, _18421_, _18420_);
  and (_18422_, _24099_, _24051_);
  and (_18423_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  or (_10976_, _18423_, _18422_);
  and (_18424_, _24219_, _24142_);
  and (_18425_, _24144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  or (_10978_, _18425_, _18424_);
  and (_18426_, _24160_, _24134_);
  and (_18427_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  or (_10980_, _18427_, _18426_);
  and (_18428_, _03281_, _24134_);
  and (_18429_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  or (_10982_, _18429_, _18428_);
  and (_18430_, _24099_, _23887_);
  and (_18431_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  or (_10984_, _18431_, _18430_);
  and (_18432_, _24320_, _24051_);
  and (_18433_, _24322_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  or (_27279_, _18433_, _18432_);
  and (_18434_, _24160_, _23996_);
  and (_18435_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  or (_10993_, _18435_, _18434_);
  and (_18436_, _24099_, _23583_);
  and (_18437_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  or (_10995_, _18437_, _18436_);
  and (_18438_, _24224_, _24089_);
  and (_18439_, _24226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  or (_27283_, _18439_, _18438_);
  and (_18440_, _10867_, _23548_);
  and (_18442_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  or (_10999_, _18442_, _18440_);
  and (_18443_, _05465_, _23996_);
  and (_18444_, _05468_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  or (_11001_, _18444_, _18443_);
  and (_18445_, _24099_, _24089_);
  and (_18446_, _24137_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  or (_11005_, _18446_, _18445_);
  and (_26840_[1], _23660_, _22731_);
  and (_18447_, _24147_, _24134_);
  and (_18448_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  or (_11011_, _18448_, _18447_);
  and (_18449_, _10867_, _23887_);
  and (_18450_, _10869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  or (_11014_, _18450_, _18449_);
  and (_18451_, _24373_, _23996_);
  and (_18452_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_11017_, _18452_, _18451_);
  and (_18453_, _16014_, _24219_);
  and (_18454_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_11021_, _18454_, _18453_);
  and (_18455_, _17032_, _24089_);
  and (_18456_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  or (_11023_, _18456_, _18455_);
  and (_18457_, _17032_, _24134_);
  and (_18458_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  or (_11024_, _18458_, _18457_);
  nand (_18459_, _02623_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_18460_, _18459_, _16094_);
  not (_18461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_18462_, _06162_, _18461_);
  and (_18463_, _06162_, _18461_);
  or (_18464_, _18463_, _18462_);
  or (_18465_, _18464_, _02617_);
  nand (_18466_, _02617_, _18461_);
  and (_18467_, _18466_, _18465_);
  or (_18468_, _18467_, _18460_);
  and (_18469_, _18468_, _02295_);
  and (_18470_, _02440_, _02689_);
  or (_11027_, _18470_, _18469_);
  and (_18471_, _24219_, _24160_);
  and (_18472_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  or (_26921_, _18472_, _18471_);
  and (_18473_, _24160_, _23548_);
  and (_18474_, _24162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  or (_11030_, _18474_, _18473_);
  and (_18475_, _24155_, _24089_);
  and (_18476_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  or (_11036_, _18476_, _18475_);
  and (_18477_, _17032_, _24051_);
  and (_18478_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  or (_11039_, _18478_, _18477_);
  and (_18479_, _17334_, _24134_);
  and (_18480_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  or (_11042_, _18480_, _18479_);
  and (_18481_, _17032_, _23887_);
  and (_18482_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  or (_11043_, _18482_, _18481_);
  and (_18483_, _24373_, _24134_);
  and (_18484_, _24375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  or (_11048_, _18484_, _18483_);
  and (_18485_, _17334_, _23996_);
  and (_18486_, _17336_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_11050_, _18486_, _18485_);
  and (_18487_, _17032_, _23583_);
  and (_18488_, _17034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  or (_27309_, _18488_, _18487_);
  and (_18489_, _24147_, _23583_);
  and (_18490_, _24149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  or (_11056_, _18490_, _18489_);
  and (_18491_, _16014_, _23887_);
  and (_18492_, _16016_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  or (_26957_, _18492_, _18491_);
  and (_18493_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  and (_18494_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  or (_18495_, _18494_, _18493_);
  and (_18496_, _18495_, _09792_);
  and (_18497_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  and (_18498_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  or (_18499_, _18498_, _18497_);
  and (_18500_, _18499_, _05549_);
  or (_18501_, _18500_, _18496_);
  or (_18502_, _18501_, _09791_);
  and (_18503_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  and (_18504_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  or (_18505_, _18504_, _18503_);
  and (_18506_, _18505_, _09792_);
  and (_18507_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  and (_18508_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  or (_18509_, _18508_, _18507_);
  and (_18510_, _18509_, _05549_);
  or (_18511_, _18510_, _18506_);
  or (_18512_, _18511_, _05535_);
  and (_18513_, _18512_, _09805_);
  and (_18514_, _18513_, _18502_);
  or (_18515_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  or (_18516_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  and (_18517_, _18516_, _18515_);
  and (_18518_, _18517_, _09792_);
  or (_18519_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  or (_18520_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  and (_18521_, _18520_, _18519_);
  and (_18522_, _18521_, _05549_);
  or (_18523_, _18522_, _18518_);
  or (_18524_, _18523_, _09791_);
  or (_18525_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  or (_18526_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  and (_18527_, _18526_, _18525_);
  and (_18528_, _18527_, _09792_);
  or (_18529_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_18530_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  and (_18531_, _18530_, _18529_);
  and (_18532_, _18531_, _05549_);
  or (_18533_, _18532_, _18528_);
  or (_18534_, _18533_, _05535_);
  and (_18535_, _18534_, _05542_);
  and (_18536_, _18535_, _18524_);
  or (_18537_, _18536_, _18514_);
  and (_18538_, _18537_, _05518_);
  and (_18539_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  and (_18540_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_18541_, _18540_, _18539_);
  and (_18542_, _18541_, _09792_);
  and (_18543_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  and (_18544_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  or (_18545_, _18544_, _18543_);
  and (_18546_, _18545_, _05549_);
  or (_18547_, _18546_, _18542_);
  or (_18548_, _18547_, _09791_);
  and (_18549_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  and (_18550_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_18551_, _18550_, _18549_);
  and (_18552_, _18551_, _09792_);
  and (_18553_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  and (_18554_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  or (_18555_, _18554_, _18553_);
  and (_18556_, _18555_, _05549_);
  or (_18557_, _18556_, _18552_);
  or (_18558_, _18557_, _05535_);
  and (_18559_, _18558_, _09805_);
  and (_18560_, _18559_, _18548_);
  or (_18561_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_18562_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  and (_18563_, _18562_, _05549_);
  and (_18564_, _18563_, _18561_);
  or (_18565_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_18566_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  and (_18567_, _18566_, _09792_);
  and (_18568_, _18567_, _18565_);
  or (_18569_, _18568_, _18564_);
  or (_18570_, _18569_, _09791_);
  or (_18571_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  or (_18572_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  and (_18573_, _18572_, _05549_);
  and (_18574_, _18573_, _18571_);
  or (_18575_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  or (_18576_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  and (_18577_, _18576_, _09792_);
  and (_18578_, _18577_, _18575_);
  or (_18579_, _18578_, _18574_);
  or (_18580_, _18579_, _05535_);
  and (_18581_, _18580_, _05542_);
  and (_18582_, _18581_, _18570_);
  or (_18583_, _18582_, _18560_);
  and (_18584_, _18583_, _09850_);
  or (_18585_, _18584_, _18538_);
  and (_18586_, _18585_, _09790_);
  and (_18587_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_18588_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_18589_, _18588_, _18587_);
  and (_18590_, _18589_, _09792_);
  and (_18591_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_18592_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  or (_18593_, _18592_, _18591_);
  and (_18594_, _18593_, _05549_);
  or (_18595_, _18594_, _18590_);
  and (_18596_, _18595_, _05535_);
  and (_18597_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_18598_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or (_18599_, _18598_, _18597_);
  and (_18600_, _18599_, _09792_);
  and (_18601_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_18602_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  or (_18603_, _18602_, _18601_);
  and (_18604_, _18603_, _05549_);
  or (_18605_, _18604_, _18600_);
  and (_18606_, _18605_, _09791_);
  or (_18607_, _18606_, _18596_);
  and (_18608_, _18607_, _09805_);
  or (_18609_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_18610_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_18611_, _18610_, _05549_);
  and (_18612_, _18611_, _18609_);
  or (_18613_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_18614_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_18615_, _18614_, _09792_);
  and (_18616_, _18615_, _18613_);
  or (_18617_, _18616_, _18612_);
  and (_18618_, _18617_, _05535_);
  or (_18619_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_18620_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_18621_, _18620_, _05549_);
  and (_18622_, _18621_, _18619_);
  or (_18623_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_18624_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_18625_, _18624_, _09792_);
  and (_18626_, _18625_, _18623_);
  or (_18627_, _18626_, _18622_);
  and (_18628_, _18627_, _09791_);
  or (_18629_, _18628_, _18618_);
  and (_18630_, _18629_, _05542_);
  or (_18631_, _18630_, _18608_);
  and (_18632_, _18631_, _09850_);
  and (_18633_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  and (_18634_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  or (_18635_, _18634_, _18633_);
  and (_18636_, _18635_, _09792_);
  and (_18637_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  and (_18638_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  or (_18639_, _18638_, _18637_);
  and (_18640_, _18639_, _05549_);
  or (_18641_, _18640_, _18636_);
  and (_18642_, _18641_, _05535_);
  and (_18643_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  and (_18644_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  or (_18645_, _18644_, _18643_);
  and (_18646_, _18645_, _09792_);
  and (_18647_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  and (_18648_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  or (_18649_, _18648_, _18647_);
  and (_18650_, _18649_, _05549_);
  or (_18651_, _18650_, _18646_);
  and (_18652_, _18651_, _09791_);
  or (_18653_, _18652_, _18642_);
  and (_18654_, _18653_, _09805_);
  or (_18655_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  or (_18656_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  and (_18657_, _18656_, _18655_);
  and (_18658_, _18657_, _09792_);
  or (_18659_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  or (_18660_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  and (_18661_, _18660_, _18659_);
  and (_18662_, _18661_, _05549_);
  or (_18663_, _18662_, _18658_);
  and (_18664_, _18663_, _05535_);
  or (_18665_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  or (_18666_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  and (_18667_, _18666_, _18665_);
  and (_18668_, _18667_, _09792_);
  or (_18669_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_18670_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  and (_18671_, _18670_, _18669_);
  and (_18672_, _18671_, _05549_);
  or (_18673_, _18672_, _18668_);
  and (_18674_, _18673_, _09791_);
  or (_18675_, _18674_, _18664_);
  and (_18676_, _18675_, _05542_);
  or (_18677_, _18676_, _18654_);
  and (_18678_, _18677_, _05518_);
  or (_18679_, _18678_, _18632_);
  and (_18680_, _18679_, _05520_);
  or (_18681_, _18680_, _18586_);
  or (_18682_, _18681_, _05526_);
  and (_18683_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  and (_18684_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  or (_18685_, _18684_, _18683_);
  and (_18686_, _18685_, _09792_);
  and (_18687_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  and (_18688_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  or (_18689_, _18688_, _18687_);
  and (_18690_, _18689_, _05549_);
  or (_18691_, _18690_, _18686_);
  or (_18692_, _18691_, _09791_);
  and (_18693_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  and (_18694_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  or (_18695_, _18694_, _18693_);
  and (_18696_, _18695_, _09792_);
  and (_18697_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  and (_18698_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  or (_18699_, _18698_, _18697_);
  and (_18700_, _18699_, _05549_);
  or (_18701_, _18700_, _18696_);
  or (_18702_, _18701_, _05535_);
  and (_18703_, _18702_, _09805_);
  and (_18704_, _18703_, _18692_);
  or (_18705_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  or (_18706_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  and (_18707_, _18706_, _05549_);
  and (_18708_, _18707_, _18705_);
  or (_18709_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  or (_18710_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  and (_18711_, _18710_, _09792_);
  and (_18712_, _18711_, _18709_);
  or (_18713_, _18712_, _18708_);
  or (_18714_, _18713_, _09791_);
  or (_18715_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  or (_18716_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  and (_18717_, _18716_, _05549_);
  and (_18718_, _18717_, _18715_);
  or (_18719_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  or (_18720_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  and (_18721_, _18720_, _09792_);
  and (_18722_, _18721_, _18719_);
  or (_18723_, _18722_, _18718_);
  or (_18724_, _18723_, _05535_);
  and (_18725_, _18724_, _05542_);
  and (_18726_, _18725_, _18714_);
  or (_18727_, _18726_, _18704_);
  and (_18728_, _18727_, _09850_);
  and (_18729_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  and (_18730_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  or (_18731_, _18730_, _18729_);
  and (_18732_, _18731_, _09792_);
  and (_18733_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  and (_18734_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  or (_18735_, _18734_, _18733_);
  and (_18736_, _18735_, _05549_);
  or (_18737_, _18736_, _18732_);
  or (_18738_, _18737_, _09791_);
  and (_18739_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  and (_18740_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  or (_18741_, _18740_, _18739_);
  and (_18742_, _18741_, _09792_);
  and (_18743_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  and (_18744_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  or (_18745_, _18744_, _18743_);
  and (_18746_, _18745_, _05549_);
  or (_18747_, _18746_, _18742_);
  or (_18748_, _18747_, _05535_);
  and (_18749_, _18748_, _09805_);
  and (_18750_, _18749_, _18738_);
  or (_18751_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  or (_18752_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  and (_18753_, _18752_, _18751_);
  and (_18754_, _18753_, _09792_);
  or (_18755_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  or (_18756_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  and (_18757_, _18756_, _18755_);
  and (_18758_, _18757_, _05549_);
  or (_18759_, _18758_, _18754_);
  or (_18760_, _18759_, _09791_);
  or (_18761_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  or (_18762_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  and (_18763_, _18762_, _18761_);
  and (_18764_, _18763_, _09792_);
  or (_18765_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  or (_18766_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  and (_18767_, _18766_, _18765_);
  and (_18768_, _18767_, _05549_);
  or (_18769_, _18768_, _18764_);
  or (_18770_, _18769_, _05535_);
  and (_18771_, _18770_, _05542_);
  and (_18772_, _18771_, _18760_);
  or (_18773_, _18772_, _18750_);
  and (_18774_, _18773_, _05518_);
  or (_18775_, _18774_, _18728_);
  and (_18776_, _18775_, _09790_);
  or (_18777_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  or (_18778_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  and (_18779_, _18778_, _18777_);
  and (_18780_, _18779_, _09792_);
  or (_18781_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  or (_18782_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  and (_18783_, _18782_, _18781_);
  and (_18784_, _18783_, _05549_);
  or (_18785_, _18784_, _18780_);
  and (_18786_, _18785_, _09791_);
  or (_18787_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  or (_18788_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  and (_18789_, _18788_, _18787_);
  and (_18790_, _18789_, _09792_);
  or (_18791_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  or (_18792_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  and (_18793_, _18792_, _18791_);
  and (_18794_, _18793_, _05549_);
  or (_18795_, _18794_, _18790_);
  and (_18796_, _18795_, _05535_);
  or (_18797_, _18796_, _18786_);
  and (_18798_, _18797_, _05542_);
  and (_18799_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  and (_18800_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  or (_18801_, _18800_, _18799_);
  and (_18802_, _18801_, _09792_);
  and (_18803_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  and (_18804_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  or (_18805_, _18804_, _18803_);
  and (_18806_, _18805_, _05549_);
  or (_18807_, _18806_, _18802_);
  and (_18808_, _18807_, _09791_);
  and (_18809_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  and (_18810_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  or (_18811_, _18810_, _18809_);
  and (_18812_, _18811_, _09792_);
  and (_18813_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  and (_18814_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  or (_18815_, _18814_, _18813_);
  and (_18816_, _18815_, _05549_);
  or (_18817_, _18816_, _18812_);
  and (_18818_, _18817_, _05535_);
  or (_18819_, _18818_, _18808_);
  and (_18820_, _18819_, _09805_);
  or (_18821_, _18820_, _18798_);
  and (_18822_, _18821_, _05518_);
  or (_18823_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or (_18824_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  and (_18825_, _18824_, _05549_);
  and (_18826_, _18825_, _18823_);
  or (_18827_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  or (_18828_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  and (_18829_, _18828_, _09792_);
  and (_18830_, _18829_, _18827_);
  or (_18831_, _18830_, _18826_);
  and (_18832_, _18831_, _09791_);
  or (_18833_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  or (_18834_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  and (_18835_, _18834_, _05549_);
  and (_18836_, _18835_, _18833_);
  or (_18837_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  or (_18838_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  and (_18839_, _18838_, _09792_);
  and (_18840_, _18839_, _18837_);
  or (_18841_, _18840_, _18836_);
  and (_18842_, _18841_, _05535_);
  or (_18843_, _18842_, _18832_);
  and (_18844_, _18843_, _05542_);
  and (_18845_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  and (_18846_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  or (_18847_, _18846_, _18845_);
  and (_18848_, _18847_, _09792_);
  and (_18849_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  and (_18850_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  or (_18851_, _18850_, _18849_);
  and (_18852_, _18851_, _05549_);
  or (_18853_, _18852_, _18848_);
  and (_18854_, _18853_, _09791_);
  and (_18855_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  and (_18856_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  or (_18857_, _18856_, _18855_);
  and (_18858_, _18857_, _09792_);
  and (_18859_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  and (_18860_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  or (_18861_, _18860_, _18859_);
  and (_18862_, _18861_, _05549_);
  or (_18863_, _18862_, _18858_);
  and (_18864_, _18863_, _05535_);
  or (_18865_, _18864_, _18854_);
  and (_18866_, _18865_, _09805_);
  or (_18867_, _18866_, _18844_);
  and (_18868_, _18867_, _09850_);
  or (_18869_, _18868_, _18822_);
  and (_18870_, _18869_, _05520_);
  or (_18871_, _18870_, _18776_);
  or (_18872_, _18871_, _10033_);
  and (_18873_, _18872_, _18682_);
  or (_18874_, _18873_, _00143_);
  and (_18875_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  and (_18876_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  or (_18877_, _18876_, _18875_);
  and (_18878_, _18877_, _09792_);
  and (_18879_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  and (_18880_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  or (_18881_, _18880_, _18879_);
  and (_18882_, _18881_, _05549_);
  or (_18883_, _18882_, _18878_);
  or (_18884_, _18883_, _09791_);
  and (_18885_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  and (_18886_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  or (_18887_, _18886_, _18885_);
  and (_18888_, _18887_, _09792_);
  and (_18889_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  and (_18890_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  or (_18891_, _18890_, _18889_);
  and (_18892_, _18891_, _05549_);
  or (_18893_, _18892_, _18888_);
  or (_18894_, _18893_, _05535_);
  and (_18895_, _18894_, _09805_);
  and (_18896_, _18895_, _18884_);
  or (_18897_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  or (_18898_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  and (_18899_, _18898_, _18897_);
  and (_18900_, _18899_, _09792_);
  or (_18901_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  or (_18902_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  and (_18903_, _18902_, _18901_);
  and (_18904_, _18903_, _05549_);
  or (_18905_, _18904_, _18900_);
  or (_18906_, _18905_, _09791_);
  or (_18907_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  or (_18908_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  and (_18909_, _18908_, _18907_);
  and (_18910_, _18909_, _09792_);
  or (_18911_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  or (_18912_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  and (_18913_, _18912_, _18911_);
  and (_18914_, _18913_, _05549_);
  or (_18915_, _18914_, _18910_);
  or (_18916_, _18915_, _05535_);
  and (_18917_, _18916_, _05542_);
  and (_18918_, _18917_, _18906_);
  or (_18919_, _18918_, _18896_);
  and (_18920_, _18919_, _05518_);
  and (_18921_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  and (_18922_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  or (_18923_, _18922_, _18921_);
  and (_18924_, _18923_, _09792_);
  and (_18925_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  and (_18926_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  or (_18927_, _18926_, _18925_);
  and (_18928_, _18927_, _05549_);
  or (_18929_, _18928_, _18924_);
  or (_18930_, _18929_, _09791_);
  and (_18931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  and (_18932_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  or (_18933_, _18932_, _18931_);
  and (_18934_, _18933_, _09792_);
  and (_18935_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  and (_18936_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  or (_18937_, _18936_, _18935_);
  and (_18938_, _18937_, _05549_);
  or (_18939_, _18938_, _18934_);
  or (_18940_, _18939_, _05535_);
  and (_18941_, _18940_, _09805_);
  and (_18942_, _18941_, _18930_);
  or (_18943_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  or (_18944_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  and (_18945_, _18944_, _05549_);
  and (_18946_, _18945_, _18943_);
  or (_18947_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  or (_18948_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  and (_18949_, _18948_, _09792_);
  and (_18951_, _18949_, _18947_);
  or (_18952_, _18951_, _18946_);
  or (_18953_, _18952_, _09791_);
  or (_18954_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  or (_18955_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  and (_18956_, _18955_, _05549_);
  and (_18957_, _18956_, _18954_);
  or (_18958_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  or (_18959_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  and (_18960_, _18959_, _09792_);
  and (_18961_, _18960_, _18958_);
  or (_18962_, _18961_, _18957_);
  or (_18963_, _18962_, _05535_);
  and (_18964_, _18963_, _05542_);
  and (_18965_, _18964_, _18953_);
  or (_18966_, _18965_, _18942_);
  and (_18967_, _18966_, _09850_);
  or (_18968_, _18967_, _18920_);
  and (_18969_, _18968_, _09790_);
  and (_18970_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  and (_18971_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or (_18972_, _18971_, _18970_);
  and (_18973_, _18972_, _09792_);
  and (_18974_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  and (_18975_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  or (_18976_, _18975_, _18974_);
  and (_18977_, _18976_, _05549_);
  or (_18978_, _18977_, _18973_);
  and (_18979_, _18978_, _05535_);
  and (_18980_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  and (_18981_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  or (_18982_, _18981_, _18980_);
  and (_18983_, _18982_, _09792_);
  and (_18984_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  and (_18985_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  or (_18986_, _18985_, _18984_);
  and (_18987_, _18986_, _05549_);
  or (_18988_, _18987_, _18983_);
  and (_18989_, _18988_, _09791_);
  or (_18990_, _18989_, _18979_);
  and (_18991_, _18990_, _09805_);
  or (_18992_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  or (_18993_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  and (_18994_, _18993_, _05549_);
  and (_18995_, _18994_, _18992_);
  or (_18996_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  or (_18997_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  and (_18998_, _18997_, _09792_);
  and (_18999_, _18998_, _18996_);
  or (_19000_, _18999_, _18995_);
  and (_19001_, _19000_, _05535_);
  or (_19002_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  or (_19003_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  and (_19004_, _19003_, _05549_);
  and (_19005_, _19004_, _19002_);
  or (_19006_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  or (_19007_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  and (_19008_, _19007_, _09792_);
  and (_19009_, _19008_, _19006_);
  or (_19010_, _19009_, _19005_);
  and (_19011_, _19010_, _09791_);
  or (_19012_, _19011_, _19001_);
  and (_19013_, _19012_, _05542_);
  or (_19014_, _19013_, _18991_);
  and (_19015_, _19014_, _09850_);
  and (_19016_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  and (_19017_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  or (_19018_, _19017_, _19016_);
  and (_19019_, _19018_, _09792_);
  and (_19020_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  and (_19021_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  or (_19022_, _19021_, _19020_);
  and (_19023_, _19022_, _05549_);
  or (_19024_, _19023_, _19019_);
  and (_19025_, _19024_, _05535_);
  and (_19026_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  and (_19027_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  or (_19028_, _19027_, _19026_);
  and (_19029_, _19028_, _09792_);
  and (_19030_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  and (_19031_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  or (_19032_, _19031_, _19030_);
  and (_19033_, _19032_, _05549_);
  or (_19034_, _19033_, _19029_);
  and (_19035_, _19034_, _09791_);
  or (_19036_, _19035_, _19025_);
  and (_19037_, _19036_, _09805_);
  or (_19038_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  or (_19039_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  and (_19040_, _19039_, _19038_);
  and (_19041_, _19040_, _09792_);
  or (_19042_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  or (_19043_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  and (_19044_, _19043_, _19042_);
  and (_19045_, _19044_, _05549_);
  or (_19046_, _19045_, _19041_);
  and (_19047_, _19046_, _05535_);
  or (_19048_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  or (_19049_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  and (_19050_, _19049_, _19048_);
  and (_19051_, _19050_, _09792_);
  or (_19052_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  or (_19053_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  and (_19054_, _19053_, _19052_);
  and (_19055_, _19054_, _05549_);
  or (_19056_, _19055_, _19051_);
  and (_19057_, _19056_, _09791_);
  or (_19058_, _19057_, _19047_);
  and (_19059_, _19058_, _05542_);
  or (_19060_, _19059_, _19037_);
  and (_19061_, _19060_, _05518_);
  or (_19062_, _19061_, _19015_);
  and (_19063_, _19062_, _05520_);
  or (_19064_, _19063_, _18969_);
  or (_19065_, _19064_, _05526_);
  and (_19066_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  and (_19067_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  or (_19068_, _19067_, _19066_);
  and (_19069_, _19068_, _09792_);
  and (_19070_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  and (_19071_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  or (_19072_, _19071_, _19070_);
  and (_19073_, _19072_, _05549_);
  or (_19074_, _19073_, _19069_);
  or (_19075_, _19074_, _09791_);
  and (_19076_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  and (_19077_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  or (_19078_, _19077_, _19076_);
  and (_19079_, _19078_, _09792_);
  and (_19080_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  and (_19081_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  or (_19082_, _19081_, _19080_);
  and (_19083_, _19082_, _05549_);
  or (_19084_, _19083_, _19079_);
  or (_19085_, _19084_, _05535_);
  and (_19086_, _19085_, _09805_);
  and (_19087_, _19086_, _19075_);
  or (_19088_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  or (_19089_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  and (_19090_, _19089_, _05549_);
  and (_19091_, _19090_, _19088_);
  or (_19092_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  or (_19093_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  and (_19094_, _19093_, _09792_);
  and (_19095_, _19094_, _19092_);
  or (_19096_, _19095_, _19091_);
  or (_19097_, _19096_, _09791_);
  or (_19098_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  or (_19099_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  and (_19100_, _19099_, _05549_);
  and (_19101_, _19100_, _19098_);
  or (_19102_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  or (_19103_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  and (_19104_, _19103_, _09792_);
  and (_19105_, _19104_, _19102_);
  or (_19106_, _19105_, _19101_);
  or (_19107_, _19106_, _05535_);
  and (_19108_, _19107_, _05542_);
  and (_19109_, _19108_, _19097_);
  or (_19110_, _19109_, _19087_);
  and (_19111_, _19110_, _09850_);
  and (_19112_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  and (_19113_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  or (_19114_, _19113_, _19112_);
  and (_19115_, _19114_, _09792_);
  and (_19116_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  and (_19117_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  or (_19118_, _19117_, _19116_);
  and (_19119_, _19118_, _05549_);
  or (_19120_, _19119_, _19115_);
  or (_19121_, _19120_, _09791_);
  and (_19122_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  and (_19123_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  or (_19124_, _19123_, _19122_);
  and (_19125_, _19124_, _09792_);
  and (_19126_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  and (_19127_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  or (_19128_, _19127_, _19126_);
  and (_19129_, _19128_, _05549_);
  or (_19130_, _19129_, _19125_);
  or (_19131_, _19130_, _05535_);
  and (_19132_, _19131_, _09805_);
  and (_19133_, _19132_, _19121_);
  or (_19134_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  or (_19135_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  and (_19136_, _19135_, _19134_);
  and (_19137_, _19136_, _09792_);
  or (_19138_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  or (_19139_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  and (_19140_, _19139_, _19138_);
  and (_19141_, _19140_, _05549_);
  or (_19142_, _19141_, _19137_);
  or (_19143_, _19142_, _09791_);
  or (_19144_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  or (_19145_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  and (_19146_, _19145_, _19144_);
  and (_19147_, _19146_, _09792_);
  or (_19148_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  or (_19149_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  and (_19150_, _19149_, _19148_);
  and (_19151_, _19150_, _05549_);
  or (_19152_, _19151_, _19147_);
  or (_19153_, _19152_, _05535_);
  and (_19154_, _19153_, _05542_);
  and (_19155_, _19154_, _19143_);
  or (_19156_, _19155_, _19133_);
  and (_19157_, _19156_, _05518_);
  or (_19158_, _19157_, _19111_);
  and (_19159_, _19158_, _09790_);
  or (_19160_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  or (_19161_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  and (_19162_, _19161_, _19160_);
  and (_19163_, _19162_, _09792_);
  or (_19164_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  or (_19165_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  and (_19166_, _19165_, _19164_);
  and (_19167_, _19166_, _05549_);
  or (_19168_, _19167_, _19163_);
  and (_19169_, _19168_, _09791_);
  or (_19170_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  or (_19171_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  and (_19172_, _19171_, _19170_);
  and (_19173_, _19172_, _09792_);
  or (_19174_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  or (_19175_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  and (_19176_, _19175_, _19174_);
  and (_19177_, _19176_, _05549_);
  or (_19178_, _19177_, _19173_);
  and (_19179_, _19178_, _05535_);
  or (_19180_, _19179_, _19169_);
  and (_19181_, _19180_, _05542_);
  and (_19182_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  and (_19183_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  or (_19184_, _19183_, _19182_);
  and (_19185_, _19184_, _09792_);
  and (_19186_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  and (_19187_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  or (_19188_, _19187_, _19186_);
  and (_19189_, _19188_, _05549_);
  or (_19190_, _19189_, _19185_);
  and (_19191_, _19190_, _09791_);
  and (_19192_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  and (_19193_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  or (_19194_, _19193_, _19192_);
  and (_19195_, _19194_, _09792_);
  and (_19196_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  and (_19197_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  or (_19198_, _19197_, _19196_);
  and (_19199_, _19198_, _05549_);
  or (_19200_, _19199_, _19195_);
  and (_19202_, _19200_, _05535_);
  or (_19203_, _19202_, _19191_);
  and (_19204_, _19203_, _09805_);
  or (_19205_, _19204_, _19181_);
  and (_19206_, _19205_, _05518_);
  or (_19207_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  or (_19208_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  and (_19209_, _19208_, _05549_);
  and (_19210_, _19209_, _19207_);
  or (_19211_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or (_19212_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  and (_19213_, _19212_, _09792_);
  and (_19214_, _19213_, _19211_);
  or (_19215_, _19214_, _19210_);
  and (_19216_, _19215_, _09791_);
  or (_19217_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  or (_19218_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  and (_19219_, _19218_, _05549_);
  and (_19220_, _19219_, _19217_);
  or (_19221_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  or (_19222_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  and (_19223_, _19222_, _09792_);
  and (_19224_, _19223_, _19221_);
  or (_19225_, _19224_, _19220_);
  and (_19226_, _19225_, _05535_);
  or (_19227_, _19226_, _19216_);
  and (_19228_, _19227_, _05542_);
  and (_19229_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  and (_19230_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  or (_19231_, _19230_, _19229_);
  and (_19232_, _19231_, _09792_);
  and (_19233_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  and (_19234_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  or (_19235_, _19234_, _19233_);
  and (_19236_, _19235_, _05549_);
  or (_19237_, _19236_, _19232_);
  and (_19238_, _19237_, _09791_);
  and (_19239_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  and (_19240_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  or (_19241_, _19240_, _19239_);
  and (_19242_, _19241_, _09792_);
  and (_19243_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  and (_19244_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  or (_19245_, _19244_, _19243_);
  and (_19246_, _19245_, _05549_);
  or (_19247_, _19246_, _19242_);
  and (_19248_, _19247_, _05535_);
  or (_19249_, _19248_, _19238_);
  and (_19250_, _19249_, _09805_);
  or (_19251_, _19250_, _19228_);
  and (_19252_, _19251_, _09850_);
  or (_19253_, _19252_, _19206_);
  and (_19254_, _19253_, _05520_);
  or (_19255_, _19254_, _19159_);
  or (_19256_, _19255_, _10033_);
  and (_19257_, _19256_, _19065_);
  or (_19258_, _19257_, _04413_);
  and (_19259_, _19258_, _18874_);
  or (_19260_, _19259_, _05563_);
  or (_19261_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_19262_, _19261_, _22731_);
  and (_11068_, _19262_, _19260_);
  and (_19263_, _16670_, _23887_);
  and (_19264_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  or (_11071_, _19264_, _19263_);
  and (_19265_, _03281_, _23887_);
  and (_19266_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  or (_27164_, _19266_, _19265_);
  and (_19267_, _15996_, _23996_);
  and (_19268_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  or (_11074_, _19268_, _19267_);
  and (_19269_, _02065_, _24134_);
  and (_19270_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  or (_11076_, _19270_, _19269_);
  and (_19271_, _24367_, _24089_);
  and (_19272_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  or (_11077_, _19272_, _19271_);
  and (_19273_, _24367_, _23887_);
  and (_19274_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  or (_11081_, _19274_, _19273_);
  and (_19275_, _24952_, _24051_);
  and (_19276_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  or (_11085_, _19276_, _19275_);
  and (_19277_, _24952_, _23583_);
  and (_19278_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  or (_11088_, _19278_, _19277_);
  and (_19279_, _24900_, _23996_);
  and (_19280_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_11091_, _19280_, _19279_);
  and (_19281_, _16670_, _23548_);
  and (_19282_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  or (_27257_, _19282_, _19281_);
  and (_19283_, _24900_, _23887_);
  and (_19284_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  or (_11103_, _19284_, _19283_);
  and (_19285_, _02065_, _24051_);
  and (_19286_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  or (_27084_, _19286_, _19285_);
  and (_19287_, _24832_, _23583_);
  and (_19288_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  or (_11106_, _19288_, _19287_);
  and (_19289_, _24813_, _23583_);
  and (_19290_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  or (_11109_, _19290_, _19289_);
  and (_19291_, _03281_, _23548_);
  and (_19292_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  or (_11111_, _19292_, _19291_);
  and (_19293_, _24735_, _24089_);
  and (_19294_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  or (_11113_, _19294_, _19293_);
  and (_19295_, _24735_, _23548_);
  and (_19296_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  or (_11115_, _19296_, _19295_);
  and (_19297_, _24694_, _24134_);
  and (_19298_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  or (_11117_, _19298_, _19297_);
  and (_19299_, _24694_, _23887_);
  and (_19300_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  or (_11121_, _19300_, _19299_);
  and (_19301_, _24503_, _23996_);
  and (_19302_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_27195_, _19302_, _19301_);
  and (_19303_, _05431_, _24134_);
  and (_19304_, _05434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  or (_27131_, _19304_, _19303_);
  and (_19305_, _16773_, _23548_);
  and (_19306_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  or (_27236_, _19306_, _19305_);
  and (_19307_, _16670_, _24051_);
  and (_19308_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  or (_11124_, _19308_, _19307_);
  and (_19309_, _24490_, _23548_);
  and (_19310_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  or (_11126_, _19310_, _19309_);
  and (_19311_, _24602_, _23996_);
  and (_19312_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  or (_11128_, _19312_, _19311_);
  and (_19313_, _02065_, _24089_);
  and (_19314_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  or (_11133_, _19314_, _19313_);
  and (_19315_, _24602_, _23887_);
  and (_19316_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  or (_11135_, _19316_, _19315_);
  and (_19317_, _16072_, _24089_);
  and (_19318_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  or (_11142_, _19318_, _19317_);
  and (_19319_, _16670_, _24089_);
  and (_19320_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  or (_11144_, _19320_, _19319_);
  and (_19321_, _24525_, _23548_);
  and (_19322_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  or (_11146_, _19322_, _19321_);
  and (_19323_, _24510_, _24134_);
  and (_19324_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  or (_27192_, _19324_, _19323_);
  and (_19325_, _16670_, _23583_);
  and (_19326_, _16672_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  or (_11156_, _19326_, _19325_);
  and (_19327_, _16072_, _23583_);
  and (_19328_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  or (_11162_, _19328_, _19327_);
  and (_19329_, _24503_, _23583_);
  and (_19330_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  or (_11167_, _19330_, _19329_);
  and (_19331_, _17581_, _23887_);
  and (_19332_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  or (_11170_, _19332_, _19331_);
  and (_19333_, _24490_, _23996_);
  and (_19334_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_11172_, _19334_, _19333_);
  and (_19335_, _24155_, _24134_);
  and (_19336_, _24157_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  or (_11173_, _19336_, _19335_);
  and (_19337_, _24952_, _23996_);
  and (_19338_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_11176_, _19338_, _19337_);
  and (_19339_, _24900_, _24089_);
  and (_19340_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  or (_11178_, _19340_, _19339_);
  and (_19341_, _24900_, _24219_);
  and (_19342_, _24903_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  or (_11180_, _19342_, _19341_);
  and (_19343_, _24302_, _24219_);
  and (_19344_, _24304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  or (_27230_, _19344_, _19343_);
  and (_19345_, _24832_, _24051_);
  and (_19346_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  or (_27199_, _19346_, _19345_);
  and (_19347_, _24832_, _24219_);
  and (_19348_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  or (_27197_, _19348_, _19347_);
  and (_19349_, _24813_, _24051_);
  and (_19350_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  or (_11188_, _19350_, _19349_);
  and (_19351_, _24813_, _23548_);
  and (_19352_, _24815_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  or (_11190_, _19352_, _19351_);
  and (_19353_, _24735_, _24134_);
  and (_19354_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  or (_11192_, _19354_, _19353_);
  and (_19355_, _17581_, _24089_);
  and (_19356_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  or (_11197_, _19356_, _19355_);
  and (_19357_, _03281_, _23583_);
  and (_19358_, _03283_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  or (_11199_, _19358_, _19357_);
  and (_19359_, _24490_, _23583_);
  and (_19360_, _24492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  or (_11200_, _19360_, _19359_);
  and (_19361_, _24602_, _24089_);
  and (_19362_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  or (_11202_, _19362_, _19361_);
  and (_19363_, _24602_, _24219_);
  and (_19364_, _24604_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  or (_11204_, _19364_, _19363_);
  and (_19365_, _24525_, _24051_);
  and (_19366_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  or (_27193_, _19366_, _19365_);
  and (_19367_, _24503_, _24219_);
  and (_19368_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  or (_11213_, _19368_, _19367_);
  and (_19369_, _24367_, _24134_);
  and (_19370_, _24369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  or (_11215_, _19370_, _19369_);
  and (_19371_, _16678_, _24051_);
  and (_19372_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  or (_11220_, _19372_, _19371_);
  and (_19373_, _24735_, _23887_);
  and (_19374_, _24737_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  or (_11222_, _19374_, _19373_);
  and (_19375_, _24694_, _23583_);
  and (_19376_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  or (_11224_, _19376_, _19375_);
  and (_19377_, _16773_, _24219_);
  and (_19378_, _16775_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  or (_11228_, _19378_, _19377_);
  and (_19379_, _24525_, _23887_);
  and (_19380_, _24527_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  or (_11232_, _19380_, _19379_);
  and (_19381_, _24503_, _24089_);
  and (_19382_, _24505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  or (_11234_, _19382_, _19381_);
  and (_19383_, _24952_, _24219_);
  and (_19384_, _24954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  or (_11237_, _19384_, _19383_);
  and (_19385_, _24832_, _23548_);
  and (_19386_, _24834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  or (_11240_, _19386_, _19385_);
  and (_19387_, _16678_, _24089_);
  and (_19388_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  or (_11242_, _19388_, _19387_);
  and (_19389_, _16678_, _23583_);
  and (_19390_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  or (_27256_, _19390_, _19389_);
  and (_19391_, _25210_, _23996_);
  and (_19392_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  or (_27156_, _19392_, _19391_);
  and (_19393_, _16072_, _24134_);
  and (_19394_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  or (_11249_, _19394_, _19393_);
  and (_19395_, _24840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_19396_, _24750_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_19397_, _24750_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_19398_, _19397_, _19396_);
  nor (_19399_, _19398_, _24781_);
  or (_19400_, _19399_, _24747_);
  or (_19401_, _19400_, _19395_);
  or (_19402_, _19398_, _24844_);
  and (_19403_, _19402_, _22731_);
  and (_11258_, _19403_, _19401_);
  and (_19404_, _16072_, _24051_);
  and (_19405_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  or (_11262_, _19405_, _19404_);
  or (_19406_, _24913_, _24851_);
  and (_19407_, _19406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_19408_, _19407_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor (_19409_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _24750_);
  not (_19410_, _19409_);
  nor (_19411_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_19412_, _19411_, _24749_);
  and (_19413_, _19412_, _19410_);
  nor (_19414_, _02137_, _02113_);
  nor (_19415_, _19414_, _24749_);
  nor (_19416_, _19415_, _19413_);
  and (_19417_, _19416_, _19408_);
  or (_19418_, _19417_, _04091_);
  and (_19419_, _19418_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_19420_, _24174_, _24187_);
  nor (_19421_, _24540_, _19420_);
  or (_19422_, _19421_, _19419_);
  nand (_19423_, _19421_, _24531_);
  and (_19424_, _19423_, _19422_);
  nand (_19425_, _19424_, _24704_);
  nand (_19426_, _24703_, _23542_);
  and (_19427_, _19426_, _22731_);
  and (_11268_, _19427_, _19425_);
  and (_11283_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _22731_);
  and (_19428_, _02232_, _24089_);
  and (_19429_, _02234_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  or (_11285_, _19429_, _19428_);
  and (_19430_, _02498_, _23548_);
  and (_19431_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  or (_11287_, _19431_, _19430_);
  and (_19432_, _02882_, _23583_);
  and (_19433_, _02884_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_11289_, _19433_, _19432_);
  and (_19434_, _02980_, _24134_);
  and (_19435_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_26972_, _19435_, _19434_);
  and (_19436_, _02980_, _23548_);
  and (_19437_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_26970_, _19437_, _19436_);
  and (_19438_, _03020_, _23583_);
  and (_19439_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_11292_, _19439_, _19438_);
  and (_19440_, _03180_, _24134_);
  and (_19441_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_11294_, _19441_, _19440_);
  and (_19442_, _03217_, _24219_);
  and (_19443_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_11296_, _19443_, _19442_);
  and (_19444_, _03343_, _24134_);
  and (_19445_, _03346_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_11298_, _19445_, _19444_);
  and (_19446_, _04608_, _24051_);
  and (_19447_, _04610_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_11300_, _19447_, _19446_);
  and (_19448_, _16678_, _23996_);
  and (_19449_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_11303_, _19449_, _19448_);
  and (_19450_, _17581_, _23583_);
  and (_19451_, _17583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  or (_11305_, _19451_, _19450_);
  not (_19452_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or (_19453_, _19407_, _19452_);
  nand (_19454_, _19414_, _19413_);
  or (_19455_, _19454_, _19453_);
  and (_19456_, _19455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_19457_, _19456_, _04687_);
  and (_19458_, _24541_, _24174_);
  and (_19459_, _19458_, _25481_);
  or (_19460_, _19459_, _19457_);
  nand (_19461_, _19459_, _23504_);
  and (_19462_, _19461_, _19460_);
  or (_19463_, _19462_, _24703_);
  nand (_19464_, _24703_, _23989_);
  and (_19465_, _19464_, _22731_);
  and (_11310_, _19465_, _19463_);
  and (_19466_, _04950_, _24134_);
  and (_19467_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  or (_27163_, _19467_, _19466_);
  and (_11315_, _26285_, _22731_);
  and (_19468_, _16072_, _24219_);
  and (_19469_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  or (_26953_, _19469_, _19468_);
  nand (_19470_, _22886_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_19471_, _19470_, _24593_);
  or (_19472_, _19471_, _03798_);
  and (_19473_, _19472_, _24699_);
  nand (_19474_, _24699_, _22886_);
  and (_19475_, _19474_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_19476_, _19475_, _24703_);
  or (_19477_, _19476_, _19473_);
  nand (_19478_, _24703_, _24126_);
  and (_19479_, _19478_, _22731_);
  and (_11322_, _19479_, _19477_);
  and (_19480_, _24089_, _23946_);
  and (_19481_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  or (_11326_, _19481_, _19480_);
  and (_19482_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nand (_19483_, _24779_, _24765_);
  and (_19484_, _19483_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_19485_, _24793_, _24809_);
  and (_19486_, _19485_, _19484_);
  or (_19487_, _19486_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor (_19488_, _24803_, _24750_);
  nand (_19489_, _19488_, _24807_);
  nor (_19490_, _24765_, _24747_);
  or (_19491_, _19490_, _24748_);
  and (_19492_, _19491_, _19489_);
  and (_19493_, _19492_, _19487_);
  or (_19494_, _19493_, _19482_);
  and (_11328_, _19494_, _22731_);
  and (_19495_, _04950_, _24051_);
  and (_19496_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  or (_11331_, _19496_, _19495_);
  and (_11332_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _22731_);
  and (_19497_, _24747_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_19498_, _19490_, _24827_);
  and (_19499_, _24804_, _24750_);
  nand (_19500_, _19499_, _24781_);
  and (_19501_, _19500_, _19498_);
  or (_19502_, _19501_, _19497_);
  and (_19503_, _19485_, _19483_);
  or (_19504_, _19503_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_19505_, _19409_, rst);
  and (_19506_, _19505_, _19504_);
  and (_11334_, _19506_, _19502_);
  and (_11336_, _26377_, _22731_);
  nor (_19507_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _17565_);
  not (_19508_, _19413_);
  and (_19509_, _19415_, _19508_);
  not (_19510_, _19509_);
  or (_19511_, _19510_, _19453_);
  and (_19512_, _19511_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_19513_, _19512_, _19507_);
  and (_19514_, _19458_, _24607_);
  or (_19515_, _19514_, _19513_);
  nand (_19516_, _19514_, _23504_);
  and (_19517_, _19516_, _19515_);
  or (_19518_, _19517_, _24703_);
  nand (_19519_, _24703_, _24043_);
  and (_19520_, _19519_, _22731_);
  and (_11347_, _19520_, _19518_);
  and (_19521_, _19458_, _24533_);
  and (_19522_, _19521_, _24531_);
  nand (_19523_, _24627_, _24188_);
  nand (_19524_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_19525_, _19509_, _19408_);
  or (_19526_, _19525_, _19524_);
  or (_19527_, _19526_, _19521_);
  nand (_19528_, _19527_, _19523_);
  or (_19529_, _19528_, _19522_);
  or (_19530_, _24704_, _23577_);
  and (_19531_, _19530_, _22731_);
  and (_11352_, _19531_, _19529_);
  and (_19532_, _25481_, _24544_);
  nand (_19533_, _19532_, _23504_);
  or (_19534_, _19532_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_19535_, _19534_, _24557_);
  and (_19536_, _19535_, _19533_);
  nor (_19537_, _24557_, _23989_);
  or (_19538_, _19537_, _19536_);
  and (_11355_, _19538_, _22731_);
  and (_19539_, _16020_, _23996_);
  and (_19540_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  or (_11357_, _19540_, _19539_);
  and (_26840_[5], _23765_, _22731_);
  nand (_19541_, _24840_, _24749_);
  nand (_19542_, _19396_, _24747_);
  and (_19543_, _19542_, _22731_);
  and (_11366_, _19543_, _19541_);
  and (_19544_, _16678_, _24134_);
  and (_19545_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  or (_11369_, _19545_, _19544_);
  and (_19546_, _24621_, _25481_);
  nand (_19547_, _19546_, _23504_);
  or (_19548_, _19546_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_19549_, _19548_, _24630_);
  and (_19550_, _19549_, _19547_);
  nor (_19551_, _24630_, _23989_);
  or (_19552_, _19551_, _19550_);
  and (_11372_, _19552_, _22731_);
  and (_19553_, _25432_, _24051_);
  and (_19554_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  or (_11375_, _19554_, _19553_);
  and (_19555_, _01832_, _23887_);
  and (_19556_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  or (_11380_, _19556_, _19555_);
  and (_19557_, _25672_, _23887_);
  and (_19558_, _25674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  or (_11383_, _19558_, _19557_);
  and (_19559_, _03324_, _24089_);
  and (_19560_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_27260_, _19560_, _19559_);
  and (_19561_, _04709_, _23887_);
  and (_19562_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_11390_, _19562_, _19561_);
  and (_19563_, _16072_, _23548_);
  and (_19564_, _16074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  or (_26954_, _19564_, _19563_);
  or (_19565_, _22740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand (_19566_, _22740_, _04912_);
  and (_19567_, _19566_, _22731_);
  and (_26863_[15], _19567_, _19565_);
  nor (_11407_, _00780_, rst);
  and (_11408_, _00352_, _22731_);
  and (_11411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _22731_);
  and (_19568_, _17545_, _23996_);
  and (_19569_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or (_11425_, _19569_, _19568_);
  and (_19570_, _04950_, _23996_);
  and (_19571_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  or (_11436_, _19571_, _19570_);
  and (_19572_, _02498_, _23887_);
  and (_19573_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  or (_11439_, _19573_, _19572_);
  and (_19574_, _03020_, _24089_);
  and (_19575_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_11440_, _19575_, _19574_);
  and (_19576_, _02767_, _24134_);
  and (_19577_, _02769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  or (_11442_, _19577_, _19576_);
  and (_19578_, _03217_, _23548_);
  and (_19579_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_27311_, _19579_, _19578_);
  and (_19580_, _04647_, _24089_);
  and (_19581_, _04649_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_11446_, _19581_, _19580_);
  and (_19582_, _01832_, _23583_);
  and (_19583_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  or (_11450_, _19583_, _19582_);
  and (_19584_, _17545_, _24134_);
  and (_19585_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  or (_11452_, _19585_, _19584_);
  and (_19586_, _03020_, _24051_);
  and (_19587_, _03022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_11455_, _19587_, _19586_);
  or (_19588_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_11462_, _19588_, _03411_);
  and (_19589_, _03404_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_11463_, _19589_, _03406_);
  or (_19590_, _03086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_11466_, _19590_, _03423_);
  and (_11475_, _00540_, _22731_);
  and (_11486_, _16453_, _24747_);
  and (_11487_, _00437_, _22731_);
  and (_19591_, _15581_, _24134_);
  and (_19592_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  or (_27210_, _19592_, _19591_);
  and (_19593_, _02045_, _23996_);
  and (_19594_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_27233_, _19594_, _19593_);
  and (_19595_, _24051_, _23946_);
  and (_19596_, _23998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  or (_11496_, _19596_, _19595_);
  and (_11510_, _00708_, _22731_);
  and (_19597_, _16020_, _23583_);
  and (_19598_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  or (_11512_, _19598_, _19597_);
  and (_11514_, _26381_, _22731_);
  and (_11517_, _00621_, _22731_);
  and (_19599_, _05491_, _23583_);
  and (_19600_, _05493_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  or (_11519_, _19600_, _19599_);
  and (_19601_, _15581_, _23996_);
  and (_19602_, _15583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  or (_11526_, _19602_, _19601_);
  and (_19603_, _24442_, _23996_);
  and (_19604_, _24444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  or (_11528_, _19604_, _19603_);
  and (_19606_, _04950_, _24219_);
  and (_19607_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  or (_11539_, _19607_, _19606_);
  and (_19608_, _01810_, _23887_);
  and (_19609_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  or (_11550_, _19609_, _19608_);
  and (_19610_, _04768_, _24051_);
  and (_19611_, _04770_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  or (_11553_, _19611_, _19610_);
  and (_19612_, _01810_, _24089_);
  and (_19613_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  or (_27217_, _19613_, _19612_);
  and (_19614_, _17545_, _24051_);
  and (_19615_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  or (_27255_, _19615_, _19614_);
  and (_19616_, _04709_, _23548_);
  and (_19617_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_11563_, _19617_, _19616_);
  and (_19618_, _04709_, _24051_);
  and (_19619_, _04711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or (_11592_, _19619_, _19618_);
  and (_19620_, _01810_, _23583_);
  and (_19621_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  or (_11594_, _19621_, _19620_);
  and (_19622_, _24889_, _23996_);
  and (_19623_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_11596_, _19623_, _19622_);
  and (_19624_, _17545_, _24089_);
  and (_19625_, _17547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  or (_11601_, _19625_, _19624_);
  and (_19626_, _03667_, _23548_);
  and (_19627_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_11603_, _19627_, _19626_);
  and (_19628_, _04950_, _23548_);
  and (_19629_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  or (_11605_, _19629_, _19628_);
  and (_19630_, _03667_, _24051_);
  and (_19631_, _03669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  or (_11611_, _19631_, _19630_);
  and (_19632_, _24889_, _24134_);
  and (_19633_, _24891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  or (_11614_, _19633_, _19632_);
  and (_19634_, _03313_, _23548_);
  and (_19635_, _03315_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  or (_27176_, _19635_, _19634_);
  and (_19636_, _16034_, _24219_);
  and (_19637_, _16036_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  or (_11627_, _19637_, _19636_);
  and (_19638_, _03324_, _23583_);
  and (_19640_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_27259_, _19640_, _19638_);
  and (_19641_, _03324_, _23548_);
  and (_19642_, _03326_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  or (_11630_, _19642_, _19641_);
  and (_19643_, _03251_, _24219_);
  and (_19644_, _03253_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_11632_, _19644_, _19643_);
  and (_19645_, _03217_, _23996_);
  and (_19646_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_11638_, _19646_, _19645_);
  and (_19647_, _16020_, _24051_);
  and (_19648_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  or (_11641_, _19648_, _19647_);
  and (_19649_, _15996_, _23583_);
  and (_19650_, _15998_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  or (_11654_, _19650_, _19649_);
  and (_19651_, _03217_, _23583_);
  and (_19652_, _03219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_11656_, _19652_, _19651_);
  and (_19653_, _01810_, _24051_);
  and (_19654_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  or (_11658_, _19654_, _19653_);
  and (_19655_, _03180_, _23887_);
  and (_19656_, _03182_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  or (_26917_, _19656_, _19655_);
  and (_19657_, _03048_, _24089_);
  and (_19658_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_11661_, _19658_, _19657_);
  and (_19659_, _03048_, _23548_);
  and (_19660_, _03050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_26932_, _19660_, _19659_);
  and (_19661_, _04950_, _23583_);
  and (_19662_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  or (_11685_, _19662_, _19661_);
  and (_19663_, _02980_, _24089_);
  and (_19664_, _02982_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  or (_11688_, _19664_, _19663_);
  and (_19665_, _02498_, _24051_);
  and (_19666_, _02500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_11691_, _19666_, _19665_);
  and (_19667_, _16678_, _23548_);
  and (_19668_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  or (_11694_, _19668_, _19667_);
  and (_19669_, _02093_, _23887_);
  and (_19670_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  or (_11696_, _19670_, _19669_);
  and (_19671_, _01832_, _23548_);
  and (_19672_, _01834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  or (_11699_, _19672_, _19671_);
  nor (_19673_, _23531_, _26401_);
  and (_19674_, _23531_, _26401_);
  or (_19675_, _19674_, _19673_);
  and (_11708_, _19675_, _22731_);
  and (_19676_, _04950_, _23887_);
  and (_19677_, _04952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  or (_11711_, _19677_, _19676_);
  and (_19678_, _02093_, _24134_);
  and (_19679_, _02095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  or (_27038_, _19679_, _19678_);
  and (_19680_, _26020_, _24219_);
  and (_19681_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  or (_11714_, _19681_, _19680_);
  and (_11716_, _01167_, _22731_);
  and (_11721_, _26457_, _22731_);
  and (_11723_, _00449_, _22731_);
  and (_11726_, _01042_, _22731_);
  and (_11728_, _01253_, _22731_);
  and (_11730_, _00364_, _22731_);
  and (_11734_, _01325_, _22731_);
  and (_11736_, _26560_, _22731_);
  and (_11738_, _01099_, _22731_);
  and (_11740_, _03830_, _22731_);
  and (_11742_, _00627_, _22731_);
  and (_11746_, _00530_, _22731_);
  and (_19682_, _26020_, _23996_);
  and (_19683_, _26022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  or (_11750_, _19683_, _19682_);
  and (_19684_, _16678_, _24219_);
  and (_19685_, _16680_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  or (_11752_, _19685_, _19684_);
  and (_19686_, _25627_, _24134_);
  and (_19687_, _25629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  or (_11754_, _19687_, _19686_);
  and (_19688_, _25432_, _24089_);
  and (_19689_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  or (_11757_, _19689_, _19688_);
  and (_19690_, _25432_, _23548_);
  and (_19691_, _25434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  or (_11759_, _19691_, _19690_);
  and (_19692_, _25314_, _23583_);
  and (_19693_, _25316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  or (_11761_, _19693_, _19692_);
  and (_19694_, _25210_, _24219_);
  and (_19695_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  or (_27154_, _19695_, _19694_);
  and (_11776_, _00715_, _22731_);
  and (_19696_, _25210_, _24089_);
  and (_19697_, _25212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  or (_11778_, _19697_, _19696_);
  and (_19698_, _24478_, _24089_);
  and (_19699_, _24480_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  or (_11792_, _19699_, _19698_);
  and (_19700_, _16020_, _24219_);
  and (_19701_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  or (_11795_, _19701_, _19700_);
  and (_19702_, _01810_, _24134_);
  and (_19703_, _01812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  or (_11902_, _19703_, _19702_);
  and (_19704_, _03287_, _23583_);
  and (_19705_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  or (_11906_, _19705_, _19704_);
  and (_19706_, _16020_, _23548_);
  and (_19707_, _16022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  or (_11909_, _19707_, _19706_);
  and (_19708_, _03309_, _23583_);
  and (_19709_, _03311_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  or (_11914_, _19709_, _19708_);
  and (_19710_, _11419_, _24219_);
  and (_19711_, _11421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  or (_11916_, _19711_, _19710_);
  and (_19712_, _07779_, _24134_);
  and (_19713_, _07781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  or (_11920_, _19713_, _19712_);
  and (_19714_, _02065_, _23996_);
  and (_19715_, _02067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  or (_11925_, _19715_, _19714_);
  and (_19716_, _08578_, _24219_);
  and (_19717_, _08580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  or (_11927_, _19717_, _19716_);
  and (_19718_, _15605_, _23548_);
  and (_19719_, _15607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  or (_27179_, _19719_, _19718_);
  and (_19720_, _16026_, _24089_);
  and (_19721_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  or (_26949_, _19721_, _19720_);
  and (_19722_, _16026_, _23583_);
  and (_19723_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  or (_11932_, _19723_, _19722_);
  and (_11934_, _01000_, _22731_);
  and (_19724_, _03287_, _24051_);
  and (_19725_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  or (_11937_, _19725_, _19724_);
  and (_19726_, _03287_, _24089_);
  and (_19727_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  or (_12092_, _19727_, _19726_);
  and (_26840_[0], _23681_, _22731_);
  and (_19728_, _16704_, _23548_);
  and (_19729_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  or (_12140_, _19729_, _19728_);
  and (_19730_, _16704_, _23583_);
  and (_19731_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  or (_12142_, _19731_, _19730_);
  and (_19732_, _03043_, _24089_);
  and (_19733_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  or (_12148_, _19733_, _19732_);
  and (_19734_, _16704_, _23887_);
  and (_19735_, _16706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  or (_12154_, _19735_, _19734_);
  nor (_19736_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_19737_, _19736_);
  and (_19738_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_19739_, _19738_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_19740_, _19738_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_19741_, _19740_, _19739_);
  not (_19742_, _19741_);
  and (_19743_, _19739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_19744_, _19739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_19745_, _19744_, _19743_);
  nor (_19746_, _19745_, _05614_);
  and (_19747_, _19745_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_19748_, _19747_, _19746_);
  nor (_19749_, _19748_, _19742_);
  nor (_19750_, _19745_, _05653_);
  and (_19751_, _19745_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_19752_, _19751_, _19750_);
  nor (_19753_, _19752_, _19741_);
  nor (_19754_, _19753_, _19749_);
  nor (_19755_, _19754_, _19737_);
  and (_19756_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _22742_);
  not (_19757_, _19756_);
  and (_19758_, _19745_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_19759_, _19745_, _05641_);
  nor (_19760_, _19759_, _19758_);
  nor (_19761_, _19760_, _19742_);
  nor (_19762_, _19745_, _05634_);
  and (_19763_, _19745_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_19764_, _19763_, _19762_);
  nor (_19765_, _19764_, _19741_);
  nor (_19766_, _19765_, _19761_);
  nor (_19767_, _19766_, _19757_);
  nor (_19768_, _19767_, _19755_);
  not (_19769_, _19738_);
  nor (_19770_, _19745_, _05660_);
  and (_19771_, _19745_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_19772_, _19771_, _19770_);
  nor (_19773_, _19772_, _19742_);
  not (_19774_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_19775_, _19745_, _19774_);
  and (_19776_, _19745_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_19777_, _19776_, _19775_);
  nor (_19778_, _19777_, _19741_);
  nor (_19779_, _19778_, _19773_);
  nor (_19780_, _19779_, _19769_);
  and (_19781_, _22747_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_19782_, _19781_);
  and (_19783_, _19745_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_19784_, _19745_, _06106_);
  nor (_19785_, _19784_, _19783_);
  nor (_19786_, _19785_, _19742_);
  not (_19787_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_19788_, _19745_, _19787_);
  and (_19789_, _19745_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_19790_, _19789_, _19788_);
  nor (_19791_, _19790_, _19741_);
  nor (_19792_, _19791_, _19786_);
  nor (_19793_, _19792_, _19782_);
  nor (_19794_, _19793_, _19780_);
  and (_19795_, _19794_, _19768_);
  and (_19796_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_19797_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor (_19798_, _19797_, _19796_);
  and (_19799_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_19800_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_19801_, _19800_, _19799_);
  and (_19802_, _19801_, _19798_);
  and (_19803_, _19802_, _19742_);
  and (_19804_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_19805_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_19806_, _19805_, _19804_);
  and (_19807_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_19808_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_19809_, _19808_, _19807_);
  and (_19810_, _19809_, _19806_);
  and (_19811_, _19810_, _19741_);
  or (_19812_, _19811_, _19745_);
  nor (_19813_, _19812_, _19803_);
  and (_19814_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_19815_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nor (_19816_, _19815_, _19814_);
  and (_19817_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_19818_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_19819_, _19818_, _19817_);
  and (_19820_, _19819_, _19816_);
  nor (_19821_, _19820_, _19741_);
  and (_19822_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_19823_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_19824_, _19823_, _19822_);
  and (_19825_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_19826_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_19827_, _19826_, _19825_);
  and (_19828_, _19827_, _19824_);
  nor (_19829_, _19828_, _19742_);
  or (_19830_, _19829_, _19821_);
  and (_19831_, _19830_, _19745_);
  nor (_19832_, _19831_, _19813_);
  nor (_19833_, _19832_, _19795_);
  and (_19834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_19835_, _19834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_19836_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_19837_, _19836_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_19838_, _19837_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_19839_, _19838_, _19835_);
  and (_19840_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_19841_, _19840_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_19842_, _19841_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_19843_, _19842_, _19839_);
  and (_19844_, _19843_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_19845_, _19844_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_19846_, _19845_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and (_19847_, _19845_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_19848_, _19847_, _19846_);
  and (_19849_, _19848_, _19833_);
  nor (_19850_, _19844_, _22802_);
  and (_19851_, _19841_, _19839_);
  and (_19852_, _19851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_19853_, _19852_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_19854_, _19853_, _22802_);
  nor (_19855_, _19854_, _19850_);
  not (_19856_, _19855_);
  and (_19857_, _19856_, _19833_);
  nor (_19858_, _19843_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_19859_, _19858_, _19844_);
  and (_19860_, _19859_, _19833_);
  nor (_19861_, _19856_, _19833_);
  nor (_19862_, _19861_, _19857_);
  nor (_19863_, _19851_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_19864_, _19863_, _19852_);
  and (_19865_, _19864_, _19833_);
  and (_19866_, _19840_, _19839_);
  nor (_19867_, _19866_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_19868_, _19867_, _19851_);
  and (_19869_, _19868_, _19833_);
  nor (_19870_, _19864_, _19833_);
  nor (_19871_, _19870_, _19865_);
  nor (_19872_, _19868_, _19833_);
  nor (_19873_, _19872_, _19869_);
  not (_19874_, _19873_);
  and (_19875_, _19839_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_19876_, _19875_, _22784_);
  nor (_19877_, _19875_, _22784_);
  nor (_19878_, _19877_, _19876_);
  not (_19879_, _19878_);
  and (_19880_, _19879_, _19833_);
  nor (_19881_, _19839_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_19882_, _19881_, _19875_);
  and (_19883_, _19882_, _19833_);
  nor (_19884_, _19879_, _19833_);
  nor (_19885_, _19884_, _19880_);
  and (_19886_, _19837_, _19835_);
  nor (_19887_, _19886_, _22776_);
  and (_19888_, _19886_, _22776_);
  nor (_19889_, _19888_, _19887_);
  not (_19890_, _19889_);
  and (_19891_, _19890_, _19833_);
  nor (_19892_, _19890_, _19833_);
  nor (_19893_, _19892_, _19891_);
  not (_19894_, _19893_);
  not (_19895_, _19795_);
  not (_19896_, _19745_);
  and (_19897_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_19898_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_19899_, _19898_, _19897_);
  and (_19900_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_19901_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_19902_, _19901_, _19900_);
  and (_19903_, _19902_, _19899_);
  and (_19904_, _19903_, _19742_);
  and (_19905_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_19906_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_19908_, _19906_, _19905_);
  and (_19909_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_19910_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_19911_, _19910_, _19909_);
  and (_19912_, _19911_, _19908_);
  and (_19913_, _19912_, _19741_);
  nor (_19914_, _19913_, _19904_);
  nor (_19915_, _19914_, _19896_);
  and (_19916_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_19917_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_19918_, _19917_, _19916_);
  and (_19919_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_19920_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_19921_, _19920_, _19919_);
  and (_19922_, _19921_, _19918_);
  and (_19923_, _19922_, _19742_);
  and (_19924_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_19925_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_19926_, _19925_, _19924_);
  and (_19927_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_19928_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_19929_, _19928_, _19927_);
  and (_19930_, _19929_, _19926_);
  and (_19931_, _19930_, _19741_);
  nor (_19932_, _19931_, _19923_);
  nor (_19933_, _19932_, _19745_);
  nor (_19934_, _19933_, _19915_);
  and (_19935_, _19934_, _19895_);
  and (_19936_, _19836_, _19835_);
  nor (_19937_, _19936_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_19938_, _19937_, _19886_);
  and (_19939_, _19938_, _19935_);
  nor (_19940_, _19938_, _19935_);
  nor (_19941_, _19940_, _19939_);
  and (_19942_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_19943_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_19944_, _19943_, _19942_);
  and (_19945_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_19946_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_19947_, _19946_, _19945_);
  and (_19948_, _19947_, _19944_);
  and (_19949_, _19948_, _19741_);
  and (_19950_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_19951_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_19952_, _19951_, _19950_);
  and (_19953_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_19954_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_19955_, _19954_, _19953_);
  and (_19956_, _19955_, _19952_);
  and (_19957_, _19956_, _19742_);
  nor (_19958_, _19957_, _19949_);
  nor (_19959_, _19958_, _19896_);
  and (_19960_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_19961_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_19962_, _19961_, _19960_);
  and (_19963_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_19964_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_19965_, _19964_, _19963_);
  and (_19966_, _19965_, _19962_);
  and (_19967_, _19966_, _19742_);
  and (_19968_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_19969_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_19970_, _19969_, _19968_);
  and (_19971_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_19972_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_19973_, _19972_, _19971_);
  and (_19974_, _19973_, _19970_);
  and (_19975_, _19974_, _19741_);
  nor (_19976_, _19975_, _19967_);
  nor (_19977_, _19976_, _19745_);
  nor (_19978_, _19977_, _19959_);
  and (_19979_, _19978_, _19895_);
  and (_19980_, _19835_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_19981_, _19980_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_19982_, _19981_, _19936_);
  and (_19983_, _19982_, _19979_);
  nor (_19984_, _19982_, _19979_);
  and (_19985_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_19986_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_19987_, _19986_, _19985_);
  and (_19988_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_19989_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_19990_, _19989_, _19988_);
  and (_19991_, _19990_, _19987_);
  and (_19992_, _19991_, _19742_);
  and (_19993_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_19994_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_19995_, _19994_, _19993_);
  and (_19996_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_19997_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_19998_, _19997_, _19996_);
  and (_19999_, _19998_, _19995_);
  and (_20000_, _19999_, _19741_);
  or (_20001_, _20000_, _19745_);
  nor (_20002_, _20001_, _19992_);
  and (_20003_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_20004_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_20005_, _20004_, _20003_);
  and (_20006_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_20007_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_20008_, _20007_, _20006_);
  and (_20009_, _20008_, _20005_);
  nor (_20010_, _20009_, _19741_);
  and (_20011_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_20012_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_20013_, _20012_, _20011_);
  and (_20014_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_20015_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_20016_, _20015_, _20014_);
  and (_20017_, _20016_, _20013_);
  nor (_20018_, _20017_, _19742_);
  or (_20019_, _20018_, _20010_);
  and (_20020_, _20019_, _19745_);
  nor (_20021_, _20020_, _20002_);
  nor (_20022_, _20021_, _19795_);
  nor (_20023_, _19835_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_20024_, _20023_, _19980_);
  and (_20025_, _20024_, _20022_);
  and (_20026_, _19834_, _22758_);
  nor (_20027_, _19834_, _22758_);
  nor (_20028_, _20027_, _20026_);
  not (_20029_, _20028_);
  and (_20030_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_20031_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_20032_, _20031_, _20030_);
  and (_20033_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_20034_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_20035_, _20034_, _20033_);
  and (_20036_, _20035_, _20032_);
  and (_20037_, _20036_, _19742_);
  and (_20038_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_20039_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_20040_, _20039_, _20038_);
  and (_20041_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_20042_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_20043_, _20042_, _20041_);
  and (_20044_, _20043_, _20040_);
  and (_20045_, _20044_, _19741_);
  or (_20046_, _20045_, _19745_);
  nor (_20047_, _20046_, _20037_);
  and (_20048_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_20049_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_20050_, _20049_, _20048_);
  and (_20051_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_20052_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_20053_, _20052_, _20051_);
  and (_20054_, _20053_, _20050_);
  nor (_20055_, _20054_, _19741_);
  and (_20056_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_20057_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_20058_, _20057_, _20056_);
  and (_20059_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_20060_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_20061_, _20060_, _20059_);
  and (_20062_, _20061_, _20058_);
  nor (_20063_, _20062_, _19742_);
  or (_20064_, _20063_, _20055_);
  and (_20065_, _20064_, _19745_);
  nor (_20066_, _20065_, _20047_);
  nor (_20067_, _20066_, _19795_);
  and (_20068_, _20067_, _20029_);
  nor (_20069_, _20067_, _20029_);
  nor (_20070_, _20069_, _20068_);
  not (_20071_, _20070_);
  and (_20072_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_20073_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_20074_, _20073_, _20072_);
  and (_20075_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_20076_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_20077_, _20076_, _20075_);
  and (_20078_, _20077_, _20074_);
  and (_20079_, _20078_, _19742_);
  and (_20080_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_20081_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_20082_, _20081_, _20080_);
  and (_20083_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_20084_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_20085_, _20084_, _20083_);
  and (_20086_, _20085_, _20082_);
  and (_20087_, _20086_, _19741_);
  nor (_20088_, _20087_, _20079_);
  nor (_20089_, _20088_, _19896_);
  and (_20090_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_20091_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_20092_, _20091_, _20090_);
  and (_20093_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_20094_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_20095_, _20094_, _20093_);
  and (_20096_, _20095_, _20092_);
  and (_20097_, _20096_, _19742_);
  and (_20098_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_20099_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_20100_, _20099_, _20098_);
  and (_20101_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_20102_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_20103_, _20102_, _20101_);
  and (_20104_, _20103_, _20100_);
  and (_20105_, _20104_, _19741_);
  nor (_20106_, _20105_, _20097_);
  nor (_20107_, _20106_, _19745_);
  nor (_20108_, _20107_, _20089_);
  and (_20109_, _20108_, _19895_);
  and (_20110_, _22752_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_20111_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _22747_);
  nor (_20112_, _20111_, _20110_);
  not (_20113_, _20112_);
  and (_20114_, _20113_, _20109_);
  and (_20115_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_20116_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_20117_, _20116_, _20115_);
  and (_20118_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_20119_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_20120_, _20119_, _20118_);
  and (_20121_, _20120_, _20117_);
  and (_20122_, _20121_, _19742_);
  and (_20123_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_20124_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_20125_, _20124_, _20123_);
  and (_20126_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_20127_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_20128_, _20127_, _20126_);
  and (_20129_, _20128_, _20125_);
  and (_20130_, _20129_, _19741_);
  or (_20131_, _20130_, _19745_);
  nor (_20132_, _20131_, _20122_);
  and (_20133_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_20134_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_20135_, _20134_, _20133_);
  and (_20136_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_20137_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_20138_, _20137_, _20136_);
  and (_20139_, _20138_, _20135_);
  nor (_20140_, _20139_, _19741_);
  and (_20141_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_20142_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_20143_, _20142_, _20141_);
  and (_20144_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_20145_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_20146_, _20145_, _20144_);
  and (_20147_, _20146_, _20143_);
  nor (_20148_, _20147_, _19742_);
  or (_20149_, _20148_, _20140_);
  and (_20150_, _20149_, _19745_);
  nor (_20151_, _20150_, _20132_);
  nor (_20152_, _20151_, _19795_);
  and (_20153_, _20152_, _22747_);
  and (_20154_, _19781_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_20155_, _19756_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor (_20156_, _20155_, _20154_);
  and (_20157_, _19736_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_20158_, _19738_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_20159_, _20158_, _20157_);
  and (_20160_, _20159_, _20156_);
  and (_20161_, _20160_, _19742_);
  and (_20162_, _19756_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_20163_, _19736_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_20164_, _20163_, _20162_);
  and (_20165_, _19781_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_20166_, _19738_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_20167_, _20166_, _20165_);
  and (_20168_, _20167_, _20164_);
  and (_20169_, _20168_, _19741_);
  or (_20170_, _20169_, _19745_);
  nor (_20171_, _20170_, _20161_);
  and (_20172_, _19756_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_20173_, _19781_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor (_20174_, _20173_, _20172_);
  and (_20175_, _19736_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_20176_, _19738_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_20177_, _20176_, _20175_);
  and (_20178_, _20177_, _20174_);
  nor (_20179_, _20178_, _19741_);
  and (_20180_, _19756_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_20181_, _19738_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_20182_, _20181_, _20180_);
  and (_20183_, _19781_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_20184_, _19736_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_20185_, _20184_, _20183_);
  and (_20186_, _20185_, _20182_);
  nor (_20187_, _20186_, _19742_);
  or (_20188_, _20187_, _20179_);
  and (_20189_, _20188_, _19745_);
  nor (_20190_, _20189_, _20171_);
  nor (_20191_, _20190_, _19795_);
  and (_20192_, _20191_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20193_, _20152_, _22747_);
  nor (_20194_, _20193_, _20153_);
  and (_20195_, _20194_, _20192_);
  nor (_20196_, _20195_, _20153_);
  nor (_20197_, _20113_, _20109_);
  nor (_20198_, _20197_, _20114_);
  not (_20199_, _20198_);
  nor (_20200_, _20199_, _20196_);
  nor (_20201_, _20200_, _20114_);
  nor (_20202_, _20201_, _20071_);
  nor (_20203_, _20202_, _20068_);
  nor (_20204_, _20024_, _20022_);
  nor (_20205_, _20204_, _20025_);
  not (_20206_, _20205_);
  nor (_20207_, _20206_, _20203_);
  nor (_20208_, _20207_, _20025_);
  nor (_20209_, _20208_, _19984_);
  or (_20210_, _20209_, _19983_);
  and (_20211_, _20210_, _19941_);
  nor (_20212_, _20211_, _19939_);
  nor (_20213_, _20212_, _19894_);
  nor (_20214_, _20213_, _19891_);
  nor (_20215_, _19882_, _19833_);
  nor (_20216_, _20215_, _19883_);
  not (_20217_, _20216_);
  nor (_20218_, _20217_, _20214_);
  and (_20219_, _20218_, _19885_);
  or (_20220_, _20219_, _19883_);
  nor (_20221_, _20220_, _19880_);
  nor (_20222_, _20221_, _19874_);
  and (_20223_, _20222_, _19871_);
  or (_20224_, _20223_, _19869_);
  nor (_20225_, _20224_, _19865_);
  nor (_20226_, _19859_, _19833_);
  nor (_20227_, _20226_, _19860_);
  not (_20228_, _20227_);
  nor (_20229_, _20228_, _20225_);
  and (_20230_, _20229_, _19862_);
  or (_20231_, _20230_, _19860_);
  nor (_20232_, _20231_, _19857_);
  nor (_20233_, _19848_, _19833_);
  nor (_20234_, _20233_, _19849_);
  not (_20235_, _20234_);
  nor (_20236_, _20235_, _20232_);
  nor (_20237_, _20236_, _19849_);
  nor (_20238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_20239_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_20240_, _20239_, _20238_);
  not (_20241_, _20240_);
  nor (_20242_, _20241_, _19847_);
  and (_20243_, _20241_, _19847_);
  nor (_20244_, _20243_, _20242_);
  not (_20245_, _20244_);
  and (_20246_, _20245_, _19833_);
  nor (_20247_, _20245_, _19833_);
  nor (_20248_, _20247_, _20246_);
  not (_20249_, _20248_);
  nand (_20250_, _20249_, _20237_);
  or (_20251_, _20249_, _20237_);
  and (_20252_, _20251_, _20250_);
  and (_20253_, _20235_, _20232_);
  nor (_20254_, _20253_, _20236_);
  nand (_20255_, _20254_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_20256_, _20254_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_20257_, _20256_, _20255_);
  nor (_20258_, _20229_, _19860_);
  nor (_20259_, _19855_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_20260_, _19855_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_20261_, _20260_, _20259_);
  nand (_20262_, _20261_, _19833_);
  or (_20263_, _20261_, _19833_);
  and (_20264_, _20263_, _20262_);
  not (_20265_, _20264_);
  nand (_20266_, _20265_, _20258_);
  or (_20267_, _20265_, _20258_);
  and (_20268_, _20267_, _20266_);
  and (_20269_, _20228_, _20225_);
  nor (_20270_, _20269_, _20229_);
  nor (_20271_, _20270_, _22797_);
  and (_20272_, _20270_, _22797_);
  nor (_20273_, _20218_, _19883_);
  and (_20274_, _20273_, _19885_);
  nor (_20275_, _20273_, _19885_);
  nor (_20276_, _20275_, _20274_);
  and (_20277_, _20276_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_20278_, _20276_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_20279_, _20217_, _20214_);
  nor (_20280_, _20279_, _20218_);
  nor (_20281_, _20280_, _22780_);
  and (_20282_, _20280_, _22780_);
  and (_20283_, _20212_, _19894_);
  nor (_20284_, _20283_, _20213_);
  and (_20285_, _20284_, _26136_);
  nor (_20286_, _20284_, _26136_);
  nor (_20287_, _19983_, _19984_);
  nor (_20288_, _20287_, _20208_);
  and (_20289_, _20287_, _20208_);
  or (_20290_, _20289_, _20288_);
  and (_20291_, _20290_, _22767_);
  nor (_20292_, _20290_, _22767_);
  and (_20293_, _20206_, _20203_);
  nor (_20294_, _20293_, _20207_);
  and (_20295_, _20294_, _22762_);
  nor (_20296_, _20294_, _22762_);
  and (_20297_, _20201_, _20071_);
  nor (_20298_, _20297_, _20202_);
  and (_20299_, _20298_, _26149_);
  nor (_20300_, _20298_, _26149_);
  and (_20301_, _20199_, _20196_);
  nor (_20302_, _20301_, _20200_);
  and (_20303_, _20302_, _26153_);
  nor (_20304_, _20302_, _26153_);
  and (_20305_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20306_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_20307_, _20306_, _20305_);
  not (_20308_, _20307_);
  nand (_20309_, _20308_, _20191_);
  or (_20310_, _20308_, _20191_);
  and (_20311_, _20310_, _20309_);
  nor (_20312_, _20194_, _20192_);
  nor (_20313_, _20312_, _20195_);
  and (_20314_, _20313_, _09640_);
  or (_20315_, _20314_, _20311_);
  nor (_20316_, _20313_, _09640_);
  or (_20317_, _20316_, _20315_);
  or (_20318_, _20317_, _20304_);
  or (_20319_, _20318_, _20303_);
  or (_20320_, _20319_, _20300_);
  or (_20321_, _20320_, _20299_);
  or (_20322_, _20321_, _20296_);
  or (_20323_, _20322_, _20295_);
  or (_20324_, _20323_, _20292_);
  or (_20325_, _20324_, _20291_);
  nor (_20326_, _20210_, _19941_);
  nor (_20327_, _20326_, _20211_);
  nor (_20328_, _20327_, _22772_);
  and (_20329_, _20327_, _22772_);
  or (_20330_, _20329_, _20328_);
  or (_20331_, _20330_, _20325_);
  or (_20332_, _20331_, _20286_);
  or (_20333_, _20332_, _20285_);
  or (_20334_, _20333_, _20282_);
  or (_20335_, _20334_, _20281_);
  or (_20336_, _20335_, _20278_);
  or (_20337_, _20336_, _20277_);
  and (_20338_, _20221_, _19874_);
  nor (_20339_, _20338_, _20222_);
  and (_20340_, _20339_, _22789_);
  nor (_20341_, _20339_, _22789_);
  or (_20342_, _20341_, _20340_);
  nor (_20343_, _20222_, _19869_);
  and (_20344_, _19871_, _22793_);
  nor (_20345_, _19871_, _22793_);
  nor (_20346_, _20345_, _20344_);
  nand (_20347_, _20346_, _20343_);
  or (_20348_, _20346_, _20343_);
  and (_20349_, _20348_, _20347_);
  or (_20350_, _20349_, _20342_);
  or (_20351_, _20350_, _20337_);
  or (_20352_, _20351_, _20272_);
  or (_20353_, _20352_, _20271_);
  or (_20354_, _20353_, _20268_);
  or (_20355_, _20354_, _20257_);
  or (_20356_, _20355_, _20252_);
  and (_20357_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_20358_, _20357_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_20359_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_20360_, _20359_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_20361_, _20360_, _20358_);
  not (_20362_, _20361_);
  not (_20363_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_20364_, _20358_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_20365_, _20358_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_20366_, _20365_, _20364_);
  nand (_20367_, _20366_, _20363_);
  or (_20368_, _20366_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_20369_, _20368_, _20367_);
  and (_20370_, _20369_, _20362_);
  not (_20371_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand (_20372_, _20366_, _20371_);
  or (_20373_, _20366_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_20374_, _20373_, _20361_);
  and (_20375_, _20374_, _20372_);
  or (_20376_, _20375_, _20370_);
  or (_20377_, _20376_, _09640_);
  and (_20378_, _26153_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_20379_, \oc8051_symbolic_cxrom1.regvalid [5], _26149_);
  and (_20380_, \oc8051_symbolic_cxrom1.regvalid [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_20381_, _20380_, _20379_);
  and (_20382_, _20381_, _20378_);
  or (_20383_, \oc8051_symbolic_cxrom1.regvalid [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_20384_, \oc8051_symbolic_cxrom1.regvalid [1], _26149_);
  and (_20385_, _20384_, _20357_);
  and (_20386_, _20385_, _20383_);
  or (_20387_, _20386_, _20382_);
  nor (_20388_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_20389_, _20388_, _26153_);
  nor (_20390_, _20389_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_20391_, _20389_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_20392_, _20391_, _20390_);
  and (_20393_, _20392_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_20394_, _20388_, _26153_);
  nor (_20395_, _20394_, _20389_);
  or (_20396_, _05641_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_20397_, _20396_, _20395_);
  or (_20398_, _20397_, _20393_);
  and (_20399_, _20398_, _09640_);
  nor (_20400_, _20392_, _05634_);
  and (_20401_, _20392_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_20402_, _20401_, _20400_);
  or (_20403_, _20402_, _20395_);
  and (_20404_, _20403_, _20399_);
  or (_20405_, _20404_, _20387_);
  and (_20406_, \oc8051_symbolic_cxrom1.regvalid [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_20407_, \oc8051_symbolic_cxrom1.regvalid [6], _26149_);
  or (_20408_, _20407_, _26153_);
  or (_20409_, _20408_, _20406_);
  or (_20410_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_20411_, \oc8051_symbolic_cxrom1.regvalid [10], _26149_);
  and (_20412_, _20411_, _20410_);
  or (_20413_, _20412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_20414_, _20413_, _20409_);
  and (_20415_, _20414_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_20416_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_20417_, \oc8051_symbolic_cxrom1.regvalid [0], _26149_);
  or (_20418_, _20417_, _20416_);
  and (_20419_, _20418_, _26153_);
  and (_20420_, \oc8051_symbolic_cxrom1.regvalid [4], _26149_);
  and (_20421_, \oc8051_symbolic_cxrom1.regvalid [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_20422_, _20421_, _20420_);
  and (_20423_, _20422_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_20424_, _20423_, _20419_);
  and (_20425_, _20424_, _09640_);
  or (_20426_, _20425_, _20415_);
  and (_20427_, _20426_, _09731_);
  and (_20428_, _20378_, _20422_);
  or (_20429_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_20430_, \oc8051_symbolic_cxrom1.regvalid [0], _26149_);
  and (_20431_, _20430_, _20357_);
  and (_20432_, _20431_, _20429_);
  or (_20433_, _20432_, _20428_);
  and (_20434_, _20414_, _09640_);
  or (_20435_, _20434_, _20433_);
  and (_20436_, _20435_, _20427_);
  not (_20437_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nand (_20438_, _20366_, _20437_);
  or (_20439_, _20366_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_20440_, _20439_, _20438_);
  and (_20441_, _20440_, _20362_);
  not (_20442_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nand (_20443_, _20366_, _20442_);
  or (_20444_, _20366_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_20445_, _20444_, _20361_);
  and (_20446_, _20445_, _20443_);
  or (_20447_, _20446_, _20441_);
  or (_20448_, _20447_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_20449_, _20448_, _20436_);
  and (_20450_, _20449_, _20405_);
  and (_20451_, _20450_, _20377_);
  or (_20452_, \oc8051_symbolic_cxrom1.regvalid [10], _09640_);
  or (_20453_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_20454_, _20453_, _20452_);
  nand (_20455_, _20454_, _20392_);
  or (_20456_, \oc8051_symbolic_cxrom1.regvalid [2], _09640_);
  or (_20457_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_20458_, _20457_, _20456_);
  or (_20459_, _20458_, _20392_);
  and (_20460_, _20459_, _20455_);
  or (_20461_, _20460_, _20395_);
  nor (_20462_, _20366_, _19774_);
  and (_20463_, _20366_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_20464_, _20463_, _20462_);
  and (_20465_, _20464_, _20362_);
  or (_20466_, _20366_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_20467_, \oc8051_symbolic_cxrom1.regvalid [12], _26149_);
  and (_20468_, _20467_, _20361_);
  and (_20469_, _20468_, _20466_);
  or (_20470_, _20469_, _09640_);
  or (_20471_, _20470_, _20465_);
  nand (_20472_, \oc8051_symbolic_cxrom1.regvalid [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_20473_, _20472_, _20396_);
  or (_20474_, _20473_, _26153_);
  or (_20475_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_20476_, \oc8051_symbolic_cxrom1.regvalid [11], _26149_);
  and (_20477_, _20476_, _20475_);
  or (_20478_, _20477_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_20479_, _20478_, _20474_);
  and (_20480_, _20479_, _20359_);
  and (_20481_, _09640_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_20482_, _20381_, _26153_);
  or (_20483_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_20484_, \oc8051_symbolic_cxrom1.regvalid [9], _26149_);
  and (_20485_, _20484_, _20483_);
  or (_20486_, _20485_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_20487_, _20486_, _20482_);
  and (_20488_, _20487_, _20481_);
  or (_20489_, _20488_, _20480_);
  and (_20490_, _20479_, _09640_);
  or (_20491_, _20490_, _20387_);
  and (_20492_, _20491_, _20489_);
  and (_20493_, _20492_, _20471_);
  and (_20494_, _20493_, _20461_);
  or (_20495_, _20366_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_20496_, \oc8051_symbolic_cxrom1.regvalid [14], _26149_);
  and (_20497_, _20496_, _20495_);
  or (_20498_, _20497_, _20362_);
  not (_20499_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand (_20500_, _20366_, _20499_);
  or (_20501_, _20366_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_20502_, _20501_, _20500_);
  or (_20503_, _20502_, _20361_);
  and (_20504_, _20503_, _20498_);
  or (_20505_, _20504_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_20506_, _20392_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_20507_, _20407_, _09640_);
  or (_20508_, _20507_, _20506_);
  and (_20509_, _20392_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_20510_, _20420_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_20511_, _20510_, _20509_);
  nand (_20512_, _20511_, _20508_);
  nand (_20513_, _20512_, _20395_);
  and (_20514_, _20513_, _20505_);
  and (_20515_, _20514_, _20494_);
  or (_20516_, _20515_, _20451_);
  nor (_20517_, _19736_, _22752_);
  and (_20518_, _20517_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20519_, _20517_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20520_, _20519_, _20518_);
  nand (_20521_, _20520_, _20371_);
  and (_20522_, _19736_, _22752_);
  nor (_20523_, _20522_, _20517_);
  nor (_20524_, \oc8051_symbolic_cxrom1.regvalid [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_20525_, _20524_);
  and (_20526_, _20525_, _20523_);
  and (_20527_, _20526_, _20521_);
  nor (_20528_, \oc8051_symbolic_cxrom1.regvalid [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_20529_, _20363_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20530_, _20529_, _20528_);
  and (_20531_, _20530_, _22752_);
  or (_20532_, _20531_, _20527_);
  and (_20533_, _20532_, _19736_);
  nand (_20534_, _20520_, _05677_);
  nor (_20535_, \oc8051_symbolic_cxrom1.regvalid [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_20536_, _20535_);
  and (_20537_, _20536_, _19738_);
  and (_20538_, _20537_, _20534_);
  nand (_20539_, _20520_, _20442_);
  nor (_20540_, \oc8051_symbolic_cxrom1.regvalid [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20541_, _20540_, _19757_);
  and (_20542_, _20541_, _20539_);
  or (_20543_, _20542_, _20538_);
  and (_20544_, _20543_, _20523_);
  or (_20545_, _20544_, _20533_);
  not (_20546_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nand (_20547_, _20520_, _20546_);
  not (_20548_, _20523_);
  nor (_20549_, \oc8051_symbolic_cxrom1.regvalid [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20550_, _20549_, _20548_);
  and (_20551_, _20550_, _20547_);
  and (_20552_, _20520_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_20553_, _20520_, _19774_);
  or (_20554_, _20553_, _20552_);
  and (_20555_, _20554_, _20548_);
  or (_20556_, _20555_, _20551_);
  and (_20557_, _20556_, _19781_);
  and (_20558_, _20520_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_20559_, _20520_, _19787_);
  or (_20560_, _20559_, _20558_);
  and (_20561_, _20560_, _19738_);
  and (_20562_, _20520_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_20563_, _20520_, _05653_);
  or (_20564_, _20563_, _20562_);
  and (_20565_, _20564_, _19756_);
  or (_20566_, _20565_, _20561_);
  and (_20567_, _20566_, _20548_);
  or (_20568_, _20567_, _20557_);
  or (_20569_, _20568_, _20545_);
  and (_20570_, _05677_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20571_, _20570_, _22752_);
  and (_20572_, _20571_, _20536_);
  and (_20573_, _20499_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20574_, \oc8051_symbolic_cxrom1.regvalid [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20575_, _20574_, _20573_);
  and (_20576_, _20575_, _22752_);
  nor (_20577_, _20576_, _20572_);
  nor (_20578_, _20577_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_20579_, _20546_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20580_, _20579_, _20549_);
  and (_20581_, _20580_, _20110_);
  and (_20582_, _19774_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20583_, \oc8051_symbolic_cxrom1.regvalid [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_20584_, _20583_, _22752_);
  nor (_20585_, _20584_, _20582_);
  and (_20586_, _20585_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_20587_, _20586_, _20581_);
  not (_20588_, _20587_);
  nor (_20589_, _20588_, _20578_);
  nor (_20590_, _20589_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_20591_, _20590_);
  and (_20592_, _20371_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20593_, _20592_, _22752_);
  and (_20594_, _20593_, _20525_);
  nor (_20595_, _20594_, _20531_);
  nor (_20596_, _20595_, _19782_);
  not (_20597_, _19739_);
  and (_20598_, \oc8051_symbolic_cxrom1.regvalid [9], _22758_);
  and (_20599_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20600_, _20599_, _20598_);
  nor (_20601_, _20600_, _20597_);
  and (_20602_, _19738_, _22752_);
  and (_20603_, _20442_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20604_, _20603_, _20540_);
  and (_20605_, _20604_, _20602_);
  nor (_20606_, _20605_, _20601_);
  not (_20607_, _20606_);
  nor (_20608_, _20607_, _20596_);
  and (_20609_, _20608_, _20591_);
  and (_20610_, _20604_, _20111_);
  nor (_20611_, _20610_, _22742_);
  nor (_20612_, _20595_, _22747_);
  nor (_20613_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_20614_, \oc8051_symbolic_cxrom1.regvalid [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_20615_, _20437_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20616_, _20615_, _20614_);
  and (_20617_, _20616_, _20613_);
  nor (_20618_, _20617_, _20612_);
  and (_20619_, _20618_, _20611_);
  nor (_20620_, _20577_, _22747_);
  nor (_20621_, \oc8051_symbolic_cxrom1.regvalid [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20622_, \oc8051_symbolic_cxrom1.regvalid [8], _22758_);
  nor (_20623_, _20622_, _20621_);
  and (_20624_, _20623_, _20613_);
  and (_20625_, _20580_, _20111_);
  or (_20626_, _20625_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_20627_, _20626_, _20624_);
  nor (_20628_, _20627_, _20620_);
  nor (_20629_, _20628_, _20619_);
  not (_20630_, _22740_);
  nor (_20631_, _20630_, first_instr);
  nand (_20632_, _20631_, _20629_);
  or (_20633_, _20632_, _20609_);
  nor (_20634_, _20633_, _19795_);
  and (_20635_, _20634_, _20569_);
  and (_20636_, _20635_, _20516_);
  nor (_20637_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20638_, _07573_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20639_, _20638_, _20637_);
  and (_20640_, _20639_, _20613_);
  or (_20641_, _20640_, _22758_);
  nor (_20642_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20643_, _08484_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20644_, _20643_, _20642_);
  and (_20645_, _20644_, _19834_);
  nor (_20646_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20647_, _08117_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20648_, _20647_, _20646_);
  and (_20649_, _20648_, _20111_);
  nor (_20650_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20651_, _07816_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20652_, _20651_, _20650_);
  and (_20653_, _20652_, _20110_);
  or (_20654_, _20653_, _20649_);
  or (_20655_, _20654_, _20645_);
  or (_20656_, _20655_, _20641_);
  nor (_20657_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20658_, _07046_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20659_, _20658_, _20657_);
  and (_20660_, _20659_, _20111_);
  nor (_20661_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20662_, _07310_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20663_, _20662_, _20661_);
  and (_20664_, _20663_, _19834_);
  or (_20665_, _20664_, _20660_);
  nor (_20666_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20667_, _06545_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20668_, _20667_, _20666_);
  and (_20669_, _20668_, _20613_);
  nor (_20670_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20671_, _06790_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20672_, _20671_, _20670_);
  and (_20673_, _20672_, _20110_);
  or (_20674_, _20673_, _20669_);
  or (_20675_, _20674_, _20665_);
  or (_20676_, _20675_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_20677_, _20676_, _20656_);
  and (_20678_, _20677_, _20629_);
  nor (_20679_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20680_, _07294_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20681_, _20680_, _20679_);
  and (_20682_, _20681_, _19834_);
  nor (_20683_, _20682_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20684_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20685_, _06518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20686_, _20685_, _20684_);
  and (_20687_, _20686_, _20613_);
  not (_20688_, _20687_);
  nor (_20689_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20690_, _06775_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20691_, _20690_, _20689_);
  and (_20692_, _20691_, _20110_);
  nor (_20693_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20694_, _07023_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20695_, _20694_, _20693_);
  and (_20696_, _20695_, _20111_);
  nor (_20697_, _20696_, _20692_);
  and (_20698_, _20697_, _20688_);
  and (_20699_, _20698_, _20683_);
  nor (_20700_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20701_, _08472_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20702_, _20701_, _20700_);
  and (_20703_, _20702_, _19834_);
  nor (_20704_, _20703_, _22758_);
  nor (_20705_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20706_, _07795_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20707_, _20706_, _20705_);
  and (_20708_, _20707_, _20110_);
  not (_20709_, _20708_);
  nor (_20710_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20711_, _08104_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20712_, _20711_, _20710_);
  and (_20713_, _20712_, _20111_);
  nor (_20714_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20715_, _07556_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20716_, _20715_, _20714_);
  and (_20717_, _20716_, _20613_);
  nor (_20718_, _20717_, _20713_);
  and (_20719_, _20718_, _20709_);
  and (_20720_, _20719_, _20704_);
  nor (_20721_, _20720_, _20699_);
  and (_20722_, _20721_, _20629_);
  nor (_20723_, _20722_, _20678_);
  nor (_20724_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20725_, _08179_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20726_, _20725_, _20724_);
  and (_20727_, _20726_, _20111_);
  nor (_20728_, _20727_, _22758_);
  nor (_20729_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20730_, _07631_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20731_, _20730_, _20729_);
  and (_20732_, _20731_, _20613_);
  nor (_20733_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20734_, _07869_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20735_, _20734_, _20733_);
  and (_20736_, _20735_, _20110_);
  nor (_20737_, _20736_, _20732_);
  nor (_20738_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20739_, _08547_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20740_, _20739_, _20738_);
  and (_20741_, _20740_, _19834_);
  not (_20742_, _20741_);
  and (_20743_, _20742_, _20737_);
  and (_20744_, _20743_, _20728_);
  nor (_20745_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20746_, _07112_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20747_, _20746_, _20745_);
  and (_20748_, _20747_, _20111_);
  nor (_20749_, _20748_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20750_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20751_, _06609_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20752_, _20751_, _20750_);
  and (_20753_, _20752_, _20613_);
  nor (_20754_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20755_, _06845_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20756_, _20755_, _20754_);
  and (_20757_, _20756_, _20110_);
  nor (_20758_, _20757_, _20753_);
  nor (_20759_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20760_, _07375_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20761_, _20760_, _20759_);
  and (_20762_, _20761_, _19834_);
  not (_20763_, _20762_);
  and (_20764_, _20763_, _20758_);
  and (_20765_, _20764_, _20749_);
  nor (_20766_, _20765_, _20744_);
  and (_20767_, _20766_, _20629_);
  nor (_20768_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20769_, _08528_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20770_, _20769_, _20768_);
  and (_20771_, _20770_, _19834_);
  nor (_20772_, _20771_, _22758_);
  nor (_20773_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20774_, _07616_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20775_, _20774_, _20773_);
  and (_20776_, _20775_, _20613_);
  not (_20777_, _20776_);
  nor (_20778_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20779_, _07854_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20780_, _20779_, _20778_);
  and (_20781_, _20780_, _20110_);
  nor (_20782_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20783_, _08162_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20784_, _20783_, _20782_);
  and (_20785_, _20784_, _20111_);
  nor (_20786_, _20785_, _20781_);
  and (_20787_, _20786_, _20777_);
  and (_20788_, _20787_, _20772_);
  nor (_20789_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20790_, _07357_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20791_, _20790_, _20789_);
  and (_20792_, _20791_, _19834_);
  nor (_20793_, _20792_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20794_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20795_, _06594_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20796_, _20795_, _20794_);
  and (_20797_, _20796_, _20613_);
  not (_20798_, _20797_);
  nor (_20799_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20800_, _06832_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20801_, _20800_, _20799_);
  and (_20802_, _20801_, _20110_);
  nor (_20803_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20804_, _07096_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20805_, _20804_, _20803_);
  and (_20806_, _20805_, _20111_);
  nor (_20807_, _20806_, _20802_);
  and (_20808_, _20807_, _20798_);
  and (_20809_, _20808_, _20793_);
  nor (_20810_, _20809_, _20788_);
  and (_20811_, _20810_, _20629_);
  nor (_20812_, _20811_, _20767_);
  and (_20813_, _20812_, _20723_);
  nor (_20814_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20815_, _06804_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20816_, _20815_, _20814_);
  and (_20817_, _20816_, _20110_);
  nor (_20818_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20819_, _07063_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20820_, _20819_, _20818_);
  and (_20821_, _20820_, _20111_);
  nor (_20822_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20823_, _06562_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20824_, _20823_, _20822_);
  and (_20825_, _20824_, _20613_);
  nor (_20826_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20827_, _07329_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20828_, _20827_, _20826_);
  and (_20829_, _20828_, _19834_);
  or (_20830_, _20829_, _20825_);
  or (_20831_, _20830_, _20821_);
  or (_20832_, _20831_, _20817_);
  and (_20833_, _20832_, _22758_);
  nor (_20834_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20835_, _07828_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20836_, _20835_, _20834_);
  and (_20837_, _20836_, _20110_);
  nor (_20838_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20839_, _08134_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20840_, _20839_, _20838_);
  and (_20841_, _20840_, _20111_);
  nor (_20842_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20843_, _07590_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20844_, _20843_, _20842_);
  and (_20845_, _20844_, _20613_);
  nor (_20846_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20847_, _08498_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20848_, _20847_, _20846_);
  and (_20849_, _20848_, _19834_);
  or (_20850_, _20849_, _20845_);
  or (_20851_, _20850_, _20841_);
  or (_20852_, _20851_, _20837_);
  and (_20853_, _20852_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_20854_, _20853_, _20833_);
  and (_20855_, _20854_, _20629_);
  nor (_20856_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20857_, _06818_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20858_, _20857_, _20856_);
  and (_20859_, _20858_, _20110_);
  nor (_20860_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20861_, _07078_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20862_, _20861_, _20860_);
  and (_20863_, _20862_, _20111_);
  nor (_20864_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20865_, _06578_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20866_, _20865_, _20864_);
  and (_20867_, _20866_, _20613_);
  nor (_20868_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20869_, _07339_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20870_, _20869_, _20868_);
  and (_20871_, _20870_, _19834_);
  or (_20872_, _20871_, _20867_);
  or (_20873_, _20872_, _20863_);
  or (_20874_, _20873_, _20859_);
  and (_20875_, _20874_, _22758_);
  nor (_20876_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20877_, _07840_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20878_, _20877_, _20876_);
  and (_20879_, _20878_, _20110_);
  nor (_20880_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20881_, _08148_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20882_, _20881_, _20880_);
  and (_20883_, _20882_, _20111_);
  nor (_20884_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20885_, _07602_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20886_, _20885_, _20884_);
  and (_20887_, _20886_, _20613_);
  nor (_20888_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20889_, _08512_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20890_, _20889_, _20888_);
  and (_20891_, _20890_, _19834_);
  or (_20892_, _20891_, _20887_);
  or (_20893_, _20892_, _20883_);
  or (_20894_, _20893_, _20879_);
  and (_20895_, _20894_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_20896_, _20895_, _20875_);
  and (_20897_, _20896_, _20629_);
  nor (_20898_, _20897_, _20855_);
  nor (_20899_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20900_, _06857_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20901_, _20900_, _20899_);
  and (_20902_, _20901_, _20110_);
  nor (_20903_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20904_, _07127_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20905_, _20904_, _20903_);
  and (_20906_, _20905_, _20111_);
  nor (_20907_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20908_, _07384_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20909_, _20908_, _20907_);
  and (_20910_, _20909_, _19834_);
  nor (_20911_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20912_, _06625_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20913_, _20912_, _20911_);
  and (_20914_, _20913_, _20613_);
  or (_20915_, _20914_, _20910_);
  or (_20916_, _20915_, _20906_);
  or (_20917_, _20916_, _20902_);
  and (_20918_, _20917_, _22758_);
  nor (_20919_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20920_, _07887_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20921_, _20920_, _20919_);
  and (_20922_, _20921_, _20110_);
  nor (_20923_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20924_, _08192_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20925_, _20924_, _20923_);
  and (_20926_, _20925_, _20111_);
  nor (_20927_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20928_, _08564_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20929_, _20928_, _20927_);
  and (_20930_, _20929_, _19834_);
  nor (_20931_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20932_, _07647_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20933_, _20932_, _20931_);
  and (_20934_, _20933_, _20613_);
  or (_20935_, _20934_, _20930_);
  or (_20936_, _20935_, _20926_);
  or (_20937_, _20936_, _20922_);
  and (_20938_, _20937_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_20939_, _20938_, _20918_);
  and (_20940_, _20939_, _20629_);
  not (_20941_, _20940_);
  nor (_20942_, \oc8051_symbolic_cxrom1.regarray[12] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20943_, _05704_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20944_, _20943_, _20942_);
  and (_20945_, _20944_, _20111_);
  nor (_20946_, _20945_, _22758_);
  nor (_20947_, \oc8051_symbolic_cxrom1.regarray[8] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20948_, _05709_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20949_, _20948_, _20947_);
  and (_20950_, _20949_, _20613_);
  nor (_20951_, \oc8051_symbolic_cxrom1.regarray[10] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20952_, _05697_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20953_, _20952_, _20951_);
  and (_20954_, _20953_, _20110_);
  nor (_20955_, _20954_, _20950_);
  nor (_20956_, \oc8051_symbolic_cxrom1.regarray[14] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20957_, _05691_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20958_, _20957_, _20956_);
  and (_20959_, _20958_, _19834_);
  not (_20960_, _20959_);
  and (_20961_, _20960_, _20955_);
  and (_20962_, _20961_, _20946_);
  nor (_20963_, \oc8051_symbolic_cxrom1.regarray[4] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20964_, _05732_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20965_, _20964_, _20963_);
  and (_20966_, _20965_, _20111_);
  nor (_20967_, _20966_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20968_, \oc8051_symbolic_cxrom1.regarray[0] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20969_, _05737_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20970_, _20969_, _20968_);
  and (_20971_, _20970_, _20613_);
  nor (_20972_, \oc8051_symbolic_cxrom1.regarray[2] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20973_, _05719_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20974_, _20973_, _20972_);
  and (_20975_, _20974_, _20110_);
  nor (_20976_, _20975_, _20971_);
  nor (_20977_, \oc8051_symbolic_cxrom1.regarray[6] [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_20978_, _05726_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20979_, _20978_, _20977_);
  and (_20980_, _20979_, _19834_);
  not (_20981_, _20980_);
  and (_20982_, _20981_, _20976_);
  and (_20983_, _20982_, _20967_);
  nor (_20984_, _20983_, _20962_);
  and (_20985_, _20984_, _20629_);
  and (_20986_, _20985_, _20941_);
  and (_20987_, _20986_, _20898_);
  and (_20988_, _20987_, _20813_);
  and (_20989_, _20988_, _20636_);
  and (_20990_, _20989_, _20356_);
  and (_20991_, _20695_, _20110_);
  or (_20992_, _20991_, _20029_);
  and (_20993_, _20686_, _19834_);
  and (_20994_, _20691_, _20613_);
  and (_20995_, _20681_, _20111_);
  or (_20996_, _20995_, _20994_);
  or (_20997_, _20996_, _20993_);
  or (_20998_, _20997_, _20992_);
  and (_20999_, _20712_, _20110_);
  or (_21000_, _20999_, _20028_);
  and (_21001_, _20707_, _20613_);
  and (_21002_, _20702_, _20111_);
  and (_21003_, _20716_, _19834_);
  or (_21004_, _21003_, _21002_);
  or (_21005_, _21004_, _21001_);
  or (_21006_, _21005_, _21000_);
  nand (_21007_, _21006_, _20998_);
  nor (_21008_, _21007_, _20609_);
  nor (_21009_, _21008_, _09731_);
  and (_21010_, _21008_, _09731_);
  or (_21011_, _21010_, _21009_);
  not (_21012_, _20609_);
  and (_21013_, _20659_, _20110_);
  and (_21014_, _20663_, _20111_);
  nor (_21015_, _21014_, _21013_);
  and (_21016_, _20668_, _19834_);
  and (_21017_, _20672_, _20613_);
  nor (_21018_, _21017_, _21016_);
  and (_21019_, _21018_, _21015_);
  and (_21020_, _21019_, _20028_);
  and (_21021_, _20644_, _20111_);
  and (_21022_, _20639_, _19834_);
  and (_21023_, _20648_, _20110_);
  or (_21024_, _21023_, _21022_);
  nor (_21025_, _21024_, _21021_);
  and (_21026_, _20652_, _20613_);
  nor (_21027_, _21026_, _20028_);
  and (_21028_, _21027_, _21025_);
  nor (_21029_, _21028_, _21020_);
  and (_21030_, _21029_, _21012_);
  nor (_21031_, _21030_, _09640_);
  and (_21032_, _21030_, _09640_);
  or (_21033_, _21032_, _21031_);
  or (_21034_, _21033_, _21011_);
  and (_21035_, _20878_, _20613_);
  and (_21036_, _20890_, _20111_);
  and (_21037_, _20882_, _20110_);
  and (_21038_, _20886_, _19834_);
  or (_21039_, _21038_, _21037_);
  or (_21040_, _21039_, _21036_);
  or (_21041_, _21040_, _21035_);
  and (_21042_, _21041_, _20029_);
  and (_21043_, _20858_, _20613_);
  and (_21044_, _20870_, _20111_);
  and (_21045_, _20866_, _19834_);
  and (_21046_, _20862_, _20110_);
  or (_21047_, _21046_, _21045_);
  or (_21048_, _21047_, _21044_);
  or (_21049_, _21048_, _21043_);
  and (_21050_, _21049_, _20028_);
  or (_21051_, _21050_, _21042_);
  and (_21052_, _21051_, _21012_);
  nand (_21053_, _21052_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21054_, _21052_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21055_, _21054_, _21053_);
  and (_21056_, _20836_, _20613_);
  and (_21057_, _20848_, _20111_);
  and (_21058_, _20844_, _19834_);
  and (_21059_, _20840_, _20110_);
  or (_21060_, _21059_, _21058_);
  or (_21061_, _21060_, _21057_);
  or (_21062_, _21061_, _21056_);
  and (_21063_, _21062_, _20029_);
  and (_21064_, _20816_, _20613_);
  and (_21065_, _20828_, _20111_);
  and (_21066_, _20824_, _19834_);
  and (_21067_, _20820_, _20110_);
  or (_21068_, _21067_, _21066_);
  or (_21069_, _21068_, _21065_);
  or (_21070_, _21069_, _21064_);
  and (_21071_, _21070_, _20028_);
  or (_21072_, _21071_, _21063_);
  and (_21073_, _21072_, _21012_);
  nor (_21074_, _21073_, _26153_);
  and (_21075_, _21073_, _26153_);
  or (_21076_, _21075_, _21074_);
  or (_21077_, _21076_, _21055_);
  or (_21078_, _21077_, _21034_);
  and (_21079_, _20958_, _20111_);
  and (_21080_, _20944_, _20110_);
  nor (_21081_, _21080_, _21079_);
  and (_21082_, _20949_, _19834_);
  and (_21083_, _20953_, _20613_);
  nor (_21084_, _21083_, _21082_);
  and (_21085_, _21084_, _21081_);
  and (_21086_, _21085_, _20029_);
  and (_21087_, _20979_, _20111_);
  and (_21088_, _20970_, _19834_);
  and (_21089_, _20965_, _20110_);
  or (_21090_, _21089_, _21088_);
  nor (_21091_, _21090_, _21087_);
  and (_21092_, _20974_, _20613_);
  nor (_21093_, _21092_, _20029_);
  and (_21094_, _21093_, _21091_);
  nor (_21095_, _21094_, _21086_);
  and (_21096_, _21095_, _21012_);
  nand (_21097_, _21096_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_21098_, _21096_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_21099_, _21098_, _21097_);
  and (_21100_, _20905_, _20110_);
  and (_21101_, _20909_, _20111_);
  and (_21102_, _20913_, _19834_);
  or (_21103_, _21102_, _21101_);
  or (_21104_, _21103_, _21100_);
  and (_21105_, _20901_, _20613_);
  or (_21106_, _21105_, _20029_);
  or (_21107_, _21106_, _21104_);
  and (_21108_, _20925_, _20110_);
  or (_21109_, _21108_, _20028_);
  and (_21110_, _20933_, _19834_);
  and (_21111_, _20921_, _20613_);
  and (_21112_, _20929_, _20111_);
  or (_21113_, _21112_, _21111_);
  or (_21114_, _21113_, _21110_);
  or (_21115_, _21114_, _21109_);
  nand (_21116_, _21115_, _21107_);
  nor (_21117_, _21116_, _20609_);
  nand (_21118_, _21117_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or (_21119_, _21117_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_21120_, _21119_, _21118_);
  or (_21121_, _21120_, _21099_);
  and (_21122_, _20747_, _20110_);
  or (_21123_, _21122_, _20029_);
  and (_21124_, _20752_, _19834_);
  and (_21125_, _20756_, _20613_);
  and (_21126_, _20761_, _20111_);
  or (_21127_, _21126_, _21125_);
  or (_21128_, _21127_, _21124_);
  or (_21129_, _21128_, _21123_);
  and (_21130_, _20740_, _20111_);
  or (_21131_, _21130_, _20028_);
  and (_21132_, _20735_, _20613_);
  and (_21133_, _20731_, _19834_);
  or (_21134_, _21133_, _21132_);
  and (_21135_, _20726_, _20110_);
  or (_21136_, _21135_, _21134_);
  or (_21137_, _21136_, _21131_);
  nand (_21138_, _21137_, _21129_);
  nor (_21139_, _21138_, _20609_);
  nand (_21140_, _21139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or (_21141_, _21139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_21142_, _21141_, _21140_);
  and (_21143_, _20805_, _20110_);
  or (_21144_, _21143_, _20029_);
  and (_21145_, _20796_, _19834_);
  and (_21146_, _20801_, _20613_);
  and (_21147_, _20791_, _20111_);
  or (_21148_, _21147_, _21146_);
  or (_21149_, _21148_, _21145_);
  or (_21150_, _21149_, _21144_);
  and (_21151_, _20784_, _20110_);
  or (_21152_, _21151_, _20028_);
  and (_21153_, _20775_, _19834_);
  and (_21154_, _20780_, _20613_);
  and (_21155_, _20770_, _20111_);
  or (_21156_, _21155_, _21154_);
  or (_21157_, _21156_, _21153_);
  or (_21158_, _21157_, _21152_);
  nand (_21159_, _21158_, _21150_);
  nor (_21160_, _21159_, _20609_);
  nor (_21161_, _21160_, _22762_);
  and (_21162_, _21160_, _22762_);
  or (_21163_, _21162_, _21161_);
  or (_21164_, _21163_, _21142_);
  or (_21165_, _21164_, _21121_);
  or (_21166_, _21165_, _21078_);
  nor (_21167_, _20152_, _26128_);
  and (_21168_, _20152_, _26128_);
  or (_21169_, _21168_, _21167_);
  and (_21170_, _20191_, _22780_);
  nor (_21171_, _20191_, _22780_);
  or (_21172_, _21171_, _21170_);
  or (_21173_, _21172_, _21169_);
  or (_21174_, _20067_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_21175_, _20067_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_21176_, _21175_, _21174_);
  nor (_21177_, _20109_, _22789_);
  and (_21178_, _20109_, _22789_);
  or (_21179_, _21178_, _21177_);
  or (_21180_, _21179_, _21176_);
  or (_21181_, _21180_, _21173_);
  or (_21182_, _19979_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_21183_, _19979_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_21184_, _21183_, _21182_);
  and (_21185_, _20022_, _22797_);
  nor (_21186_, _20022_, _22797_);
  or (_21187_, _21186_, _21185_);
  or (_21188_, _21187_, _21184_);
  nor (_21189_, _19833_, _04912_);
  and (_21190_, _19833_, _04912_);
  or (_21191_, _21190_, _21189_);
  nor (_21192_, _19935_, _22806_);
  and (_21193_, _19935_, _22806_);
  or (_21194_, _21193_, _21192_);
  or (_21195_, _21194_, _21191_);
  or (_21196_, _21195_, _21188_);
  or (_21197_, _21196_, _21181_);
  or (_21198_, _21197_, _21166_);
  nor (_21199_, _20985_, _20940_);
  not (_21200_, _20767_);
  not (_21201_, _20722_);
  and (_21202_, _20898_, _21201_);
  and (_21203_, _21202_, _20678_);
  and (_21204_, _21203_, _21200_);
  and (_21205_, _21204_, _21199_);
  and (_21206_, _21205_, _20636_);
  and (_21207_, _21206_, _21198_);
  nor (_21208_, _20152_, _09640_);
  and (_21209_, _20152_, _09640_);
  or (_21210_, _21209_, _21208_);
  nor (_21211_, _19935_, _22772_);
  nor (_21212_, _20767_, _22780_);
  and (_21213_, _20767_, _22780_);
  or (_21214_, _21213_, _21212_);
  nor (_21215_, _20940_, _26128_);
  and (_21216_, _20940_, _26128_);
  or (_21217_, _21216_, _21215_);
  or (_21218_, _21217_, _21214_);
  or (_21219_, _19864_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_21220_, _19864_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_21221_, _21220_, _21219_);
  and (_21222_, _20985_, _22789_);
  nor (_21223_, _20985_, _22789_);
  or (_21224_, _21223_, _21222_);
  or (_21225_, _21224_, _21221_);
  or (_21226_, _21225_, _21218_);
  or (_21227_, _21226_, _21211_);
  or (_21228_, _21227_, _21210_);
  and (_21229_, _20022_, _22762_);
  nor (_21230_, _20022_, _22762_);
  or (_21231_, _21230_, _21229_);
  nor (_21232_, _19859_, _22797_);
  and (_21233_, _19859_, _22797_);
  or (_21234_, _21233_, _21232_);
  or (_21235_, _21234_, _20261_);
  and (_21236_, _19848_, _22806_);
  nor (_21237_, _19848_, _22806_);
  or (_21238_, _21237_, _21236_);
  or (_21239_, _21238_, _20245_);
  or (_21240_, _21239_, _21235_);
  or (_21241_, _21240_, _21231_);
  or (_21242_, _21241_, _21228_);
  and (_21243_, _19935_, _22772_);
  and (_21244_, _19833_, _26136_);
  nor (_21245_, _19833_, _26136_);
  or (_21246_, _21245_, _21244_);
  or (_21247_, _21246_, _21243_);
  nor (_21248_, _20067_, _26149_);
  and (_21249_, _20109_, _26153_);
  or (_21250_, _21249_, _21248_);
  and (_21251_, _20067_, _26149_);
  nor (_21252_, _19979_, _22767_);
  or (_21253_, _21252_, _21251_);
  or (_21254_, _21253_, _21250_);
  and (_21255_, _20191_, _09731_);
  nor (_21256_, _20109_, _26153_);
  or (_21257_, _21256_, _21255_);
  nor (_21258_, _20191_, _09731_);
  and (_21259_, _19979_, _22767_);
  or (_21260_, _21259_, _21258_);
  or (_21261_, _21260_, _21257_);
  or (_21262_, _21261_, _21254_);
  or (_21263_, _21262_, _21247_);
  or (_21264_, _21263_, _21242_);
  not (_21265_, _20678_);
  and (_21266_, _20722_, _21265_);
  and (_21267_, _21266_, _20898_);
  and (_21268_, _21267_, _21264_);
  not (_21269_, _20985_);
  and (_21270_, _20855_, _20678_);
  and (_21271_, _21270_, _20811_);
  and (_21272_, _21271_, _20767_);
  not (_21273_, _20896_);
  and (_21274_, _21273_, _20855_);
  and (_21275_, _21274_, _20723_);
  and (_21276_, _20811_, _20766_);
  and (_21277_, _21276_, _20896_);
  or (_21278_, _21277_, _21275_);
  or (_21279_, _21278_, _21203_);
  or (_21280_, _21279_, _21272_);
  and (_21281_, _21280_, _20940_);
  and (_21282_, _21274_, _21265_);
  and (_21283_, _20941_, _20767_);
  and (_21284_, _21283_, _21282_);
  and (_21285_, _21282_, _20722_);
  and (_21286_, _21285_, _21200_);
  or (_21287_, _21286_, _21284_);
  or (_21288_, _21287_, _21281_);
  and (_21289_, _21288_, _21269_);
  and (_21290_, _20940_, _21200_);
  and (_21291_, _21290_, _21202_);
  or (_21292_, _21291_, _21204_);
  not (_21293_, _20766_);
  and (_21294_, _20811_, _21293_);
  and (_21295_, _21282_, _21294_);
  and (_21296_, _21202_, _20766_);
  not (_21297_, _20810_);
  and (_21298_, _20897_, _21297_);
  not (_21299_, _20811_);
  and (_21300_, _21270_, _21299_);
  or (_21301_, _21300_, _21298_);
  or (_21302_, _21301_, _21296_);
  or (_21303_, _21302_, _21295_);
  and (_21304_, _21303_, _20941_);
  or (_21305_, _21304_, _21292_);
  and (_21306_, _21305_, _20985_);
  and (_21307_, _21285_, _20940_);
  nand (_21308_, _20985_, _20767_);
  nand (_21309_, _21308_, _20810_);
  and (_21310_, _21309_, _21307_);
  or (_21311_, _21310_, _21306_);
  or (_21312_, _21311_, _21289_);
  nor (_21313_, _19868_, _22789_);
  nor (_21314_, _19982_, _22767_);
  and (_21315_, _19982_, _22767_);
  or (_21316_, _21315_, _21314_);
  nor (_21317_, _19889_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_21318_, _19889_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_21319_, _21318_, _21317_);
  or (_21320_, _21319_, _21316_);
  or (_21321_, _21320_, _21313_);
  or (_21322_, _19882_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_21323_, _19882_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_21324_, _21323_, _21322_);
  and (_21325_, _19868_, _22789_);
  or (_21326_, _21325_, _21324_);
  or (_21327_, _21326_, _21321_);
  or (_21328_, _19878_, _26128_);
  nand (_21329_, _19878_, _26128_);
  and (_21330_, _21329_, _21328_);
  nor (_21331_, _19938_, _22772_);
  and (_21332_, _20028_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_21333_, _20028_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_21334_, _21333_, _21332_);
  nor (_21335_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_21336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_21337_, _21336_, _21335_);
  nand (_21338_, _21337_, _20307_);
  nor (_21339_, _20112_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21340_, _20112_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_21341_, _21340_, _21339_);
  or (_21342_, _21341_, _21338_);
  or (_21343_, _21342_, _21334_);
  nor (_21344_, _20024_, _22762_);
  and (_21345_, _20024_, _22762_);
  or (_21346_, _21345_, _21344_);
  or (_21347_, _21346_, _21343_);
  and (_21348_, _19938_, _22772_);
  or (_21349_, _21348_, _21347_);
  or (_21350_, _21349_, _21331_);
  or (_21351_, _21350_, _21221_);
  or (_21352_, _21351_, _21330_);
  or (_21353_, _21352_, _21327_);
  or (_21354_, _21353_, _21240_);
  and (_21355_, _21354_, _21312_);
  and (_21356_, _20898_, _20723_);
  and (_21357_, _21356_, _21294_);
  and (_21358_, _21286_, _21297_);
  or (_21359_, _21358_, _21357_);
  and (_21360_, _21359_, _20986_);
  not (_21361_, _21276_);
  or (_21362_, _21307_, _21361_);
  and (_21363_, _20722_, _20678_);
  and (_21364_, _21363_, _20898_);
  and (_21365_, _21364_, _20940_);
  or (_21366_, _21365_, _21276_);
  and (_21367_, _21366_, _21269_);
  and (_21368_, _21367_, _21362_);
  or (_21369_, _21368_, _21360_);
  and (_21370_, _20518_, _19838_);
  and (_21371_, _21370_, _19842_);
  and (_21372_, _21371_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_21373_, _21372_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_21374_, _21373_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_21375_, _21373_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_21376_, _21375_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_21377_, _21376_, _20240_);
  nor (_21378_, _21377_, _21374_);
  and (_21379_, _21374_, _20241_);
  and (_21380_, _20518_, _19837_);
  nor (_21381_, _21380_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_21382_, _21381_, _21370_);
  and (_21383_, _21382_, _26136_);
  nor (_21384_, _21382_, _26136_);
  or (_21385_, _21384_, _21383_);
  and (_21386_, _20518_, _19836_);
  nor (_21387_, _21386_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_21389_, _21387_, _21380_);
  nor (_21390_, _21389_, _22772_);
  and (_21391_, _21370_, _19840_);
  and (_21392_, _21370_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_21393_, _21392_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_21394_, _21393_, _21391_);
  nor (_21395_, _21394_, _26128_);
  and (_21396_, _21389_, _22772_);
  or (_21397_, _21396_, _21395_);
  or (_21398_, _21397_, _21390_);
  and (_21399_, _20518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_21400_, _20518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_21401_, _21400_, _21399_);
  nand (_21402_, _21401_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_21403_, _21401_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_21404_, _21403_, _21402_);
  nor (_21405_, _21370_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_21406_, _21405_, _21392_);
  and (_21407_, _21406_, _22780_);
  or (_21408_, _21407_, _21404_);
  nor (_21409_, _21399_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_21410_, _21409_, _21386_);
  and (_21411_, _21410_, _22767_);
  nor (_21412_, _21410_, _22767_);
  or (_21413_, _21412_, _21411_);
  or (_21414_, _21413_, _21408_);
  and (_21415_, _21394_, _26128_);
  nor (_21416_, _21406_, _22780_);
  or (_21417_, _20520_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_21418_, _20520_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21419_, _21418_, _21417_);
  nor (_21420_, _19756_, _19781_);
  nor (_21421_, _21420_, _09640_);
  and (_21422_, _21420_, _09640_);
  nor (_21423_, _21422_, _21421_);
  nand (_21424_, _21423_, _20308_);
  nor (_21425_, _20523_, _26153_);
  and (_21426_, _20523_, _26153_);
  or (_21427_, _21426_, _21425_);
  or (_21428_, _21427_, _21424_);
  or (_21429_, _21428_, _21419_);
  or (_21430_, _21429_, _21416_);
  or (_21431_, _21430_, _21415_);
  or (_21432_, _21431_, _21414_);
  or (_21433_, _21432_, _21398_);
  or (_21434_, _21433_, _21385_);
  or (_21435_, _21434_, _21379_);
  nor (_21436_, _21372_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_21437_, _21436_, _21373_);
  nor (_21438_, _21437_, _26114_);
  and (_21439_, _21437_, _26114_);
  or (_21440_, _21439_, _21438_);
  or (_21441_, _21440_, _21435_);
  or (_21442_, _21375_, _21374_);
  and (_21443_, _21442_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_21444_, _21371_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_21445_, _21444_, _21372_);
  nor (_21446_, _21445_, _22797_);
  and (_21447_, _21445_, _22797_);
  and (_21448_, _21370_, _19841_);
  or (_21449_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nand (_21450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_21451_, _21450_, _21449_);
  or (_21452_, _21451_, _21448_);
  nand (_21453_, _21451_, _21448_);
  and (_21454_, _21453_, _21452_);
  nor (_21455_, _21391_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_21456_, _21455_, _21448_);
  nor (_21457_, _21456_, _22789_);
  and (_21458_, _21456_, _22789_);
  or (_21459_, _21458_, _21457_);
  or (_21460_, _21459_, _21454_);
  or (_21461_, _21460_, _21447_);
  or (_21462_, _21461_, _21446_);
  or (_21463_, _21462_, _21443_);
  or (_21464_, _21463_, _21441_);
  or (_21465_, _21464_, _21378_);
  and (_21466_, _21465_, _21369_);
  nor (_21467_, _20897_, _20767_);
  and (_21468_, _21467_, _21271_);
  not (_21469_, _20984_);
  or (_21470_, _21294_, _21469_);
  and (_21471_, _20941_, _20897_);
  and (_21472_, _21471_, _21470_);
  or (_21473_, _21472_, _21468_);
  and (_21474_, _21469_, _20897_);
  not (_21475_, _20721_);
  and (_21476_, _20855_, _21475_);
  and (_21477_, _21476_, _21199_);
  or (_21478_, _21477_, _21474_);
  and (_21479_, _21478_, _21293_);
  and (_21480_, _21298_, _20940_);
  or (_21481_, _20896_, _21475_);
  nand (_21482_, _20984_, _20678_);
  nor (_21483_, _21482_, _21481_);
  or (_21484_, _21483_, _21300_);
  and (_21485_, _21484_, _20940_);
  or (_21486_, _21485_, _21480_);
  or (_21487_, _21486_, _21479_);
  or (_21488_, _21487_, _21473_);
  and (_21489_, _21284_, _21299_);
  or (_21490_, _21274_, _20767_);
  and (_21491_, _21481_, _20940_);
  and (_21492_, _21491_, _21490_);
  or (_21493_, _21492_, _21489_);
  and (_21494_, _21493_, _20985_);
  and (_21495_, _21275_, _20812_);
  or (_21496_, _21495_, _21364_);
  or (_21497_, _21270_, _20813_);
  and (_21498_, _21497_, _21269_);
  or (_21499_, _21498_, _21496_);
  and (_21500_, _21499_, _20941_);
  or (_21501_, _21500_, _21494_);
  or (_21502_, _21501_, _21488_);
  and (_21503_, _19852_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21504_, _21503_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_21505_, _21504_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_21506_, _21505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_21507_, _21505_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_21508_, _21507_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_21509_, _21508_, _20240_);
  nor (_21510_, _21509_, _21506_);
  nand (_21511_, _20240_, _22806_);
  and (_21512_, _21511_, _21506_);
  and (_21513_, _19838_, _19743_);
  and (_21514_, _21513_, _19842_);
  and (_21515_, _21514_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_21516_, _21515_, _22802_);
  and (_21517_, _21515_, _22802_);
  nor (_21518_, _21517_, _21516_);
  and (_21520_, _21518_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_21521_, _21507_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_21522_, _21521_, _21520_);
  or (_21523_, _21522_, _21512_);
  nor (_21524_, _21503_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_21525_, _21524_, _21504_);
  and (_21526_, _21525_, _22797_);
  nor (_21527_, _21525_, _22797_);
  and (_21528_, _21513_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_21529_, _21513_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_21530_, _21529_, _21528_);
  nand (_21531_, _21530_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  or (_21532_, _21530_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_21533_, _21532_, _21531_);
  and (_21534_, _19886_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_21535_, _19836_, _19743_);
  nor (_21536_, _21535_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_21537_, _21536_, _21534_);
  nor (_21538_, _21537_, _22772_);
  and (_21539_, _21537_, _22772_);
  or (_21540_, _21539_, _21538_);
  and (_21541_, _19743_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_21542_, _19743_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_21543_, _21542_, _21541_);
  nand (_21544_, _21543_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_21545_, _21543_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_21546_, _21545_, _21544_);
  or (_21547_, _19745_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_21548_, _19745_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_21549_, _21548_, _21547_);
  or (_21550_, _21549_, _21546_);
  or (_21551_, _21550_, _21540_);
  or (_21552_, _21551_, _21533_);
  and (_21553_, _21513_, _19841_);
  and (_21554_, _21513_, _19840_);
  nor (_21555_, _21554_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_21556_, _21555_, _21553_);
  nor (_21557_, _21556_, _22789_);
  and (_21558_, _21556_, _22789_);
  or (_21559_, _21558_, _21557_);
  or (_21560_, _21559_, _21552_);
  or (_21561_, _21560_, _21527_);
  or (_21562_, _21561_, _21526_);
  nor (_21563_, _21518_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_21564_, _21528_, _22784_);
  and (_21565_, _21528_, _22784_);
  nor (_21566_, _21565_, _21564_);
  nor (_21567_, _21566_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_21568_, _21566_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_21569_, _21534_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_21570_, _21569_, _21513_);
  nor (_21571_, _21570_, _26136_);
  or (_21572_, _19741_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_21573_, _19741_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_21574_, _21573_, _21572_);
  nor (_21575_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_21576_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or (_21577_, _21576_, _21575_);
  and (_21578_, _21577_, _21541_);
  nor (_21579_, _21577_, _21541_);
  or (_21580_, _21579_, _21578_);
  or (_21581_, _21423_, _20307_);
  or (_21582_, _21581_, _21580_);
  or (_21583_, _21582_, _21574_);
  or (_21584_, _21583_, _21571_);
  and (_21585_, _21570_, _26136_);
  or (_21586_, _21553_, _21451_);
  nand (_21587_, _21553_, _21451_);
  and (_21588_, _21587_, _21586_);
  or (_21589_, _21588_, _21585_);
  or (_21590_, _21589_, _21584_);
  or (_21591_, _21590_, _21568_);
  or (_21592_, _21591_, _21567_);
  or (_21593_, _21592_, _21563_);
  or (_21594_, _21593_, _21562_);
  or (_21595_, _21594_, _21523_);
  or (_21596_, _21595_, _21510_);
  and (_21597_, _21596_, _21502_);
  or (_21598_, _21597_, _21466_);
  or (_21599_, _21598_, _21355_);
  or (_21600_, _21599_, _21268_);
  and (_21601_, _21600_, _20636_);
  or (_21602_, _21601_, _21207_);
  or (property_invalid, _21602_, _20990_);
  and (_21603_, _24017_, _23548_);
  and (_21604_, _24053_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  or (_12202_, _21604_, _21603_);
  and (_21605_, _20630_, first_instr);
  or (_00000_, _21605_, rst);
  and (_21606_, _16026_, _24051_);
  and (_21607_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  or (_12224_, _21607_, _21606_);
  and (_21608_, _03033_, _23996_);
  and (_21609_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or (_12251_, _21609_, _21608_);
  and (_21610_, _16008_, _23996_);
  and (_21611_, _16010_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  or (_12261_, _21611_, _21610_);
  and (_21612_, _03033_, _24134_);
  and (_21613_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  or (_12268_, _21613_, _21612_);
  and (_21614_, _05442_, _23583_);
  and (_21615_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  or (_12274_, _21615_, _21614_);
  and (_21616_, _05438_, _23996_);
  and (_21617_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_12280_, _21617_, _21616_);
  and (_21618_, _05438_, _23583_);
  and (_21619_, _05440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  or (_12293_, _21619_, _21618_);
  and (_21621_, _02964_, _24051_);
  and (_21622_, _02966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  or (_27186_, _21622_, _21621_);
  and (_21623_, _03355_, _23996_);
  and (_21624_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_12301_, _21624_, _21623_);
  or (_21625_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_21626_, _21625_, _22731_);
  nand (_21627_, _24189_, _23542_);
  and (_12316_, _21627_, _21626_);
  nand (_21628_, _24210_, _24184_);
  or (_21629_, _24184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_21630_, _21629_, _22731_);
  and (_12325_, _21630_, _21628_);
  and (_21631_, _05442_, _24134_);
  and (_21632_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  or (_12332_, _21632_, _21631_);
  and (_21633_, _03287_, _24219_);
  and (_21634_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  or (_12334_, _21634_, _21633_);
  and (_21635_, _03287_, _23548_);
  and (_21636_, _03289_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  or (_12340_, _21636_, _21635_);
  and (_21637_, _05485_, _23583_);
  and (_21638_, _05487_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  or (_12342_, _21638_, _21637_);
  and (_21639_, _16026_, _23548_);
  and (_21640_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  or (_12344_, _21640_, _21639_);
  and (_21641_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  and (_21643_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  or (_21644_, _21643_, _21641_);
  and (_21645_, _21644_, _09792_);
  and (_21646_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  and (_21647_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  or (_21648_, _21647_, _21646_);
  and (_21649_, _21648_, _05549_);
  or (_21650_, _21649_, _21645_);
  or (_21651_, _21650_, _09791_);
  and (_21652_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  and (_21653_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  or (_21654_, _21653_, _21652_);
  and (_21655_, _21654_, _09792_);
  and (_21656_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  and (_21657_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  or (_21658_, _21657_, _21656_);
  and (_21659_, _21658_, _05549_);
  or (_21660_, _21659_, _21655_);
  or (_21661_, _21660_, _05535_);
  and (_21662_, _21661_, _09805_);
  and (_21663_, _21662_, _21651_);
  or (_21664_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  or (_21665_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  and (_21666_, _21665_, _21664_);
  and (_21667_, _21666_, _09792_);
  or (_21668_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  or (_21669_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  and (_21670_, _21669_, _21668_);
  and (_21671_, _21670_, _05549_);
  or (_21672_, _21671_, _21667_);
  or (_21673_, _21672_, _09791_);
  or (_21674_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  or (_21675_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  and (_21676_, _21675_, _21674_);
  and (_21677_, _21676_, _09792_);
  or (_21678_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  or (_21679_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  and (_21680_, _21679_, _21678_);
  and (_21681_, _21680_, _05549_);
  or (_21682_, _21681_, _21677_);
  or (_21683_, _21682_, _05535_);
  and (_21684_, _21683_, _05542_);
  and (_21685_, _21684_, _21673_);
  or (_21686_, _21685_, _21663_);
  and (_21687_, _21686_, _05518_);
  and (_21688_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  and (_21689_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  or (_21690_, _21689_, _21688_);
  and (_21691_, _21690_, _09792_);
  and (_21692_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  and (_21693_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  or (_21694_, _21693_, _21692_);
  and (_21695_, _21694_, _05549_);
  or (_21696_, _21695_, _21691_);
  or (_21697_, _21696_, _09791_);
  and (_21698_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  and (_21699_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  or (_21700_, _21699_, _21698_);
  and (_21701_, _21700_, _09792_);
  and (_21702_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  and (_21703_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  or (_21704_, _21703_, _21702_);
  and (_21705_, _21704_, _05549_);
  or (_21706_, _21705_, _21701_);
  or (_21707_, _21706_, _05535_);
  and (_21708_, _21707_, _09805_);
  and (_21709_, _21708_, _21697_);
  or (_21710_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  or (_21711_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  and (_21712_, _21711_, _05549_);
  and (_21713_, _21712_, _21710_);
  or (_21714_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  or (_21715_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  and (_21716_, _21715_, _09792_);
  and (_21717_, _21716_, _21714_);
  or (_21718_, _21717_, _21713_);
  or (_21719_, _21718_, _09791_);
  or (_21720_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  or (_21721_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  and (_21722_, _21721_, _05549_);
  and (_21723_, _21722_, _21720_);
  or (_21724_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  or (_21725_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  and (_21726_, _21725_, _09792_);
  and (_21727_, _21726_, _21724_);
  or (_21728_, _21727_, _21723_);
  or (_21729_, _21728_, _05535_);
  and (_21730_, _21729_, _05542_);
  and (_21731_, _21730_, _21719_);
  or (_21732_, _21731_, _21709_);
  and (_21733_, _21732_, _09850_);
  or (_21734_, _21733_, _21687_);
  and (_21735_, _21734_, _09790_);
  and (_21736_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_21737_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_21738_, _21737_, _21736_);
  and (_21739_, _21738_, _09792_);
  and (_21740_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  and (_21741_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  or (_21742_, _21741_, _21740_);
  and (_21743_, _21742_, _05549_);
  or (_21744_, _21743_, _21739_);
  and (_21745_, _21744_, _05535_);
  and (_21746_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_21747_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_21748_, _21747_, _21746_);
  and (_21749_, _21748_, _09792_);
  and (_21750_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_21751_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  or (_21752_, _21751_, _21750_);
  and (_21753_, _21752_, _05549_);
  or (_21754_, _21753_, _21749_);
  and (_21755_, _21754_, _09791_);
  or (_21756_, _21755_, _21745_);
  and (_21757_, _21756_, _09805_);
  or (_21758_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_21759_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_21760_, _21759_, _05549_);
  and (_21761_, _21760_, _21758_);
  or (_21762_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_21763_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_21764_, _21763_, _09792_);
  and (_21765_, _21764_, _21762_);
  or (_21766_, _21765_, _21761_);
  and (_21767_, _21766_, _05535_);
  or (_21768_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  or (_21769_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and (_21770_, _21769_, _05549_);
  and (_21771_, _21770_, _21768_);
  or (_21772_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_21773_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_21774_, _21773_, _09792_);
  and (_21775_, _21774_, _21772_);
  or (_21776_, _21775_, _21771_);
  and (_21777_, _21776_, _09791_);
  or (_21778_, _21777_, _21767_);
  and (_21779_, _21778_, _05542_);
  or (_21780_, _21779_, _21757_);
  and (_21781_, _21780_, _09850_);
  and (_21782_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  and (_21783_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  or (_21784_, _21783_, _21782_);
  and (_21785_, _21784_, _09792_);
  and (_21786_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  and (_21787_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  or (_21788_, _21787_, _21786_);
  and (_21789_, _21788_, _05549_);
  or (_21790_, _21789_, _21785_);
  and (_21791_, _21790_, _05535_);
  and (_21792_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  and (_21793_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  or (_21794_, _21793_, _21792_);
  and (_21795_, _21794_, _09792_);
  and (_21796_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  and (_21797_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  or (_21798_, _21797_, _21796_);
  and (_21799_, _21798_, _05549_);
  or (_21800_, _21799_, _21795_);
  and (_21801_, _21800_, _09791_);
  or (_21802_, _21801_, _21791_);
  and (_21803_, _21802_, _09805_);
  or (_21804_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  or (_21805_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  and (_21806_, _21805_, _21804_);
  and (_21807_, _21806_, _09792_);
  or (_21808_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  or (_21809_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  and (_21810_, _21809_, _21808_);
  and (_21811_, _21810_, _05549_);
  or (_21812_, _21811_, _21807_);
  and (_21813_, _21812_, _05535_);
  or (_21814_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  or (_21815_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  and (_21816_, _21815_, _21814_);
  and (_21817_, _21816_, _09792_);
  or (_21818_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  or (_21819_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  and (_21820_, _21819_, _21818_);
  and (_21821_, _21820_, _05549_);
  or (_21822_, _21821_, _21817_);
  and (_21823_, _21822_, _09791_);
  or (_21824_, _21823_, _21813_);
  and (_21825_, _21824_, _05542_);
  or (_21826_, _21825_, _21803_);
  and (_21827_, _21826_, _05518_);
  or (_21828_, _21827_, _21781_);
  and (_21829_, _21828_, _05520_);
  or (_21830_, _21829_, _21735_);
  or (_21831_, _21830_, _05526_);
  and (_21832_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  and (_21833_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  or (_21834_, _21833_, _21832_);
  and (_21835_, _21834_, _09792_);
  and (_21836_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  and (_21837_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  or (_21838_, _21837_, _21836_);
  and (_21839_, _21838_, _05549_);
  or (_21840_, _21839_, _21835_);
  or (_21841_, _21840_, _09791_);
  and (_21842_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  and (_21843_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  or (_21844_, _21843_, _21842_);
  and (_21845_, _21844_, _09792_);
  and (_21846_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  and (_21847_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  or (_21848_, _21847_, _21846_);
  and (_21849_, _21848_, _05549_);
  or (_21850_, _21849_, _21845_);
  or (_21851_, _21850_, _05535_);
  and (_21852_, _21851_, _09805_);
  and (_21853_, _21852_, _21841_);
  or (_21854_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  or (_21855_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  and (_21856_, _21855_, _05549_);
  and (_21857_, _21856_, _21854_);
  or (_21858_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  or (_21859_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  and (_21860_, _21859_, _09792_);
  and (_21861_, _21860_, _21858_);
  or (_21862_, _21861_, _21857_);
  or (_21863_, _21862_, _09791_);
  or (_21864_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  or (_21865_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  and (_21866_, _21865_, _05549_);
  and (_21867_, _21866_, _21864_);
  or (_21868_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  or (_21869_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  and (_21870_, _21869_, _09792_);
  and (_21871_, _21870_, _21868_);
  or (_21872_, _21871_, _21867_);
  or (_21873_, _21872_, _05535_);
  and (_21874_, _21873_, _05542_);
  and (_21875_, _21874_, _21863_);
  or (_21876_, _21875_, _21853_);
  and (_21877_, _21876_, _09850_);
  and (_21878_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  and (_21879_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  or (_21880_, _21879_, _21878_);
  and (_21881_, _21880_, _09792_);
  and (_21882_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  and (_21883_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  or (_21884_, _21883_, _21882_);
  and (_21885_, _21884_, _05549_);
  or (_21886_, _21885_, _21881_);
  or (_21887_, _21886_, _09791_);
  and (_21888_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  and (_21889_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  or (_21890_, _21889_, _21888_);
  and (_21891_, _21890_, _09792_);
  and (_21892_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  and (_21893_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  or (_21894_, _21893_, _21892_);
  and (_21895_, _21894_, _05549_);
  or (_21896_, _21895_, _21891_);
  or (_21897_, _21896_, _05535_);
  and (_21898_, _21897_, _09805_);
  and (_21899_, _21898_, _21887_);
  or (_21900_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  or (_21901_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  and (_21902_, _21901_, _21900_);
  and (_21903_, _21902_, _09792_);
  or (_21904_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  or (_21905_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  and (_21906_, _21905_, _21904_);
  and (_21907_, _21906_, _05549_);
  or (_21908_, _21907_, _21903_);
  or (_21909_, _21908_, _09791_);
  or (_21910_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  or (_21911_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  and (_21912_, _21911_, _21910_);
  and (_21913_, _21912_, _09792_);
  or (_21914_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  or (_21915_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  and (_21916_, _21915_, _21914_);
  and (_21917_, _21916_, _05549_);
  or (_21918_, _21917_, _21913_);
  or (_21919_, _21918_, _05535_);
  and (_21920_, _21919_, _05542_);
  and (_21921_, _21920_, _21909_);
  or (_21922_, _21921_, _21899_);
  and (_21923_, _21922_, _05518_);
  or (_21924_, _21923_, _21877_);
  and (_21925_, _21924_, _09790_);
  or (_21926_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  or (_21927_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  and (_21928_, _21927_, _21926_);
  and (_21929_, _21928_, _09792_);
  or (_21930_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  or (_21931_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  and (_21932_, _21931_, _21930_);
  and (_21933_, _21932_, _05549_);
  or (_21934_, _21933_, _21929_);
  and (_21935_, _21934_, _09791_);
  or (_21936_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  or (_21937_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  and (_21938_, _21937_, _21936_);
  and (_21939_, _21938_, _09792_);
  or (_21940_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  or (_21941_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  and (_21942_, _21941_, _21940_);
  and (_21943_, _21942_, _05549_);
  or (_21944_, _21943_, _21939_);
  and (_21945_, _21944_, _05535_);
  or (_21946_, _21945_, _21935_);
  and (_21947_, _21946_, _05542_);
  and (_21948_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  and (_21949_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  or (_21950_, _21949_, _21948_);
  and (_21951_, _21950_, _09792_);
  and (_21952_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  and (_21953_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  or (_21954_, _21953_, _21952_);
  and (_21955_, _21954_, _05549_);
  or (_21956_, _21955_, _21951_);
  and (_21957_, _21956_, _09791_);
  and (_21958_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  and (_21959_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  or (_21960_, _21959_, _21958_);
  and (_21961_, _21960_, _09792_);
  and (_21962_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  and (_21963_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  or (_21964_, _21963_, _21962_);
  and (_21965_, _21964_, _05549_);
  or (_21966_, _21965_, _21961_);
  and (_21967_, _21966_, _05535_);
  or (_21968_, _21967_, _21957_);
  and (_21969_, _21968_, _09805_);
  or (_21970_, _21969_, _21947_);
  and (_21971_, _21970_, _05518_);
  or (_21972_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  or (_21973_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  and (_21974_, _21973_, _05549_);
  and (_21975_, _21974_, _21972_);
  or (_21976_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  or (_21977_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  and (_21978_, _21977_, _09792_);
  and (_21979_, _21978_, _21976_);
  or (_21980_, _21979_, _21975_);
  and (_21981_, _21980_, _09791_);
  or (_21982_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  or (_21983_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  and (_21984_, _21983_, _05549_);
  and (_21985_, _21984_, _21982_);
  or (_21986_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  or (_21987_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  and (_21988_, _21987_, _09792_);
  and (_21989_, _21988_, _21986_);
  or (_21990_, _21989_, _21985_);
  and (_21991_, _21990_, _05535_);
  or (_21992_, _21991_, _21981_);
  and (_21993_, _21992_, _05542_);
  and (_21994_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  and (_21995_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  or (_21996_, _21995_, _21994_);
  and (_21997_, _21996_, _09792_);
  and (_21998_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  and (_21999_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  or (_22000_, _21999_, _21998_);
  and (_22001_, _22000_, _05549_);
  or (_22002_, _22001_, _21997_);
  and (_22003_, _22002_, _09791_);
  and (_22004_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  and (_22005_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  or (_22006_, _22005_, _22004_);
  and (_22007_, _22006_, _09792_);
  and (_22008_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  and (_22009_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  or (_22010_, _22009_, _22008_);
  and (_22011_, _22010_, _05549_);
  or (_22012_, _22011_, _22007_);
  and (_22013_, _22012_, _05535_);
  or (_22014_, _22013_, _22003_);
  and (_22015_, _22014_, _09805_);
  or (_22016_, _22015_, _21993_);
  and (_22017_, _22016_, _09850_);
  or (_22018_, _22017_, _21971_);
  and (_22019_, _22018_, _05520_);
  or (_22020_, _22019_, _21925_);
  or (_22021_, _22020_, _10033_);
  and (_22022_, _22021_, _21831_);
  or (_22023_, _22022_, _00143_);
  and (_22024_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  and (_22025_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  or (_22026_, _22025_, _22024_);
  and (_22027_, _22026_, _09792_);
  and (_22028_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  and (_22029_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  or (_22030_, _22029_, _22028_);
  and (_22031_, _22030_, _05549_);
  or (_22032_, _22031_, _22027_);
  or (_22033_, _22032_, _09791_);
  and (_22034_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  and (_22035_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  or (_22036_, _22035_, _22034_);
  and (_22037_, _22036_, _09792_);
  and (_22038_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  and (_22039_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  or (_22040_, _22039_, _22038_);
  and (_22041_, _22040_, _05549_);
  or (_22042_, _22041_, _22037_);
  or (_22043_, _22042_, _05535_);
  and (_22044_, _22043_, _09805_);
  and (_22045_, _22044_, _22033_);
  or (_22046_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  or (_22047_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  and (_22048_, _22047_, _22046_);
  and (_22049_, _22048_, _09792_);
  or (_22050_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  or (_22051_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  and (_22052_, _22051_, _22050_);
  and (_22053_, _22052_, _05549_);
  or (_22054_, _22053_, _22049_);
  or (_22055_, _22054_, _09791_);
  or (_22056_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  or (_22057_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  and (_22058_, _22057_, _22056_);
  and (_22059_, _22058_, _09792_);
  or (_22060_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  or (_22061_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  and (_22062_, _22061_, _22060_);
  and (_22063_, _22062_, _05549_);
  or (_22064_, _22063_, _22059_);
  or (_22065_, _22064_, _05535_);
  and (_22066_, _22065_, _05542_);
  and (_22067_, _22066_, _22055_);
  or (_22068_, _22067_, _22045_);
  and (_22069_, _22068_, _05518_);
  and (_22070_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  and (_22071_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  or (_22072_, _22071_, _22070_);
  and (_22073_, _22072_, _09792_);
  and (_22074_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  and (_22075_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  or (_22076_, _22075_, _22074_);
  and (_22077_, _22076_, _05549_);
  or (_22078_, _22077_, _22073_);
  or (_22079_, _22078_, _09791_);
  and (_22080_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  and (_22081_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  or (_22082_, _22081_, _22080_);
  and (_22083_, _22082_, _09792_);
  and (_22084_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  and (_22085_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  or (_22086_, _22085_, _22084_);
  and (_22087_, _22086_, _05549_);
  or (_22088_, _22087_, _22083_);
  or (_22089_, _22088_, _05535_);
  and (_22090_, _22089_, _09805_);
  and (_22091_, _22090_, _22079_);
  or (_22092_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  or (_22093_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  and (_22094_, _22093_, _05549_);
  and (_22095_, _22094_, _22092_);
  or (_22096_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  or (_22097_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  and (_22098_, _22097_, _09792_);
  and (_22099_, _22098_, _22096_);
  or (_22100_, _22099_, _22095_);
  or (_22101_, _22100_, _09791_);
  or (_22102_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  or (_22103_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  and (_22104_, _22103_, _05549_);
  and (_22105_, _22104_, _22102_);
  or (_22106_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  or (_22107_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  and (_22108_, _22107_, _09792_);
  and (_22109_, _22108_, _22106_);
  or (_22110_, _22109_, _22105_);
  or (_22111_, _22110_, _05535_);
  and (_22112_, _22111_, _05542_);
  and (_22113_, _22112_, _22101_);
  or (_22114_, _22113_, _22091_);
  and (_22115_, _22114_, _09850_);
  or (_22116_, _22115_, _22069_);
  and (_22117_, _22116_, _09790_);
  and (_22118_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  and (_22119_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  or (_22120_, _22119_, _22118_);
  and (_22121_, _22120_, _09792_);
  and (_22122_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  and (_22123_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  or (_22124_, _22123_, _22122_);
  and (_22125_, _22124_, _05549_);
  or (_22126_, _22125_, _22121_);
  and (_22127_, _22126_, _05535_);
  and (_22128_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  and (_22129_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  or (_22130_, _22129_, _22128_);
  and (_22131_, _22130_, _09792_);
  and (_22132_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  and (_22133_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  or (_22134_, _22133_, _22132_);
  and (_22135_, _22134_, _05549_);
  or (_22136_, _22135_, _22131_);
  and (_22137_, _22136_, _09791_);
  or (_22138_, _22137_, _22127_);
  and (_22139_, _22138_, _09805_);
  or (_22140_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  or (_22141_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  and (_22142_, _22141_, _05549_);
  and (_22143_, _22142_, _22140_);
  or (_22144_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  or (_22145_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  and (_22146_, _22145_, _09792_);
  and (_22147_, _22146_, _22144_);
  or (_22148_, _22147_, _22143_);
  and (_22149_, _22148_, _05535_);
  or (_22150_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  or (_22151_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  and (_22152_, _22151_, _05549_);
  and (_22153_, _22152_, _22150_);
  or (_22154_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  or (_22155_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  and (_22156_, _22155_, _09792_);
  and (_22157_, _22156_, _22154_);
  or (_22158_, _22157_, _22153_);
  and (_22159_, _22158_, _09791_);
  or (_22160_, _22159_, _22149_);
  and (_22161_, _22160_, _05542_);
  or (_22162_, _22161_, _22139_);
  and (_22163_, _22162_, _09850_);
  and (_22164_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  and (_22165_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  or (_22166_, _22165_, _22164_);
  and (_22167_, _22166_, _09792_);
  and (_22168_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  and (_22169_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  or (_22170_, _22169_, _22168_);
  and (_22171_, _22170_, _05549_);
  or (_22172_, _22171_, _22167_);
  and (_22173_, _22172_, _05535_);
  and (_22174_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  and (_22175_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  or (_22176_, _22175_, _22174_);
  and (_22177_, _22176_, _09792_);
  and (_22178_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  and (_22179_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  or (_22180_, _22179_, _22178_);
  and (_22181_, _22180_, _05549_);
  or (_22182_, _22181_, _22177_);
  and (_22183_, _22182_, _09791_);
  or (_22184_, _22183_, _22173_);
  and (_22185_, _22184_, _09805_);
  or (_22186_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  or (_22187_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  and (_22188_, _22187_, _22186_);
  and (_22189_, _22188_, _09792_);
  or (_22190_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  or (_22191_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  and (_22192_, _22191_, _22190_);
  and (_22193_, _22192_, _05549_);
  or (_22194_, _22193_, _22189_);
  and (_22195_, _22194_, _05535_);
  or (_22196_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  or (_22197_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  and (_22198_, _22197_, _22196_);
  and (_22199_, _22198_, _09792_);
  or (_22200_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  or (_22201_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  and (_22202_, _22201_, _22200_);
  and (_22203_, _22202_, _05549_);
  or (_22204_, _22203_, _22199_);
  and (_22205_, _22204_, _09791_);
  or (_22206_, _22205_, _22195_);
  and (_22207_, _22206_, _05542_);
  or (_22208_, _22207_, _22185_);
  and (_22209_, _22208_, _05518_);
  or (_22210_, _22209_, _22163_);
  and (_22211_, _22210_, _05520_);
  or (_22212_, _22211_, _22117_);
  or (_22213_, _22212_, _05526_);
  and (_22214_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  and (_22215_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  or (_22216_, _22215_, _22214_);
  and (_22217_, _22216_, _09792_);
  and (_22218_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  and (_22219_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  or (_22220_, _22219_, _22218_);
  and (_22221_, _22220_, _05549_);
  or (_22222_, _22221_, _22217_);
  or (_22223_, _22222_, _09791_);
  and (_22224_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  and (_22225_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  or (_22226_, _22225_, _22224_);
  and (_22227_, _22226_, _09792_);
  and (_22228_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  and (_22229_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  or (_22230_, _22229_, _22228_);
  and (_22231_, _22230_, _05549_);
  or (_22232_, _22231_, _22227_);
  or (_22233_, _22232_, _05535_);
  and (_22234_, _22233_, _09805_);
  and (_22235_, _22234_, _22223_);
  or (_22236_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  or (_22237_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  and (_22238_, _22237_, _05549_);
  and (_22239_, _22238_, _22236_);
  or (_22240_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  or (_22241_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  and (_22242_, _22241_, _09792_);
  and (_22243_, _22242_, _22240_);
  or (_22244_, _22243_, _22239_);
  or (_22245_, _22244_, _09791_);
  or (_22246_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  or (_22247_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  and (_22248_, _22247_, _05549_);
  and (_22249_, _22248_, _22246_);
  or (_22250_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  or (_22251_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  and (_22252_, _22251_, _09792_);
  and (_22253_, _22252_, _22250_);
  or (_22254_, _22253_, _22249_);
  or (_22255_, _22254_, _05535_);
  and (_22256_, _22255_, _05542_);
  and (_22257_, _22256_, _22245_);
  or (_22258_, _22257_, _22235_);
  and (_22259_, _22258_, _09850_);
  and (_22260_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  and (_22261_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  or (_22262_, _22261_, _22260_);
  and (_22263_, _22262_, _09792_);
  and (_22264_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  and (_22265_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  or (_22266_, _22265_, _22264_);
  and (_22267_, _22266_, _05549_);
  or (_22268_, _22267_, _22263_);
  or (_22269_, _22268_, _09791_);
  and (_22270_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  and (_22271_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  or (_22272_, _22271_, _22270_);
  and (_22273_, _22272_, _09792_);
  and (_22274_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  and (_22275_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  or (_22276_, _22275_, _22274_);
  and (_22277_, _22276_, _05549_);
  or (_22278_, _22277_, _22273_);
  or (_22279_, _22278_, _05535_);
  and (_22280_, _22279_, _09805_);
  and (_22281_, _22280_, _22269_);
  or (_22282_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  or (_22283_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  and (_22284_, _22283_, _22282_);
  and (_22285_, _22284_, _09792_);
  or (_22286_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  or (_22287_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  and (_22288_, _22287_, _22286_);
  and (_22289_, _22288_, _05549_);
  or (_22290_, _22289_, _22285_);
  or (_22291_, _22290_, _09791_);
  or (_22292_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  or (_22293_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  and (_22294_, _22293_, _22292_);
  and (_22295_, _22294_, _09792_);
  or (_22296_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  or (_22297_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  and (_22298_, _22297_, _22296_);
  and (_22299_, _22298_, _05549_);
  or (_22300_, _22299_, _22295_);
  or (_22301_, _22300_, _05535_);
  and (_22302_, _22301_, _05542_);
  and (_22303_, _22302_, _22291_);
  or (_22304_, _22303_, _22281_);
  and (_22305_, _22304_, _05518_);
  or (_22306_, _22305_, _22259_);
  and (_22307_, _22306_, _09790_);
  or (_22308_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  or (_22309_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  and (_22310_, _22309_, _22308_);
  and (_22311_, _22310_, _09792_);
  or (_22312_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  or (_22313_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  and (_22314_, _22313_, _22312_);
  and (_22315_, _22314_, _05549_);
  or (_22316_, _22315_, _22311_);
  and (_22317_, _22316_, _09791_);
  or (_22318_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  or (_22319_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  and (_22320_, _22319_, _22318_);
  and (_22321_, _22320_, _09792_);
  or (_22322_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  or (_22323_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  and (_22324_, _22323_, _22322_);
  and (_22325_, _22324_, _05549_);
  or (_22326_, _22325_, _22321_);
  and (_22327_, _22326_, _05535_);
  or (_22328_, _22327_, _22317_);
  and (_22329_, _22328_, _05542_);
  and (_22330_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  and (_22331_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  or (_22332_, _22331_, _22330_);
  and (_22333_, _22332_, _09792_);
  and (_22334_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  and (_22335_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  or (_22336_, _22335_, _22334_);
  and (_22337_, _22336_, _05549_);
  or (_22338_, _22337_, _22333_);
  and (_22339_, _22338_, _09791_);
  and (_22340_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  and (_22341_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  or (_22342_, _22341_, _22340_);
  and (_22343_, _22342_, _09792_);
  and (_22344_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  and (_22345_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  or (_22346_, _22345_, _22344_);
  and (_22347_, _22346_, _05549_);
  or (_22348_, _22347_, _22343_);
  and (_22349_, _22348_, _05535_);
  or (_22350_, _22349_, _22339_);
  and (_22351_, _22350_, _09805_);
  or (_22352_, _22351_, _22329_);
  and (_22353_, _22352_, _05518_);
  or (_22354_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  or (_22355_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  and (_22356_, _22355_, _05549_);
  and (_22357_, _22356_, _22354_);
  or (_22358_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  or (_22359_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  and (_22360_, _22359_, _09792_);
  and (_22361_, _22360_, _22358_);
  or (_22362_, _22361_, _22357_);
  and (_22363_, _22362_, _09791_);
  or (_22364_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  or (_22365_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  and (_22366_, _22365_, _05549_);
  and (_22367_, _22366_, _22364_);
  or (_22368_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  or (_22369_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  and (_22370_, _22369_, _09792_);
  and (_22371_, _22370_, _22368_);
  or (_22372_, _22371_, _22367_);
  and (_22373_, _22372_, _05535_);
  or (_22374_, _22373_, _22363_);
  and (_22375_, _22374_, _05542_);
  and (_22376_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  and (_22377_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  or (_22378_, _22377_, _22376_);
  and (_22379_, _22378_, _09792_);
  and (_22380_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  and (_22381_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  or (_22382_, _22381_, _22380_);
  and (_22383_, _22382_, _05549_);
  or (_22384_, _22383_, _22379_);
  and (_22385_, _22384_, _09791_);
  and (_22386_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  and (_22387_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  or (_22388_, _22387_, _22386_);
  and (_22389_, _22388_, _09792_);
  and (_22390_, _09793_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  and (_22391_, _05514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  or (_22392_, _22391_, _22390_);
  and (_22393_, _22392_, _05549_);
  or (_22394_, _22393_, _22389_);
  and (_22395_, _22394_, _05535_);
  or (_22396_, _22395_, _22385_);
  and (_22397_, _22396_, _09805_);
  or (_22398_, _22397_, _22375_);
  and (_22399_, _22398_, _09850_);
  or (_22400_, _22399_, _22353_);
  and (_22401_, _22400_, _05520_);
  or (_22402_, _22401_, _22307_);
  or (_22403_, _22402_, _10033_);
  and (_22404_, _22403_, _22213_);
  or (_22405_, _22404_, _04413_);
  and (_22406_, _22405_, _22023_);
  or (_22407_, _22406_, _05563_);
  or (_22408_, _10735_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_22409_, _22408_, _22731_);
  and (_12348_, _22409_, _22407_);
  and (_22410_, _02205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_22411_, _22410_, _02306_);
  and (_22412_, _22411_, _02195_);
  nor (_22413_, _22412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_22414_, _22412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_22415_, _22414_, _22413_);
  and (_22416_, _22415_, _02198_);
  and (_22417_, _01818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_22418_, _22417_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_22419_, _11221_);
  and (_22420_, _01829_, _22419_);
  and (_22421_, _22420_, _22418_);
  or (_22422_, _11203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_22423_, _11211_, _02320_);
  and (_22424_, _22423_, _22422_);
  or (_22425_, _22424_, _22421_);
  or (_22426_, _22425_, _22416_);
  or (_22427_, _22426_, _01814_);
  nand (_22428_, _01814_, _23542_);
  and (_22429_, _22428_, _22427_);
  or (_22430_, _22429_, _01816_);
  or (_22431_, _02300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_22432_, _22431_, _22731_);
  and (_12351_, _22432_, _22430_);
  and (_22433_, _02488_, _24134_);
  and (_22434_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  or (_12353_, _22434_, _22433_);
  nand (_22435_, _01814_, _24210_);
  and (_22436_, _08225_, _02195_);
  or (_22437_, _22436_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_22438_, _11205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_22439_, _22438_, _02198_);
  and (_22440_, _22439_, _22437_);
  or (_22441_, _01818_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_22442_, _22441_, _01829_);
  nor (_22443_, _22442_, _22417_);
  or (_22444_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_22445_, _11203_, _02320_);
  and (_22446_, _22445_, _22444_);
  or (_22447_, _22446_, _22443_);
  or (_22448_, _22447_, _22440_);
  or (_22449_, _22448_, _01814_);
  and (_22450_, _22449_, _22435_);
  or (_22451_, _22450_, _01816_);
  or (_22452_, _02300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_22453_, _22452_, _22731_);
  and (_12355_, _22453_, _22451_);
  and (_22454_, _12438_, _23996_);
  and (_22455_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  or (_12357_, _22455_, _22454_);
  and (_22456_, _12438_, _24219_);
  and (_22457_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  or (_27190_, _22457_, _22456_);
  and (_22458_, _16026_, _24219_);
  and (_22459_, _16028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  or (_12369_, _22459_, _22458_);
  and (_22460_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_22461_, _01814_, _24126_);
  and (_22462_, _01825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_22463_, _22462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_22464_, _22462_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_22465_, _22464_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_22466_, _22465_, _22463_);
  and (_22467_, _02210_, _02302_);
  or (_22468_, _22467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_22469_, _02318_, _02320_);
  and (_22470_, _22469_, _22468_);
  and (_22471_, _08225_, _02302_);
  or (_22472_, _22471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_22473_, _02308_, _02197_);
  and (_22474_, _22473_, _22472_);
  or (_22475_, _22474_, _22470_);
  or (_22476_, _22475_, _22466_);
  or (_22477_, _22476_, _01814_);
  and (_22478_, _22477_, _02300_);
  and (_22479_, _22478_, _22461_);
  or (_22480_, _22479_, _22460_);
  and (_12384_, _22480_, _22731_);
  and (_22481_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_22482_, _01814_, _24043_);
  nand (_22483_, _08225_, _01823_);
  nor (_22484_, _22483_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_22485_, _22484_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not (_22486_, _22471_);
  or (_22487_, _22486_, _02196_);
  and (_22488_, _22487_, _02198_);
  and (_22489_, _22488_, _22485_);
  or (_22490_, _01824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not (_22491_, _01825_);
  and (_22492_, _01829_, _22491_);
  and (_22493_, _22492_, _22490_);
  and (_22494_, _02210_, _01823_);
  or (_22495_, _22494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_22496_, _22467_, _02320_);
  and (_22497_, _22496_, _22495_);
  or (_22498_, _22497_, _22493_);
  or (_22499_, _22498_, _22489_);
  or (_22500_, _22499_, _01814_);
  and (_22501_, _22500_, _02300_);
  and (_22502_, _22501_, _22482_);
  or (_22503_, _22502_, _22481_);
  and (_12387_, _22503_, _22731_);
  and (_22504_, _01816_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_22505_, _01814_, _24082_);
  and (_22506_, _08225_, _01822_);
  or (_22507_, _22506_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_22508_, _22483_, _02197_);
  and (_22509_, _22508_, _22507_);
  and (_22510_, _02210_, _01822_);
  or (_22511_, _22510_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_22512_, _22494_, _02320_);
  and (_22513_, _22512_, _22511_);
  and (_22514_, _01822_, _01818_);
  and (_22515_, _22514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_22516_, _22515_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_22517_, _01824_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_22518_, _22517_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_22519_, _22518_, _22516_);
  or (_22520_, _22519_, _22513_);
  or (_22521_, _22520_, _22509_);
  or (_22522_, _22521_, _01814_);
  and (_22523_, _22522_, _02300_);
  and (_22524_, _22523_, _22505_);
  or (_22525_, _22524_, _22504_);
  and (_12390_, _22525_, _22731_);
  not (_22526_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_22527_, _22414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_22528_, _22527_, _22526_);
  and (_22529_, _22527_, _22526_);
  or (_22530_, _22529_, _22528_);
  and (_22531_, _22530_, _02198_);
  or (_22532_, _11218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_22533_, _22514_);
  and (_22534_, _01829_, _22533_);
  and (_22535_, _22534_, _22532_);
  or (_22536_, _11214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_22537_, _22510_, _02320_);
  and (_22538_, _22537_, _22536_);
  or (_22539_, _22538_, _22535_);
  or (_22540_, _22539_, _01814_);
  or (_22541_, _22540_, _22531_);
  or (_22542_, _02193_, _23577_);
  and (_22543_, _22542_, _22541_);
  or (_22544_, _22543_, _01816_);
  nand (_22545_, _01816_, _22526_);
  and (_22546_, _22545_, _22731_);
  and (_12391_, _22546_, _22544_);
  and (_22547_, _25637_, _23583_);
  and (_22548_, _25640_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  or (_12393_, _22548_, _22547_);
  and (_22549_, _12438_, _23583_);
  and (_22550_, _12440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  or (_12397_, _22550_, _22549_);
  and (_22551_, _05442_, _24219_);
  and (_22552_, _05444_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  or (_12399_, _22552_, _22551_);
  and (_22553_, _03355_, _23583_);
  and (_22554_, _03357_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  or (_12404_, _22554_, _22553_);
  and (_22555_, _03033_, _23887_);
  and (_22556_, _03035_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  or (_27161_, _22556_, _22555_);
  or (_22557_, _02300_, _23880_);
  nor (_22558_, _11184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_22559_, _22558_, _11185_);
  and (_22560_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_22561_, _22560_, _22559_);
  nor (_22562_, _22561_, _01814_);
  and (_22563_, _01814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_22564_, _22563_, _22562_);
  or (_22565_, _22564_, _01816_);
  and (_22566_, _22565_, _22731_);
  and (_12412_, _22566_, _22557_);
  nand (_22567_, _01816_, _23542_);
  and (_22568_, _02205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_22569_, _22568_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_22570_, _22569_, _11184_);
  and (_22571_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_22572_, _22571_, _22570_);
  nor (_22573_, _22572_, _01814_);
  and (_22574_, _01814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_22575_, _22574_, _22573_);
  or (_22576_, _22575_, _01816_);
  and (_22577_, _22576_, _22731_);
  and (_12413_, _22577_, _22567_);
  and (_22578_, _02488_, _24051_);
  and (_22579_, _02490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  or (_12416_, _22579_, _22578_);
  nor (_22580_, _02205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_22581_, _22580_, _22568_);
  and (_22582_, _11205_, _02196_);
  nor (_22583_, _22582_, _22581_);
  nor (_22584_, _22583_, _01814_);
  and (_22585_, _01814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or (_22586_, _22585_, _22584_);
  or (_22587_, _22586_, _01816_);
  nand (_22588_, _01816_, _24210_);
  and (_22589_, _22588_, _22731_);
  and (_12417_, _22589_, _22587_);
  and (_22590_, _02045_, _24219_);
  and (_22591_, _02047_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  or (_12420_, _22591_, _22590_);
  and (_22592_, _24510_, _24219_);
  and (_22593_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  or (_12422_, _22593_, _22592_);
  and (_22594_, _24510_, _23583_);
  and (_22595_, _24512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  or (_12424_, _22595_, _22594_);
  and (_22596_, _12429_, _24219_);
  and (_22597_, _12431_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  or (_27182_, _22597_, _22596_);
  nand (_22598_, _01816_, _24082_);
  nand (_22599_, _08226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_22600_, _02210_);
  nand (_22601_, _11191_, _22600_);
  and (_22602_, _22601_, _22599_);
  nor (_22603_, _22602_, _01814_);
  or (_22604_, _22600_, _01814_);
  and (_22605_, _22604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_22606_, _22605_, _22603_);
  or (_22607_, _22606_, _01816_);
  and (_22608_, _22607_, _22731_);
  and (_12432_, _22608_, _22598_);
  and (_22609_, _03043_, _23996_);
  and (_22610_, _03045_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  or (_27252_, _22610_, _22609_);
  dff (first_instr, _00000_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _26823_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _26823_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _26823_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _26823_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _26823_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _26823_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _26823_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _26823_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _26839_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _26822_[1]);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _26822_[2]);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _26822_[3]);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _26822_[4]);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _26822_[5]);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _26822_[6]);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _26822_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _26822_[8]);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _26822_[9]);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _26822_[10]);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _26822_[11]);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _26822_[12]);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _26822_[13]);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _26822_[14]);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _26822_[15]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _26830_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _26830_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _26830_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _26830_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _26830_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _26830_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _26830_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _26830_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _26831_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _26831_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _26831_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _26831_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _26831_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _26831_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _26831_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _26831_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _26832_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _26832_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _26832_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _26832_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _26832_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _26832_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _26832_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _26832_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _26833_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _26833_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _26833_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _26833_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _26833_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _26833_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _26833_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _26833_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _26834_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _26834_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _26834_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _26834_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _26834_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _26834_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _26834_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _26834_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _26835_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _26835_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _26835_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _26835_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _26835_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _26835_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _26835_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _26835_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _26836_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _26836_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _26836_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _26836_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _26836_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _26836_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _26836_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _26836_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _26837_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _26837_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _26837_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _26837_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _26837_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _26837_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _26837_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _26837_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _26838_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _26838_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _26838_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _26838_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _26838_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _26838_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _26838_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _26838_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _26824_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _26824_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _26824_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _26824_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _26824_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _26824_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _26824_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _26824_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _26825_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _26825_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _26825_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _26825_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _26825_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _26825_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _26825_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _26825_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _26826_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _26826_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _26826_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _26826_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _26826_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _26826_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _26826_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _26826_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _26827_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _26827_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _26827_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _26827_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _26827_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _26827_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _26827_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _26827_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _26828_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _26828_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _26828_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _26828_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _26828_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _26828_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _26828_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _26828_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _26829_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _26829_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _26829_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _26829_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _26829_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _26829_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _26829_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _26829_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _11336_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _11315_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _09141_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _11283_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _11332_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _09148_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _09152_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _09133_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _11514_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _11408_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _11487_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _11475_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _11517_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _11510_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _11407_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _09145_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11708_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22676_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _11721_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _11934_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _11726_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _11738_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _11716_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11728_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _11734_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _11740_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _11736_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _11730_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _11723_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _11746_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _11742_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _11776_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _26840_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _26840_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _26840_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _26840_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _26840_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _26840_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _26840_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _26840_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _26867_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _26867_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _26867_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _26867_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _26867_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _26867_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _26867_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _26867_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _26877_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _26877_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _26877_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _26877_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _26877_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _26877_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _26877_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _26877_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _26847_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _26847_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _26848_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _26848_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _26848_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _26849_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _26849_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _26849_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _26850_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _26850_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _26851_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _26851_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _26851_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _26851_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _26852_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _26852_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _26853_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _26841_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _26841_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _26841_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _26842_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _26842_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _26842_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _26843_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _26843_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _26844_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _26844_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _26844_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _26844_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _26844_[4]);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _26844_[5]);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _26844_[6]);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _26844_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _26845_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _26846_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _26846_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _26892_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _26854_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _26854_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _26854_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _26854_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _26854_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _26854_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _26854_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _26854_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _26855_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _26855_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _26855_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _26855_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _26855_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _26855_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _26855_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _26855_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _26856_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _26856_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _26856_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _26856_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _26856_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _26856_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _26856_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _26856_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _26857_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _26857_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _26857_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _26857_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _26857_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _26857_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _26857_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _26857_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _26858_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _26858_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _26858_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _26858_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _26858_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _26858_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _26858_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _26858_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _26859_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _26859_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _26859_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _26859_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _26859_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _26859_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _26859_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _26859_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _26860_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _26860_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _26860_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _26860_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _26860_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _26860_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _26860_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _26860_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _26861_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _26861_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _26861_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _26861_[3]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _26861_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _26861_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _26861_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _26861_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _26865_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _26865_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _26865_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _26865_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _26865_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _26862_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _26862_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _26862_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _26862_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _26862_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _26862_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _26862_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _26862_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _26862_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _26862_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _26862_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _26862_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _26862_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _26862_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _26862_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _26862_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _26863_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _26863_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _26863_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _26863_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _26863_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _26863_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _26863_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _26863_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _26863_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _26863_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _26863_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _26863_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _26863_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _26863_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _26863_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _26863_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _26883_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _26883_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _26883_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _26883_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _26883_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _26883_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _26883_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _26883_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _26883_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _26883_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _26883_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _26883_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _26883_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _26883_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _26883_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _26883_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _26883_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _26883_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _26883_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _26883_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _26883_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _26883_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _26883_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _26883_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _26883_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _26883_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _26883_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _26883_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _26883_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _26883_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _26883_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _26883_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _26864_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _26866_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _26866_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _26866_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _26866_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _26866_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _26866_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _26866_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _26866_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _26868_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _26869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _26870_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _26870_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _26870_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _26870_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _26870_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _26870_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _26870_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _26870_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _26870_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _26870_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _26870_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _26870_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _26870_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _26870_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _26870_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _26870_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _26871_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _26871_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _26871_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _26871_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _26871_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _26871_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _26871_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _26871_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _26871_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _26871_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _26871_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _26871_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _26871_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _26871_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _26871_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _26871_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _26872_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _26874_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _26873_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _26875_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _26875_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _26875_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _26875_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _26875_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _26875_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _26875_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _26875_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _26876_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _26876_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _26876_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _26878_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _26879_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _26879_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _26879_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _26879_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _26879_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _26879_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _26879_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _26879_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _26880_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _26881_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _26882_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _26882_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _26882_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _26882_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _26884_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _26884_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _26884_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _26884_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _26884_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _26884_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _26884_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _26884_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _26884_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _26884_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _26884_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _26884_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _26884_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _26884_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _26884_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _26884_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _26884_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _26884_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _26884_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _26884_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _26884_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _26884_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _26884_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _26884_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _26884_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _26884_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _26884_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _26884_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _26884_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _26884_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _26884_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _26884_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _26885_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _26886_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _26887_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _26888_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _26888_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _26888_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _26888_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _26889_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _26890_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _26891_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _26891_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _26891_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _26891_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _26891_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _26891_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _26891_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _26891_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _26893_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _26893_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _26893_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _23339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _26970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _23165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _23153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _11688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _26971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _26972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _23014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _23431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _26951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _23435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _11292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _11440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _11455_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _23303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _26952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _23725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _26932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _23866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _23849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _11661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _23394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _23389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _26933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _23956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _23942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _26917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _24010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _24046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _24012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _11294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _23678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _22955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _23046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _23077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _11289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _22770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _26986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _22729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _22873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _11296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _27311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _24090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _11656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _27312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _24168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _24138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _11638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _04945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _27171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _10382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _10250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _11792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _05029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _05024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _05093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _27154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _10796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _10780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _10764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _11778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _11161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _27155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _27156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _12637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _15619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _15213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _11761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _27122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _11589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _12266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _12243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _09970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _07588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _08947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _27209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _10001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _04842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _27210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _11526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _08369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _08381_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _27207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _27208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _22681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _08629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _08634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _09980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _27205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _26065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _11383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _07499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _06869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _21620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _09230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _27206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _09896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _27203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _09891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _03584_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _27204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _06614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _07503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _03063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _09600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _09745_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _11081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _09809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _11077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _09986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _11215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _27202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _11237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _27201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _09448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _11088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _09479_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _11085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _09499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _11176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _11180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _09008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _11103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _09032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _11178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _09093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _27200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _11091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _27197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _11240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _08606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _11106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _27198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _27199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _08724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _08971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _08294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _11190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _08378_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _11109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _08397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _11188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _08490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _27196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _08087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _11115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _11222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _08123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _11113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _08142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _11192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _08169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _07645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _07762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _11121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _11224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _07812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _07923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _11117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _07944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _27305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _07972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _27306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _08275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _27307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _27308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _10812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _07968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _27300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _27301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _10720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _27302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _07975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _08814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _27303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _27304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _10607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _27299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _07983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _10656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _07981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _10671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _08290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _10688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _10534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _10562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _07990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _10583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _07988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _27298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _08694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _08855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _07997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _10379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _10446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _07995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _27296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _07993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _10508_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _27297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _10173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _27295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _08005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _10186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _10196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _10242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _08002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _10260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _08851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _09770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _27292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _09844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _08247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _27293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _08809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _27294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _10115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _08799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _10126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _10140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _09226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _27291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _09748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _09211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _03196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _06574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _27246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _27247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _22743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _22787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _22677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _22679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _08847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _10040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _10061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _08802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _10070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _27287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _08012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _27288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _10428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _26904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _10461_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _10523_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _08932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _09180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _10528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _26905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _08986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _10201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _09112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _26902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _10337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _26903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _09198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _10375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _10166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _08992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _10170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _09113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _10179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _26901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _08989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _09183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _09191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _09768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _09810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _09048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _26899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _26900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _09854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _09130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _10964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _22616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _22688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _11056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _23972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _26923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _11011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _23949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _10978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _22611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _08728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _05116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _10933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _08393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _22620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _10967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _26921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _11030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _23787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _26922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _10951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _10944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _10980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _10993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _24326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _27176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _26004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _27177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _06994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _26026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _26009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _24429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _25883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _24483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _25972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _04929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _25966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _22724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _23502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _22668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _25927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _10560_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _10899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _25953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _24432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _25993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _24423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _02554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _07425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _27174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _07399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _01662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _24390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _24498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _11442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _27175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _07511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _07501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _07550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _27172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _07554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _24191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _27173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _07306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _27169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _24199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _07868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _07646_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _27170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _08240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _07904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _24195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _09224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _09220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _09159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _24205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _08272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _08261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _08256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _08903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _24222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _27166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _27167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _27168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _00541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _09061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _09059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _09004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _10705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _10703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _00302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _10810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _24227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _10175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _00527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _27165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _24241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _11111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _27164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _11199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _10915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _10893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _10982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _00215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _11539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _11605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _11711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _11685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _26105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _11331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _27163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _11436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _12334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _12340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _24280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _11906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _12092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _11937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _24252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _24466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _02342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _05861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _27244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _22944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _10686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _22667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _27245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _10713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _26075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _26030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _27161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _26046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _23326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _27162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _12268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _12251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _02457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _12065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _02454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _27159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _27160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _02721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _10936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _10910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _06923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _02466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _07214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _02464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _05330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _27157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _11920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _27158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _22664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _22662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _02477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _22661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _27151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _27152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _27153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _02725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _27147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _22669_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _27148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _02487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _27149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _02482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _22666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _27150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _27144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _27145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _22678_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _02496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _22672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _02493_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _22671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _27146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _27142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _02736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _22723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _22686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _02510_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _22685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _02506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _27143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _25079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _27140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _22929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _02529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _22915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _27141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _22860_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _22739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _09328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _27137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _02747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _27138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _02538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _25774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _27139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _25762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _27133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _10690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _27134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _12342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _27135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _00019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _27136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _07444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _00994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _10681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _01254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _01235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _10675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _07540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _19907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _06071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _02547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _26621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _27129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _26604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _27130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _02741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _27131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _27132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _00007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _02559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _26785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _27125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _27126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _27127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _26746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _27128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _05450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _05383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _10609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _03511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _03297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _03262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _04262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _27242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _07370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _01407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _01392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _10658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _02099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _01495_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _10650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _00985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _02575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _00515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _27123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _11519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _00087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _02567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _27124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _00032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _27118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _27119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _05764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _27120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _04562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _08410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _02579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _27121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _27117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _04931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _24445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _04934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _05168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _24477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _24488_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _05052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _07544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _09691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _09688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _10589_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _09721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _07391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _05783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _05703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _06787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _07103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _27241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _07870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _07961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _04889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _04839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _04811_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _27234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _12140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _12154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _12142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _07403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _27235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _10958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _10941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _11228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _27236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _10513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _07546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _10833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _27237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _27238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _27239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _25887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _25904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _25889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _27080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _25949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _11553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _25731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _25742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _12420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _00074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _22663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _27232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _22628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _22635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _07414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _27233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _11463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _04174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _11462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _04075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _04101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _11466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _03992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _26894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _25399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _25389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _25439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _27213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _25427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _11300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _25317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _25304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _25537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _25530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _25570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _25559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _11446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _25468_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _25464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _25498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _25857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _11563_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _11390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _25667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _25653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _11592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _25702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _27189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _27258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _11630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _24435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _27259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _27260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _24338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _24335_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _24356_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _24463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _24456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _27243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _24524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _24506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _24501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _11298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _24366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _25348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _11603_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _25239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _25237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _25031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _11611_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _27228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _25265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _11632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _27289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _27290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _24211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _24202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _24288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _24285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _24256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _04958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _04962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _05005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _04954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _24213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _04863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _24215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _24183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _03336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _04487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _03509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _05113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _27116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _05089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _04873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _04914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _03352_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _04381_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _27114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _04424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _03345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _27115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _04455_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _03339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _04310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _27111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _04316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _03519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _04324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _27112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _27113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _03598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _03389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _27109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _03533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _04254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _04271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _03529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _04282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _27110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _27108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _04171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _04189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _03401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _03605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _04194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _04208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _03399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _27106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _04087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _04112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _03427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _04116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _03539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _27107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _04162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _03749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _27101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _27102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _27103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _27104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _04040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _04068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _27105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _03673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _27098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _03671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _03507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _03695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _03718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _03498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _03726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _03921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _03948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _03560_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _27097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _03969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _03989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _04007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _03456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _03477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _03848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _03475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _03854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _03627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _03864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _03918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _03467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _03761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _03486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _03768_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _03573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _03780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _03800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _03817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _03483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _04968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _25245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _25087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _24958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _27095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _25282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _25273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _27096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _25437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _04960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _25324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _25337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _25326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _04972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _25373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _27094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _04883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _24135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _24128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _24103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _24316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _24282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _24242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _27093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _25871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _25853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _25906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _24329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _24344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _04906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _24359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _24370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _25471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _05154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _27091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _25525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _27092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _25733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _25725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _25717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _23180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _02770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _25562_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _25555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _25676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _25671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _25641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _25476_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _01070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _01307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _01379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _04473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _22684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _09347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _27089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _24235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _04445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _02165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _02081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _27088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _03766_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _03648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _02773_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _01196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _04432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _09686_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _09103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _02781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _05027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _04850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _04776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _05648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _10154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _04417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _10622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _10668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _04408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _07449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _07100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _05935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _11916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _04369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _27085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _27086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _27087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _04398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _10886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _10891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _22627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _22665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _04354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _03116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _11133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _27084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _11076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _11925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _24363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _22720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _22714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _04346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _22680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _12416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _12353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _04359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _25379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _04321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _01500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _27083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _04318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _03117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _25095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _13109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _01925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _02151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _02042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _04313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _04490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _04422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _03609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _02797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _08865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _27081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _05217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _04870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _04307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _27082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _07123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _04299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _09096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _09317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _27078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _04269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _08782_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _27079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _04294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _08873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _09416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _09402_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _09391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _10048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _09743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _09544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _02808_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _09270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _11927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _27076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _27077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _10736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _10630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _10918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _10925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _02828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _08767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _05290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _04218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _22687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _04205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _03130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _11614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _11596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _03268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _02052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _02261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _02128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _04200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _04515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _04731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _04600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _04177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _06555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _07427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _06604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _04191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _10844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _09613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _04187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _08667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _02864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _27074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _01799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _23384_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _27075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _03079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _11528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _26771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _00044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _00079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _27073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _08738_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _04168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _08650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _08655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _27070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _03932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _04198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _27071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _03160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _27072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _08597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _08602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _00172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _27067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _26774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _27068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _27069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _04107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _03426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _11001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _06349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _12202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _07226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _22659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _04097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _18267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _06239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _04089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _04072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _08817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _04050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _27063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _25114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _23315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _27064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _27065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _04026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _27057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _27058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _27059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _27060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _27061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _27062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _18155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _27056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _23993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _25749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _25595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _11326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _11496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _04037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _09147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _27053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _23200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _27054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _03099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _27055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _03753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _03741_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _03240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _08023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _09950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _09966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _09974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _27285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _10008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _08020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _27286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _25624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _25474_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _25419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _10968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _27284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _09886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _09908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _08238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _25843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _27280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _27281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _27282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _27283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _24901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _24796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _24683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _00972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _05091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _10950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _22622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _27278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _27279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _25824_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _25943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _10948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _03395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _06732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _04137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _10938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _22614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _25847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _10955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _27274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _27275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _27276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _27277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _11036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _22689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _11173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _09287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _27268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _27269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _27270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _27271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _27272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _27273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _11048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _11017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _10838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _07338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _07626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _27263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _27264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _27265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _27266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _27267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _10901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _10999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _11014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _27261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _03548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _27262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _10820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _10866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _07346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _27257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _11071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _11156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _11144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _11124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _07344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _10897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _11752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _11694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _07353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _27256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _11242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _11220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _11369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _11303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _27253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _09331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _09427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _27254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _11601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _27255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _11452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _11425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _09666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _09662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _09649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _27251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _12148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _23365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _07355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _27252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _27249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _27250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _08400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _08408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _08949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _26817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _00022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _00082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _27248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _07360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _26728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _26685_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _26725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _25076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _25082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _25747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _22623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _10090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _11550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _11594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _27217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _11658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _11902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _10111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _11213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _05882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _05940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _11167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _11234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _07386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _07614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _27195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _27214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _23135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _00674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _27215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _07565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _27216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _26078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _10097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _07199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _11126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _07223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _11200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _07276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _07366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _05608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _11172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _10059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _07580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _03443_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _27212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _04814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _07462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _04780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _22645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _11204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _06772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _11135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _06814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _11202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _06894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _07047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _11128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _07898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _10818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _10928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _23110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _10043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _06806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _27211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _09412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _06304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _11146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _11232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _06382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _06622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _27193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _27194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _06722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _12422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _04624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _04621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _12424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _06025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _06076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _27192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _06235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _12399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _26661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _04365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _12274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _04371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _04588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _12332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _04591_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _27190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _27191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _04655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _12397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _04728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _04720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _04713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _12357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _04857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _04788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _04784_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _04771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _27188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _04836_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _04834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _04822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _04296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _04284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _04415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _04411_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _04391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _27186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _04351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _27187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _27185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _04453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _04457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _12293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _04509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _04546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _04511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _12280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _27182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _27183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _27184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _05143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _05206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _05187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _09513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _04618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _05064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _27179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _04922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _04919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _04911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _27180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _04963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _27181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _22658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _27019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _22674_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _22673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _11285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _22651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _27020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _27021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _27099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _11759_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _18441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _18950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _11757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _11375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _12748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _27100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _10953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _10942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _10984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _10995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _11005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _10976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _27310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _09884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _03123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _27023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _05607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _03125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _03154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _05189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _03163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _03179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _05466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _25452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _22879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _23021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _22959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _03095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _27024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _22798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _06948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _06955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _27008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _03418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _26029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _05445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _26033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _27009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _10923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _06340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _06086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _10431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _10434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _06346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _10739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _26959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _26960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _10151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _06350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _26961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _10194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _05917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _06179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _12261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _11021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _06336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _26957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _05932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _10828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _10864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _10831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _26958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _26934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _10506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _07043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _10539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _07197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _10569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _26935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _07037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _07965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _08812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _11043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _27309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _11023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _11039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _11024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _10946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _10881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _27240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _10883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _07397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _10599_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _10574_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _10716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _10711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _27230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _25352_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _06338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _03576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _14268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _27231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _08017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _04393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _01504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _01404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _23102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _22939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _10366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _25037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _25170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _27229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _27224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _09017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _09014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _10181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _07180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _27225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _10190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _07513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _02030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _10244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _02327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _03156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _10214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _26052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _00657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _00289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _27226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _04504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _04525_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _04506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _05470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _05135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _10198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _27227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _23171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _27219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _24346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _25875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _25960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _09807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _27220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _09846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _27222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _09268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _09256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _10177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _27223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _09276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _07433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _08825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _06088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _06268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _01224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _07506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _07910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _09367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _09357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _27221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _10613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _10577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _10551_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _09063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _09735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _09996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _09218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _06207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _18176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _07515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _10974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _12393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _09214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _01301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _09207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _07912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _19605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _27090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _19639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _21642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _21519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _21388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _11754_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _17998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _11714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _22615_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _22613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _22612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _22621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _22619_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _22618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _11750_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _22657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _22655_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _11696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _27037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _22638_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _22637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _27038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _22648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _22647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _11699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _11380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _11450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _27066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _22625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _22630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _22634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _27007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _11287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _11439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _22683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _22682_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _11691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _22721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _22717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _03664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _03300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _03704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _23428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _03701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _23307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _27052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _23332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _26270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _26134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _27047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _27048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _27049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _04005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _03177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _23852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _23961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _03675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _27050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _27051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _03103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _24049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _24007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _24084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _27042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _03971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _27043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _27044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _03999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _27045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _27046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _03994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _27036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _12616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _12515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _03056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _10727_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _10814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _11416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _03924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _27039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _03961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _06056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _06601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _03051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _27040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _27041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _03986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _07894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _08331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _08103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _10347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _10107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _10012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _03053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _05303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _27033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _03856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _03216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _15234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _15162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _03907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _27034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _27035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _03827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _22636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _03064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _27030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _27031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _22617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _27032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _19201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _03804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _22646_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _27028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _27029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _22654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _22650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _03812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _22626_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _05238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _03069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _05474_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _05714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _03076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _27022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _05222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _03112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _03092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _27025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _22675_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _27026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _22713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _27027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _22656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _22660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _27016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _02853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _02878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _27017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _05644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _27018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _05272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _02933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _03000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _05252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _03012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _05503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _03027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _05245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _03047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _05483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _01604_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _27014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _01606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _27015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _05283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _05650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _02822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _02850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _00299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _05336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _00305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _05557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _00310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _00596_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _05325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _01600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _27013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _00270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _05354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _00276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _05564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _00280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _00291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _05346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _05581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _00203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _05369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _00209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _05575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _00212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _00262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _05357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _05729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _25996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _26012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _05452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _26015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _26019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _05447_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _05695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _27012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _05588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _26086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _05390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _26096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _05586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _26117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _00103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _03422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _03415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _06558_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _03480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _03472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _05778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _27005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _27006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _05433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _27010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _27011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _26056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _05423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _26062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _05590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _26069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _03342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _03321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _25946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _25939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _06569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _03223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _03206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _06564_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _03820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _05781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _03553_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _27002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _03631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _27003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _27004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _03440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _04013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _27001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _03974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _05786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _03659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _03716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _03697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _03836_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _04055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _04185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _04165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _04159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _06530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _27000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _03867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _03900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _04279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _04273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _26998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _26999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _04386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _06519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _04109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _04092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _07117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _07083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _01698_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _27178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _01688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _06928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _06897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _01729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _26995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _04492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _04471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _26996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _04576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _04571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _26997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _06147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _06485_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _26993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _26994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _04679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _04664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _04734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _04765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _04740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _05166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _06477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _05241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _05220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _05812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _06149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _26988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _04966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _26989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _26990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _26991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _04817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _04845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _26992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _04927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _04917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _05740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _05718_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _05320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _26987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _05794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _05788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _06467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _05172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _06457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _06059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _05820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _05840_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _05833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _06462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _05928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _06459_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _06123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _06107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _26984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _26985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _05825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _06151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _06021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _05998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _06434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _06380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _06408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _06396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _06444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _26982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _06465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _06439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _06280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _06266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _06248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _26983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _06333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _06327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _06314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _06445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _06428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _06068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _26980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _06547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _06541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _06436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _26981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _06627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _06886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _06881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _06420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _06667_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _06707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _06744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _06760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _26979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _07010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _07049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _07039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _26976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _26977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _06823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _06817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _26978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _06401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _07270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _07266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _07251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _07349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _07341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _26974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _05859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _07125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _07115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _07089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _07204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _07185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _26975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _06964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _06960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _07607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _07586_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _05866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _26973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _07407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _07394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _06403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _07471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _06169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _07648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _26969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _07908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _07902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _06390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _07542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _07528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _09056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _09002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _05909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _08253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _08249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _08280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _08278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _06373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _06225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _06214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _26966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _26967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _10003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _10050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _26968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _05913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _09122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _09069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _09788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _09232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _09228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _06355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _08905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _08862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _01388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _26963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _04126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _26964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _26965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _00184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _25957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _02533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _26962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _06229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _10970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _11914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _06232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _06120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _06243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _10653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _26953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _26954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _26955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _11162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _11142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _11262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _11249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _26956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _11795_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _11909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _05945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _11512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _06309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _11641_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _26950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _11357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _12369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _12344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _05951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _11932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _26949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _12224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _06297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _06095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _11627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _06285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _26948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _06288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _10420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _05974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _10921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _10694_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _08780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _24419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _05960_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _12404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _24475_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _05676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _05954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _12301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _05892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _06275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _05981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _11654_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _06282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _06277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _26947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _11074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _26942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _26943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _06983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _26944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _06978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _26945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _26946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _10826_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _07317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _10639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _07033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _26936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _07194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _10648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _10692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _26937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _10723_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _10734_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _26938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _07003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _26939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _07188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _26940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _26941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _09119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _07061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _09157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _07059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _09196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _07201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _09201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _09755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _07216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _07959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _08259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _07075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _07297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _08284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _08912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _26931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _07081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _07300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _05175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _26926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _07164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _05163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _26927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _05379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _26928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _26929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _26930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _05978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _07245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _07324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _07535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _07952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _07221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _07293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _07232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _07418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _07456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _07094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _07469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _07092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _07113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _07051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _26924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _07054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _26925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _07145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _07107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _07177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _06045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _07141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _06054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _06065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _06414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _07130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _07309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _06416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _26918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _09057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _26919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _26920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _08887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _09139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _11042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _11050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _26911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _08896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _26912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _26913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _26914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _26915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _08892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _26916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _10645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _26906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _26907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _26908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _10696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _26909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _10747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _26910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _10093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _10113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _26897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _10144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _08995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _09216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _26898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _09209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _27218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _10853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _11170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _11305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _11197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _09977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _09664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _09630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _09108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _10572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _10601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _08925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _09177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _10618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _08923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _10624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _10018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _09034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _09188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _10045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _09009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _10055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _26896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _08999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _26895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _09939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _09953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _09042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _09961_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _09972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _09038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _10006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _11068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _04666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _04746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _04805_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _04717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _04460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _27313_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _12348_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _27314_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _27315_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _27315_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _27315_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _27315_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _27316_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _27317_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _27318_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _27318_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _27318_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _27318_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _27318_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _27318_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _27318_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _27318_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _10454_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _10442_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _10266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _10304_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _10358_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _10324_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _10220_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _10147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _06501_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _06506_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _06504_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _06511_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _06517_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _06514_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _06526_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _05463_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _09920_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _09918_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _09881_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _09875_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _09864_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _09741_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _09959_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _09766_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _09776_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _09911_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _09837_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _09800_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _09916_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _09914_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _09835_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _09929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _11411_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _22640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _09539_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _09650_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _09621_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _09580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _09560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _22639_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _11486_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _08845_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _11258_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _11366_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _08746_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _22642_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _11334_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _09118_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _22641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _11328_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _08233_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _08572_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _11352_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _11268_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _11347_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _11310_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _07742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _07723_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _07703_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _11322_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _07156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _06967_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _07135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _07072_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _07024_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _22643_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _07479_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _11372_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _06560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _06536_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _06510_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _06442_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _22644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _06793_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _06752_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _11355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _11669_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _11644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _11618_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _05791_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _11994_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _11891_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _11973_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _10870_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _11035_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _10987_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _10960_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _10934_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _05805_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _11356_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _11255_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _10857_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _10592_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _10460_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _10565_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _10541_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _10516_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _10482_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _05816_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _10753_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _09922_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _09894_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _09868_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _09786_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _05843_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _10293_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _10136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _10842_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _10161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _10130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _10118_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _10102_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _10120_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _10132_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _09826_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _06681_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _06980_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _06974_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _06992_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _06988_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _06990_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _06999_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _06997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _06701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _22716_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _03359_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _04010_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _05666_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _05602_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _04002_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _01093_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _11027_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _10620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _22697_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _04015_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _05476_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _05019_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _09955_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _08662_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _06161_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _22670_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _09079_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _22652_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _09462_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _12417_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _12413_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _12412_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _04044_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _12432_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _07109_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _02667_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _22649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _12355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _12351_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _04046_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _12391_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _12390_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _12387_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _12384_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _22653_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _22624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _12325_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _12316_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _04077_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _05477_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _26179_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _09136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _24427_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _02924_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _18134_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _18119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _18105_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _17956_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _08907_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02719_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _07409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _08711_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _08701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _08288_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02751_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _17942_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02766_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _08270_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _08268_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _08266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02763_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _08242_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _08237_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _17922_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _17853_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _07896_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _07891_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _07889_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02788_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _07917_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _07905_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _07914_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _17818_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _07875_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _07884_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _07881_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _07879_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _07877_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02791_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _07624_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _17768_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _17752_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _07639_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02805_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _07577_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _07562_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _07558_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02843_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _07603_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _17618_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _22883_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _22895_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _22892_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _22889_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _22722_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _22765_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _22715_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _22718_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _22719_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _22725_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _22727_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01368_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _01336_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _25690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _25688_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _01421_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _25708_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _25706_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _22748_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _01409_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _22726_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _22728_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _22807_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _01334_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _22632_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _22633_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _22842_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _22631_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _22870_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _22819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _22848_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _01355_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _25655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _25638_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _25646_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _01426_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _22730_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _22754_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _22756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _25680_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _22712_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _22711_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _22710_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _22709_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _22708_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _22707_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _22706_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _22705_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _22704_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _22703_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _25678_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _22702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _22701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _22629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _22700_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _26109_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _22699_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _22698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _01423_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _22696_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _22695_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _22694_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _22693_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _22692_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _22691_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _22690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _01332_);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
endmodule
