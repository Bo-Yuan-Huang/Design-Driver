
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, property_invalid_rom_pc, property_invalid_dec_rom_pc, property_invalid_pc, property_invalid_acc, property_invalid_b_reg, property_invalid_dpl, property_invalid_dph, property_invalid_iram, property_invalid_p0, property_invalid_p1, property_invalid_p2, property_invalid_p3, property_invalid_psw, property_invalid_sp);
  wire _00000_;
  wire _00001_;
  wire [7:0] _00002_;
  wire [7:0] _00003_;
  wire [7:0] _00004_;
  wire [7:0] _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire [7:0] _35582_;
  wire _35583_;
  wire [7:0] _35584_;
  wire _35585_;
  wire [7:0] _35586_;
  wire _35587_;
  wire [7:0] _35588_;
  wire _35589_;
  wire [7:0] _35590_;
  wire _35591_;
  wire [7:0] _35592_;
  wire _35593_;
  wire [7:0] _35594_;
  wire _35595_;
  wire [7:0] _35596_;
  wire _35597_;
  wire [7:0] _35598_;
  wire _35599_;
  wire [7:0] _35600_;
  wire _35601_;
  wire [7:0] _35602_;
  wire _35603_;
  wire [7:0] _35604_;
  wire _35605_;
  wire [7:0] _35606_;
  wire _35607_;
  wire [7:0] _35608_;
  wire _35609_;
  wire [7:0] _35610_;
  wire _35611_;
  wire [7:0] _35612_;
  wire _35613_;
  wire [7:0] _35614_;
  wire [7:0] _35615_;
  wire [7:0] _35616_;
  wire [7:0] _35617_;
  wire [7:0] _35618_;
  wire [7:0] _35619_;
  wire [7:0] _35620_;
  wire [7:0] _35621_;
  wire [7:0] _35622_;
  wire [7:0] _35623_;
  wire [7:0] _35624_;
  wire [7:0] _35625_;
  wire [7:0] _35626_;
  wire [7:0] _35627_;
  wire [7:0] _35628_;
  wire [15:0] _35629_;
  wire [7:0] _35630_;
  wire [7:0] _35631_;
  wire [7:0] _35632_;
  wire [7:0] _35633_;
  wire [7:0] _35634_;
  wire [7:0] _35635_;
  wire [7:0] _35636_;
  wire [7:0] _35637_;
  wire [7:0] _35638_;
  wire [7:0] _35639_;
  wire [15:0] _35640_;
  wire [7:0] _35641_;
  wire [7:0] _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire [1:0] _35771_;
  wire [5:0] _35772_;
  wire [7:0] _35773_;
  wire [1:0] _35774_;
  wire [15:0] _35775_;
  wire [7:0] _35776_;
  wire [7:0] _35777_;
  wire [7:0] _35778_;
  wire [2:0] _35779_;
  wire [2:0] _35780_;
  wire [1:0] _35781_;
  wire [7:0] _35782_;
  wire _35783_;
  wire [1:0] _35784_;
  wire [1:0] _35785_;
  wire [2:0] _35786_;
  wire [2:0] _35787_;
  wire [1:0] _35788_;
  wire [3:0] _35789_;
  wire [1:0] _35790_;
  wire _35791_;
  wire _35792_;
  wire [15:0] _35793_;
  wire [15:0] _35794_;
  wire _35795_;
  wire [4:0] _35796_;
  wire [7:0] _35797_;
  wire [7:0] _35798_;
  wire [7:0] _35799_;
  wire _35800_;
  wire _35801_;
  wire [7:0] _35802_;
  wire [15:0] _35803_;
  wire [15:0] _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire [7:0] _35808_;
  wire [2:0] _35809_;
  wire [7:0] _35810_;
  wire [7:0] _35811_;
  wire _35812_;
  wire [7:0] _35813_;
  wire _35814_;
  wire _35815_;
  wire [3:0] _35816_;
  wire [31:0] _35817_;
  wire [31:0] _35818_;
  wire [7:0] _35819_;
  wire _35820_;
  wire _35821_;
  wire [15:0] _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire [15:0] _35826_;
  wire _35827_;
  wire _35828_;
  wire [7:0] _35829_;
  wire _35830_;
  wire [2:0] _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire [7:0] _35960_;
  wire _35961_;
  wire _35962_;
  wire [7:0] _35963_;
  wire _35964_;
  wire [7:0] _35965_;
  wire [7:0] _35966_;
  wire [7:0] _35967_;
  wire [7:0] _35968_;
  wire [7:0] _35969_;
  wire [7:0] _35970_;
  wire [7:0] _35971_;
  wire [7:0] _35972_;
  wire [6:0] _35973_;
  wire _35974_;
  wire [7:0] _35975_;
  wire [7:0] ACC_gm;
  wire [7:0] B_gm;
  wire [7:0] DPH_gm;
  wire [7:0] DPL_gm;
  wire [7:0] IE_gm;
  wire [7:0] IE_gm_next;
  wire [7:0] IP_gm;
  wire [7:0] IP_gm_next;
  wire [7:0] P0_gm;
  wire [7:0] P1_gm;
  wire [7:0] P2_gm;
  wire [7:0] P3_gm;
  wire [7:0] PCON_gm;
  wire [7:0] PCON_gm_next;
  wire [15:0] PC_gm;
  wire [7:0] PSW_gm;
  wire [7:0] SBUF_gm;
  wire [7:0] SBUF_gm_next;
  wire [7:0] SCON_gm;
  wire [7:0] SCON_gm_next;
  wire [7:0] SP_gm;
  wire [7:0] TCON_gm;
  wire [7:0] TCON_gm_next;
  wire [7:0] TH0_gm;
  wire [7:0] TH0_gm_next;
  wire [7:0] TH1_gm;
  wire [7:0] TH1_gm_next;
  wire [7:0] TL0_gm;
  wire [7:0] TL0_gm_next;
  wire [7:0] TL1_gm;
  wire [7:0] TL1_gm_next;
  wire [7:0] TMOD_gm;
  wire [7:0] TMOD_gm_next;
  wire [7:0] acc_impl;
  wire [7:0] b_reg_impl;
  input clk;
  wire [31:0] cxrom_data_out;
  wire [15:0] dptr_impl;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e0 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e2 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e3 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e7 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IE_next ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IP_next ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P0INREG ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P1INREG ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P2INREG ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [7:0] \oc8051_golden_model_1.P3INREG ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [7:0] \oc8051_golden_model_1.PCON_next ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_00 ;
  wire [7:0] \oc8051_golden_model_1.PSW_01 ;
  wire [7:0] \oc8051_golden_model_1.PSW_02 ;
  wire [7:0] \oc8051_golden_model_1.PSW_03 ;
  wire [7:0] \oc8051_golden_model_1.PSW_04 ;
  wire [7:0] \oc8051_golden_model_1.PSW_06 ;
  wire [7:0] \oc8051_golden_model_1.PSW_07 ;
  wire [7:0] \oc8051_golden_model_1.PSW_08 ;
  wire [7:0] \oc8051_golden_model_1.PSW_09 ;
  wire [7:0] \oc8051_golden_model_1.PSW_0a ;
  wire [7:0] \oc8051_golden_model_1.PSW_0b ;
  wire [7:0] \oc8051_golden_model_1.PSW_0c ;
  wire [7:0] \oc8051_golden_model_1.PSW_0d ;
  wire [7:0] \oc8051_golden_model_1.PSW_0e ;
  wire [7:0] \oc8051_golden_model_1.PSW_0f ;
  wire [7:0] \oc8051_golden_model_1.PSW_11 ;
  wire [7:0] \oc8051_golden_model_1.PSW_12 ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_14 ;
  wire [7:0] \oc8051_golden_model_1.PSW_16 ;
  wire [7:0] \oc8051_golden_model_1.PSW_17 ;
  wire [7:0] \oc8051_golden_model_1.PSW_18 ;
  wire [7:0] \oc8051_golden_model_1.PSW_19 ;
  wire [7:0] \oc8051_golden_model_1.PSW_1a ;
  wire [7:0] \oc8051_golden_model_1.PSW_1b ;
  wire [7:0] \oc8051_golden_model_1.PSW_1c ;
  wire [7:0] \oc8051_golden_model_1.PSW_1d ;
  wire [7:0] \oc8051_golden_model_1.PSW_1e ;
  wire [7:0] \oc8051_golden_model_1.PSW_1f ;
  wire [7:0] \oc8051_golden_model_1.PSW_20 ;
  wire [7:0] \oc8051_golden_model_1.PSW_21 ;
  wire [7:0] \oc8051_golden_model_1.PSW_22 ;
  wire [7:0] \oc8051_golden_model_1.PSW_23 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_30 ;
  wire [7:0] \oc8051_golden_model_1.PSW_31 ;
  wire [7:0] \oc8051_golden_model_1.PSW_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_40 ;
  wire [7:0] \oc8051_golden_model_1.PSW_41 ;
  wire [7:0] \oc8051_golden_model_1.PSW_42 ;
  wire [7:0] \oc8051_golden_model_1.PSW_44 ;
  wire [7:0] \oc8051_golden_model_1.PSW_45 ;
  wire [7:0] \oc8051_golden_model_1.PSW_46 ;
  wire [7:0] \oc8051_golden_model_1.PSW_47 ;
  wire [7:0] \oc8051_golden_model_1.PSW_48 ;
  wire [7:0] \oc8051_golden_model_1.PSW_49 ;
  wire [7:0] \oc8051_golden_model_1.PSW_4a ;
  wire [7:0] \oc8051_golden_model_1.PSW_4b ;
  wire [7:0] \oc8051_golden_model_1.PSW_4c ;
  wire [7:0] \oc8051_golden_model_1.PSW_4d ;
  wire [7:0] \oc8051_golden_model_1.PSW_4e ;
  wire [7:0] \oc8051_golden_model_1.PSW_4f ;
  wire [7:0] \oc8051_golden_model_1.PSW_50 ;
  wire [7:0] \oc8051_golden_model_1.PSW_51 ;
  wire [7:0] \oc8051_golden_model_1.PSW_52 ;
  wire [7:0] \oc8051_golden_model_1.PSW_54 ;
  wire [7:0] \oc8051_golden_model_1.PSW_55 ;
  wire [7:0] \oc8051_golden_model_1.PSW_56 ;
  wire [7:0] \oc8051_golden_model_1.PSW_57 ;
  wire [7:0] \oc8051_golden_model_1.PSW_58 ;
  wire [7:0] \oc8051_golden_model_1.PSW_59 ;
  wire [7:0] \oc8051_golden_model_1.PSW_5a ;
  wire [7:0] \oc8051_golden_model_1.PSW_5b ;
  wire [7:0] \oc8051_golden_model_1.PSW_5c ;
  wire [7:0] \oc8051_golden_model_1.PSW_5d ;
  wire [7:0] \oc8051_golden_model_1.PSW_5e ;
  wire [7:0] \oc8051_golden_model_1.PSW_5f ;
  wire [7:0] \oc8051_golden_model_1.PSW_60 ;
  wire [7:0] \oc8051_golden_model_1.PSW_61 ;
  wire [7:0] \oc8051_golden_model_1.PSW_64 ;
  wire [7:0] \oc8051_golden_model_1.PSW_65 ;
  wire [7:0] \oc8051_golden_model_1.PSW_66 ;
  wire [7:0] \oc8051_golden_model_1.PSW_67 ;
  wire [7:0] \oc8051_golden_model_1.PSW_68 ;
  wire [7:0] \oc8051_golden_model_1.PSW_69 ;
  wire [7:0] \oc8051_golden_model_1.PSW_6a ;
  wire [7:0] \oc8051_golden_model_1.PSW_6b ;
  wire [7:0] \oc8051_golden_model_1.PSW_6c ;
  wire [7:0] \oc8051_golden_model_1.PSW_6d ;
  wire [7:0] \oc8051_golden_model_1.PSW_6e ;
  wire [7:0] \oc8051_golden_model_1.PSW_6f ;
  wire [7:0] \oc8051_golden_model_1.PSW_70 ;
  wire [7:0] \oc8051_golden_model_1.PSW_71 ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_73 ;
  wire [7:0] \oc8051_golden_model_1.PSW_74 ;
  wire [7:0] \oc8051_golden_model_1.PSW_76 ;
  wire [7:0] \oc8051_golden_model_1.PSW_77 ;
  wire [7:0] \oc8051_golden_model_1.PSW_78 ;
  wire [7:0] \oc8051_golden_model_1.PSW_79 ;
  wire [7:0] \oc8051_golden_model_1.PSW_7a ;
  wire [7:0] \oc8051_golden_model_1.PSW_7b ;
  wire [7:0] \oc8051_golden_model_1.PSW_7c ;
  wire [7:0] \oc8051_golden_model_1.PSW_7d ;
  wire [7:0] \oc8051_golden_model_1.PSW_7e ;
  wire [7:0] \oc8051_golden_model_1.PSW_7f ;
  wire [7:0] \oc8051_golden_model_1.PSW_80 ;
  wire [7:0] \oc8051_golden_model_1.PSW_81 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_83 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_90 ;
  wire [7:0] \oc8051_golden_model_1.PSW_91 ;
  wire [7:0] \oc8051_golden_model_1.PSW_93 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_aa ;
  wire [7:0] \oc8051_golden_model_1.PSW_ab ;
  wire [7:0] \oc8051_golden_model_1.PSW_ac ;
  wire [7:0] \oc8051_golden_model_1.PSW_ad ;
  wire [7:0] \oc8051_golden_model_1.PSW_ae ;
  wire [7:0] \oc8051_golden_model_1.PSW_af ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_c9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ca ;
  wire [7:0] \oc8051_golden_model_1.PSW_cb ;
  wire [7:0] \oc8051_golden_model_1.PSW_cc ;
  wire [7:0] \oc8051_golden_model_1.PSW_cd ;
  wire [7:0] \oc8051_golden_model_1.PSW_ce ;
  wire [7:0] \oc8051_golden_model_1.PSW_cf ;
  wire [7:0] \oc8051_golden_model_1.PSW_d1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_da ;
  wire [7:0] \oc8051_golden_model_1.PSW_db ;
  wire [7:0] \oc8051_golden_model_1.PSW_dc ;
  wire [7:0] \oc8051_golden_model_1.PSW_dd ;
  wire [7:0] \oc8051_golden_model_1.PSW_de ;
  wire [7:0] \oc8051_golden_model_1.PSW_df ;
  wire [7:0] \oc8051_golden_model_1.PSW_e0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_e9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ea ;
  wire [7:0] \oc8051_golden_model_1.PSW_eb ;
  wire [7:0] \oc8051_golden_model_1.PSW_ec ;
  wire [7:0] \oc8051_golden_model_1.PSW_ed ;
  wire [7:0] \oc8051_golden_model_1.PSW_ee ;
  wire [7:0] \oc8051_golden_model_1.PSW_ef ;
  wire [7:0] \oc8051_golden_model_1.PSW_f0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f1 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_f9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_fa ;
  wire [7:0] \oc8051_golden_model_1.PSW_fb ;
  wire [7:0] \oc8051_golden_model_1.PSW_fc ;
  wire [7:0] \oc8051_golden_model_1.PSW_fd ;
  wire [7:0] \oc8051_golden_model_1.PSW_fe ;
  wire [7:0] \oc8051_golden_model_1.PSW_ff ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SBUF_next ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SCON_next ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TCON_next ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH0_next ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TH1_next ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL0_next ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TL1_next ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire [7:0] \oc8051_golden_model_1.TMOD_next ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_e0 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_e2 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_e3 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_f0 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_f2 ;
  wire [15:0] \oc8051_golden_model_1.XRAM_ADDR_f3 ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_IN ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT_f0 ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT_f2 ;
  wire [7:0] \oc8051_golden_model_1.XRAM_DATA_OUT_f3 ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0573 ;
  wire [7:0] \oc8051_golden_model_1.n0606 ;
  wire [15:0] \oc8051_golden_model_1.n0713 ;
  wire [15:0] \oc8051_golden_model_1.n0745 ;
  wire [6:0] \oc8051_golden_model_1.n1002 ;
  wire \oc8051_golden_model_1.n1003 ;
  wire \oc8051_golden_model_1.n1004 ;
  wire \oc8051_golden_model_1.n1005 ;
  wire \oc8051_golden_model_1.n1006 ;
  wire \oc8051_golden_model_1.n1007 ;
  wire \oc8051_golden_model_1.n1008 ;
  wire \oc8051_golden_model_1.n1009 ;
  wire \oc8051_golden_model_1.n1010 ;
  wire \oc8051_golden_model_1.n1017 ;
  wire [7:0] \oc8051_golden_model_1.n1018 ;
  wire [7:0] \oc8051_golden_model_1.n1025 ;
  wire \oc8051_golden_model_1.n1026 ;
  wire \oc8051_golden_model_1.n1027 ;
  wire \oc8051_golden_model_1.n1028 ;
  wire \oc8051_golden_model_1.n1029 ;
  wire \oc8051_golden_model_1.n1030 ;
  wire \oc8051_golden_model_1.n1031 ;
  wire \oc8051_golden_model_1.n1032 ;
  wire \oc8051_golden_model_1.n1033 ;
  wire \oc8051_golden_model_1.n1040 ;
  wire [7:0] \oc8051_golden_model_1.n1041 ;
  wire \oc8051_golden_model_1.n1057 ;
  wire [7:0] \oc8051_golden_model_1.n1058 ;
  wire [3:0] \oc8051_golden_model_1.n1139 ;
  wire [3:0] \oc8051_golden_model_1.n1141 ;
  wire [3:0] \oc8051_golden_model_1.n1143 ;
  wire [3:0] \oc8051_golden_model_1.n1144 ;
  wire [3:0] \oc8051_golden_model_1.n1145 ;
  wire [3:0] \oc8051_golden_model_1.n1146 ;
  wire [3:0] \oc8051_golden_model_1.n1147 ;
  wire [3:0] \oc8051_golden_model_1.n1148 ;
  wire [3:0] \oc8051_golden_model_1.n1149 ;
  wire \oc8051_golden_model_1.n1195 ;
  wire \oc8051_golden_model_1.n1237 ;
  wire [8:0] \oc8051_golden_model_1.n1238 ;
  wire [8:0] \oc8051_golden_model_1.n1239 ;
  wire [7:0] \oc8051_golden_model_1.n1240 ;
  wire \oc8051_golden_model_1.n1241 ;
  wire [2:0] \oc8051_golden_model_1.n1242 ;
  wire \oc8051_golden_model_1.n1243 ;
  wire [1:0] \oc8051_golden_model_1.n1244 ;
  wire [7:0] \oc8051_golden_model_1.n1245 ;
  wire [6:0] \oc8051_golden_model_1.n1246 ;
  wire \oc8051_golden_model_1.n1247 ;
  wire \oc8051_golden_model_1.n1248 ;
  wire \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1251 ;
  wire \oc8051_golden_model_1.n1252 ;
  wire \oc8051_golden_model_1.n1253 ;
  wire \oc8051_golden_model_1.n1254 ;
  wire \oc8051_golden_model_1.n1261 ;
  wire [7:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1278 ;
  wire [7:0] \oc8051_golden_model_1.n1279 ;
  wire [15:0] \oc8051_golden_model_1.n1310 ;
  wire [7:0] \oc8051_golden_model_1.n1312 ;
  wire \oc8051_golden_model_1.n1313 ;
  wire \oc8051_golden_model_1.n1314 ;
  wire \oc8051_golden_model_1.n1315 ;
  wire \oc8051_golden_model_1.n1316 ;
  wire \oc8051_golden_model_1.n1317 ;
  wire \oc8051_golden_model_1.n1318 ;
  wire \oc8051_golden_model_1.n1319 ;
  wire \oc8051_golden_model_1.n1320 ;
  wire \oc8051_golden_model_1.n1327 ;
  wire [7:0] \oc8051_golden_model_1.n1328 ;
  wire [8:0] \oc8051_golden_model_1.n1330 ;
  wire [8:0] \oc8051_golden_model_1.n1334 ;
  wire \oc8051_golden_model_1.n1335 ;
  wire [3:0] \oc8051_golden_model_1.n1336 ;
  wire [4:0] \oc8051_golden_model_1.n1337 ;
  wire [4:0] \oc8051_golden_model_1.n1341 ;
  wire \oc8051_golden_model_1.n1342 ;
  wire [8:0] \oc8051_golden_model_1.n1343 ;
  wire \oc8051_golden_model_1.n1351 ;
  wire [7:0] \oc8051_golden_model_1.n1352 ;
  wire [6:0] \oc8051_golden_model_1.n1353 ;
  wire \oc8051_golden_model_1.n1368 ;
  wire [7:0] \oc8051_golden_model_1.n1369 ;
  wire [8:0] \oc8051_golden_model_1.n1392 ;
  wire \oc8051_golden_model_1.n1393 ;
  wire [4:0] \oc8051_golden_model_1.n1398 ;
  wire \oc8051_golden_model_1.n1399 ;
  wire \oc8051_golden_model_1.n1407 ;
  wire [7:0] \oc8051_golden_model_1.n1408 ;
  wire [6:0] \oc8051_golden_model_1.n1409 ;
  wire \oc8051_golden_model_1.n1424 ;
  wire [7:0] \oc8051_golden_model_1.n1425 ;
  wire [8:0] \oc8051_golden_model_1.n1427 ;
  wire [8:0] \oc8051_golden_model_1.n1429 ;
  wire \oc8051_golden_model_1.n1430 ;
  wire [3:0] \oc8051_golden_model_1.n1431 ;
  wire [4:0] \oc8051_golden_model_1.n1432 ;
  wire [4:0] \oc8051_golden_model_1.n1434 ;
  wire \oc8051_golden_model_1.n1435 ;
  wire [8:0] \oc8051_golden_model_1.n1436 ;
  wire \oc8051_golden_model_1.n1443 ;
  wire [7:0] \oc8051_golden_model_1.n1444 ;
  wire [6:0] \oc8051_golden_model_1.n1445 ;
  wire \oc8051_golden_model_1.n1460 ;
  wire [7:0] \oc8051_golden_model_1.n1461 ;
  wire [8:0] \oc8051_golden_model_1.n1463 ;
  wire \oc8051_golden_model_1.n1464 ;
  wire \oc8051_golden_model_1.n1471 ;
  wire [7:0] \oc8051_golden_model_1.n1472 ;
  wire [6:0] \oc8051_golden_model_1.n1473 ;
  wire [7:0] \oc8051_golden_model_1.n1474 ;
  wire [8:0] \oc8051_golden_model_1.n1476 ;
  wire [8:0] \oc8051_golden_model_1.n1478 ;
  wire \oc8051_golden_model_1.n1479 ;
  wire [4:0] \oc8051_golden_model_1.n1480 ;
  wire [4:0] \oc8051_golden_model_1.n1482 ;
  wire \oc8051_golden_model_1.n1483 ;
  wire [8:0] \oc8051_golden_model_1.n1484 ;
  wire \oc8051_golden_model_1.n1491 ;
  wire [7:0] \oc8051_golden_model_1.n1492 ;
  wire [6:0] \oc8051_golden_model_1.n1493 ;
  wire \oc8051_golden_model_1.n1508 ;
  wire [7:0] \oc8051_golden_model_1.n1509 ;
  wire [4:0] \oc8051_golden_model_1.n1511 ;
  wire \oc8051_golden_model_1.n1512 ;
  wire [7:0] \oc8051_golden_model_1.n1513 ;
  wire [6:0] \oc8051_golden_model_1.n1514 ;
  wire [7:0] \oc8051_golden_model_1.n1515 ;
  wire [8:0] \oc8051_golden_model_1.n1517 ;
  wire \oc8051_golden_model_1.n1518 ;
  wire \oc8051_golden_model_1.n1525 ;
  wire [7:0] \oc8051_golden_model_1.n1526 ;
  wire [6:0] \oc8051_golden_model_1.n1527 ;
  wire [7:0] \oc8051_golden_model_1.n1528 ;
  wire [8:0] \oc8051_golden_model_1.n1531 ;
  wire [8:0] \oc8051_golden_model_1.n1532 ;
  wire [7:0] \oc8051_golden_model_1.n1533 ;
  wire [7:0] \oc8051_golden_model_1.n1534 ;
  wire [6:0] \oc8051_golden_model_1.n1535 ;
  wire \oc8051_golden_model_1.n1536 ;
  wire \oc8051_golden_model_1.n1537 ;
  wire \oc8051_golden_model_1.n1538 ;
  wire \oc8051_golden_model_1.n1539 ;
  wire \oc8051_golden_model_1.n1540 ;
  wire \oc8051_golden_model_1.n1541 ;
  wire \oc8051_golden_model_1.n1542 ;
  wire \oc8051_golden_model_1.n1543 ;
  wire \oc8051_golden_model_1.n1550 ;
  wire [7:0] \oc8051_golden_model_1.n1551 ;
  wire [7:0] \oc8051_golden_model_1.n1552 ;
  wire [8:0] \oc8051_golden_model_1.n1555 ;
  wire [8:0] \oc8051_golden_model_1.n1557 ;
  wire \oc8051_golden_model_1.n1558 ;
  wire [4:0] \oc8051_golden_model_1.n1559 ;
  wire [4:0] \oc8051_golden_model_1.n1561 ;
  wire \oc8051_golden_model_1.n1562 ;
  wire \oc8051_golden_model_1.n1569 ;
  wire [7:0] \oc8051_golden_model_1.n1570 ;
  wire [6:0] \oc8051_golden_model_1.n1571 ;
  wire \oc8051_golden_model_1.n1586 ;
  wire [7:0] \oc8051_golden_model_1.n1587 ;
  wire [8:0] \oc8051_golden_model_1.n1591 ;
  wire \oc8051_golden_model_1.n1592 ;
  wire [4:0] \oc8051_golden_model_1.n1594 ;
  wire \oc8051_golden_model_1.n1595 ;
  wire \oc8051_golden_model_1.n1602 ;
  wire [7:0] \oc8051_golden_model_1.n1603 ;
  wire [6:0] \oc8051_golden_model_1.n1604 ;
  wire \oc8051_golden_model_1.n1619 ;
  wire [7:0] \oc8051_golden_model_1.n1620 ;
  wire [8:0] \oc8051_golden_model_1.n1624 ;
  wire \oc8051_golden_model_1.n1625 ;
  wire [4:0] \oc8051_golden_model_1.n1627 ;
  wire \oc8051_golden_model_1.n1628 ;
  wire \oc8051_golden_model_1.n1635 ;
  wire [7:0] \oc8051_golden_model_1.n1636 ;
  wire [6:0] \oc8051_golden_model_1.n1637 ;
  wire \oc8051_golden_model_1.n1652 ;
  wire [7:0] \oc8051_golden_model_1.n1653 ;
  wire [8:0] \oc8051_golden_model_1.n1657 ;
  wire \oc8051_golden_model_1.n1658 ;
  wire [4:0] \oc8051_golden_model_1.n1660 ;
  wire \oc8051_golden_model_1.n1661 ;
  wire \oc8051_golden_model_1.n1668 ;
  wire [7:0] \oc8051_golden_model_1.n1669 ;
  wire [6:0] \oc8051_golden_model_1.n1670 ;
  wire \oc8051_golden_model_1.n1685 ;
  wire [7:0] \oc8051_golden_model_1.n1686 ;
  wire [7:0] \oc8051_golden_model_1.n1700 ;
  wire [6:0] \oc8051_golden_model_1.n1701 ;
  wire [7:0] \oc8051_golden_model_1.n1702 ;
  wire \oc8051_golden_model_1.n1746 ;
  wire [7:0] \oc8051_golden_model_1.n1747 ;
  wire \oc8051_golden_model_1.n1763 ;
  wire [7:0] \oc8051_golden_model_1.n1764 ;
  wire \oc8051_golden_model_1.n1780 ;
  wire [7:0] \oc8051_golden_model_1.n1781 ;
  wire \oc8051_golden_model_1.n1797 ;
  wire [7:0] \oc8051_golden_model_1.n1798 ;
  wire [7:0] \oc8051_golden_model_1.n1810 ;
  wire [6:0] \oc8051_golden_model_1.n1811 ;
  wire [7:0] \oc8051_golden_model_1.n1812 ;
  wire \oc8051_golden_model_1.n1856 ;
  wire [7:0] \oc8051_golden_model_1.n1857 ;
  wire \oc8051_golden_model_1.n1873 ;
  wire [7:0] \oc8051_golden_model_1.n1874 ;
  wire \oc8051_golden_model_1.n1890 ;
  wire [7:0] \oc8051_golden_model_1.n1891 ;
  wire \oc8051_golden_model_1.n1907 ;
  wire [7:0] \oc8051_golden_model_1.n1908 ;
  wire \oc8051_golden_model_1.n1983 ;
  wire [7:0] \oc8051_golden_model_1.n1984 ;
  wire \oc8051_golden_model_1.n2000 ;
  wire [7:0] \oc8051_golden_model_1.n2001 ;
  wire \oc8051_golden_model_1.n2017 ;
  wire [7:0] \oc8051_golden_model_1.n2018 ;
  wire \oc8051_golden_model_1.n2034 ;
  wire [7:0] \oc8051_golden_model_1.n2035 ;
  wire \oc8051_golden_model_1.n2039 ;
  wire [6:0] \oc8051_golden_model_1.n2040 ;
  wire [7:0] \oc8051_golden_model_1.n2041 ;
  wire [6:0] \oc8051_golden_model_1.n2042 ;
  wire [7:0] \oc8051_golden_model_1.n2043 ;
  wire \oc8051_golden_model_1.n2058 ;
  wire [7:0] \oc8051_golden_model_1.n2059 ;
  wire \oc8051_golden_model_1.n2087 ;
  wire [7:0] \oc8051_golden_model_1.n2088 ;
  wire [6:0] \oc8051_golden_model_1.n2089 ;
  wire [7:0] \oc8051_golden_model_1.n2090 ;
  wire [3:0] \oc8051_golden_model_1.n2097 ;
  wire \oc8051_golden_model_1.n2098 ;
  wire [7:0] \oc8051_golden_model_1.n2099 ;
  wire [6:0] \oc8051_golden_model_1.n2100 ;
  wire \oc8051_golden_model_1.n2115 ;
  wire [7:0] \oc8051_golden_model_1.n2116 ;
  wire [7:0] \oc8051_golden_model_1.n2273 ;
  wire \oc8051_golden_model_1.n2276 ;
  wire \oc8051_golden_model_1.n2278 ;
  wire \oc8051_golden_model_1.n2284 ;
  wire [7:0] \oc8051_golden_model_1.n2285 ;
  wire [6:0] \oc8051_golden_model_1.n2286 ;
  wire \oc8051_golden_model_1.n2301 ;
  wire [7:0] \oc8051_golden_model_1.n2302 ;
  wire \oc8051_golden_model_1.n2306 ;
  wire \oc8051_golden_model_1.n2308 ;
  wire \oc8051_golden_model_1.n2314 ;
  wire [7:0] \oc8051_golden_model_1.n2315 ;
  wire [6:0] \oc8051_golden_model_1.n2316 ;
  wire \oc8051_golden_model_1.n2331 ;
  wire [7:0] \oc8051_golden_model_1.n2332 ;
  wire \oc8051_golden_model_1.n2336 ;
  wire \oc8051_golden_model_1.n2338 ;
  wire \oc8051_golden_model_1.n2344 ;
  wire [7:0] \oc8051_golden_model_1.n2345 ;
  wire [6:0] \oc8051_golden_model_1.n2346 ;
  wire \oc8051_golden_model_1.n2361 ;
  wire [7:0] \oc8051_golden_model_1.n2362 ;
  wire \oc8051_golden_model_1.n2366 ;
  wire \oc8051_golden_model_1.n2368 ;
  wire \oc8051_golden_model_1.n2374 ;
  wire [7:0] \oc8051_golden_model_1.n2375 ;
  wire [6:0] \oc8051_golden_model_1.n2376 ;
  wire \oc8051_golden_model_1.n2391 ;
  wire [7:0] \oc8051_golden_model_1.n2392 ;
  wire \oc8051_golden_model_1.n2394 ;
  wire [7:0] \oc8051_golden_model_1.n2395 ;
  wire [6:0] \oc8051_golden_model_1.n2396 ;
  wire [7:0] \oc8051_golden_model_1.n2397 ;
  wire [7:0] \oc8051_golden_model_1.n2398 ;
  wire [6:0] \oc8051_golden_model_1.n2399 ;
  wire [7:0] \oc8051_golden_model_1.n2400 ;
  wire [15:0] \oc8051_golden_model_1.n2404 ;
  wire \oc8051_golden_model_1.n2410 ;
  wire [7:0] \oc8051_golden_model_1.n2411 ;
  wire [6:0] \oc8051_golden_model_1.n2412 ;
  wire \oc8051_golden_model_1.n2427 ;
  wire [7:0] \oc8051_golden_model_1.n2428 ;
  wire \oc8051_golden_model_1.n2430 ;
  wire [7:0] \oc8051_golden_model_1.n2431 ;
  wire [6:0] \oc8051_golden_model_1.n2432 ;
  wire [7:0] \oc8051_golden_model_1.n2433 ;
  wire \oc8051_golden_model_1.n2461 ;
  wire [7:0] \oc8051_golden_model_1.n2462 ;
  wire [6:0] \oc8051_golden_model_1.n2463 ;
  wire [7:0] \oc8051_golden_model_1.n2464 ;
  wire \oc8051_golden_model_1.n2469 ;
  wire [7:0] \oc8051_golden_model_1.n2470 ;
  wire [6:0] \oc8051_golden_model_1.n2471 ;
  wire [7:0] \oc8051_golden_model_1.n2472 ;
  wire \oc8051_golden_model_1.n2477 ;
  wire [7:0] \oc8051_golden_model_1.n2478 ;
  wire [6:0] \oc8051_golden_model_1.n2479 ;
  wire [7:0] \oc8051_golden_model_1.n2480 ;
  wire \oc8051_golden_model_1.n2485 ;
  wire [7:0] \oc8051_golden_model_1.n2486 ;
  wire [6:0] \oc8051_golden_model_1.n2487 ;
  wire [7:0] \oc8051_golden_model_1.n2488 ;
  wire \oc8051_golden_model_1.n2493 ;
  wire [7:0] \oc8051_golden_model_1.n2494 ;
  wire [6:0] \oc8051_golden_model_1.n2495 ;
  wire [7:0] \oc8051_golden_model_1.n2496 ;
  wire [7:0] \oc8051_golden_model_1.n2517 ;
  wire [6:0] \oc8051_golden_model_1.n2518 ;
  wire [7:0] \oc8051_golden_model_1.n2519 ;
  wire [3:0] \oc8051_golden_model_1.n2520 ;
  wire [7:0] \oc8051_golden_model_1.n2521 ;
  wire \oc8051_golden_model_1.n2522 ;
  wire \oc8051_golden_model_1.n2523 ;
  wire \oc8051_golden_model_1.n2524 ;
  wire \oc8051_golden_model_1.n2525 ;
  wire \oc8051_golden_model_1.n2526 ;
  wire \oc8051_golden_model_1.n2527 ;
  wire \oc8051_golden_model_1.n2528 ;
  wire \oc8051_golden_model_1.n2529 ;
  wire \oc8051_golden_model_1.n2536 ;
  wire [7:0] \oc8051_golden_model_1.n2537 ;
  wire [7:0] \oc8051_golden_model_1.n2546 ;
  wire [6:0] \oc8051_golden_model_1.n2547 ;
  wire \oc8051_golden_model_1.n2562 ;
  wire [7:0] \oc8051_golden_model_1.n2563 ;
  wire \oc8051_golden_model_1.n2564 ;
  wire \oc8051_golden_model_1.n2565 ;
  wire \oc8051_golden_model_1.n2566 ;
  wire \oc8051_golden_model_1.n2567 ;
  wire \oc8051_golden_model_1.n2568 ;
  wire \oc8051_golden_model_1.n2569 ;
  wire \oc8051_golden_model_1.n2570 ;
  wire \oc8051_golden_model_1.n2571 ;
  wire \oc8051_golden_model_1.n2578 ;
  wire [7:0] \oc8051_golden_model_1.n2579 ;
  wire \oc8051_golden_model_1.n2580 ;
  wire \oc8051_golden_model_1.n2581 ;
  wire \oc8051_golden_model_1.n2582 ;
  wire \oc8051_golden_model_1.n2583 ;
  wire \oc8051_golden_model_1.n2584 ;
  wire \oc8051_golden_model_1.n2585 ;
  wire \oc8051_golden_model_1.n2586 ;
  wire \oc8051_golden_model_1.n2587 ;
  wire \oc8051_golden_model_1.n2594 ;
  wire [7:0] \oc8051_golden_model_1.n2595 ;
  wire [7:0] \oc8051_golden_model_1.n2625 ;
  wire [6:0] \oc8051_golden_model_1.n2626 ;
  wire [7:0] \oc8051_golden_model_1.n2627 ;
  wire \oc8051_golden_model_1.n2646 ;
  wire [7:0] \oc8051_golden_model_1.n2647 ;
  wire [6:0] \oc8051_golden_model_1.n2648 ;
  wire \oc8051_golden_model_1.n2663 ;
  wire [7:0] \oc8051_golden_model_1.n2664 ;
  wire [7:0] \oc8051_golden_model_1.n2668 ;
  wire [3:0] \oc8051_golden_model_1.n2669 ;
  wire [7:0] \oc8051_golden_model_1.n2670 ;
  wire \oc8051_golden_model_1.n2671 ;
  wire \oc8051_golden_model_1.n2672 ;
  wire \oc8051_golden_model_1.n2673 ;
  wire \oc8051_golden_model_1.n2674 ;
  wire \oc8051_golden_model_1.n2675 ;
  wire \oc8051_golden_model_1.n2676 ;
  wire \oc8051_golden_model_1.n2677 ;
  wire \oc8051_golden_model_1.n2678 ;
  wire \oc8051_golden_model_1.n2685 ;
  wire [7:0] \oc8051_golden_model_1.n2686 ;
  wire \oc8051_golden_model_1.n2690 ;
  wire \oc8051_golden_model_1.n2691 ;
  wire \oc8051_golden_model_1.n2692 ;
  wire \oc8051_golden_model_1.n2693 ;
  wire \oc8051_golden_model_1.n2694 ;
  wire \oc8051_golden_model_1.n2695 ;
  wire \oc8051_golden_model_1.n2696 ;
  wire \oc8051_golden_model_1.n2697 ;
  wire \oc8051_golden_model_1.n2704 ;
  wire [7:0] \oc8051_golden_model_1.n2705 ;
  wire [15:0] \oc8051_golden_model_1.n2706 ;
  wire \oc8051_golden_model_1.n2721 ;
  wire [7:0] \oc8051_golden_model_1.n2722 ;
  wire [7:0] \oc8051_golden_model_1.n2723 ;
  wire \oc8051_golden_model_1.n2739 ;
  wire [7:0] \oc8051_golden_model_1.n2740 ;
  wire [7:0] \oc8051_golden_model_1.n2741 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [7:0] \oc8051_top_1.b_reg ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [15:0] \oc8051_top_1.dptr ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw_next ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  wire [7:0] p0in_reg;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  wire [7:0] p1in_reg;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  wire [7:0] p2in_reg;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [7:0] p3in_reg;
  wire [15:0] pc_impl;
  output property_invalid_acc;
  output property_invalid_b_reg;
  output property_invalid_dec_rom_pc;
  output property_invalid_dph;
  output property_invalid_dpl;
  output property_invalid_iram;
  output property_invalid_p0;
  output property_invalid_p1;
  output property_invalid_p2;
  output property_invalid_p3;
  output property_invalid_pc;
  output property_invalid_psw;
  wire property_invalid_psw_1_r;
  output property_invalid_rom_pc;
  output property_invalid_sp;
  wire property_invalid_sp_1_r;
  wire [7:0] psw_impl;
  wire [15:0] rd_rom_0_addr;
  input rst;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not (_35583_, rst);
  not (_15082_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not (_15093_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_15104_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _15093_);
  and (_15115_, _15104_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_15126_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _15093_);
  and (_15137_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _15093_);
  nor (_15148_, _15137_, _15126_);
  and (_15159_, _15148_, _15115_);
  nor (_15170_, _15159_, _15082_);
  and (_15181_, _15082_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_15192_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and (_15203_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _15192_);
  nor (_15214_, _15203_, _15181_);
  not (_15225_, _15214_);
  and (_15236_, _15225_, _15159_);
  or (_15247_, _15236_, _15170_);
  and (_35774_[1], _15247_, _35583_);
  nor (_15268_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not (_15279_, _15268_);
  and (_15290_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and (_15301_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_15312_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_15322_, _15312_);
  not (_15333_, _15203_);
  nor (_15344_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not (_15355_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_15366_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _15355_);
  nor (_15377_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not (_15388_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_15399_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _15388_);
  nor (_15409_, _15399_, _15377_);
  nor (_15420_, _15409_, _15366_);
  not (_15431_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_15442_, _15366_, _15431_);
  nor (_15453_, _15442_, _15420_);
  and (_15464_, _15453_, _15344_);
  not (_15475_, _15464_);
  and (_15486_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_15496_, _15486_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not (_15507_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_15518_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _15507_);
  and (_15529_, _15518_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_15540_, _15529_, _15496_);
  and (_15551_, _15540_, _15475_);
  nor (_15562_, _15551_, _15333_);
  not (_15573_, _15181_);
  nor (_15584_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor (_15594_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _15388_);
  nor (_15605_, _15594_, _15584_);
  nor (_15616_, _15605_, _15366_);
  not (_15627_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_15638_, _15366_, _15627_);
  nor (_15649_, _15638_, _15616_);
  and (_15660_, _15649_, _15344_);
  not (_15671_, _15660_);
  and (_15681_, _15486_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_15692_, _15518_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_15703_, _15692_, _15681_);
  and (_15714_, _15703_, _15671_);
  nor (_15725_, _15714_, _15573_);
  nor (_15736_, _15725_, _15562_);
  nor (_15747_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor (_15758_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _15388_);
  nor (_15769_, _15758_, _15747_);
  nor (_15779_, _15769_, _15366_);
  not (_15790_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_15801_, _15366_, _15790_);
  nor (_15812_, _15801_, _15779_);
  and (_15823_, _15812_, _15344_);
  not (_15834_, _15823_);
  and (_15845_, _15486_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_15856_, _15518_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_15866_, _15856_, _15845_);
  and (_15877_, _15866_, _15834_);
  nor (_15888_, _15877_, _15225_);
  nor (_15899_, _15888_, _15268_);
  and (_15910_, _15899_, _15736_);
  nor (_15921_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor (_15932_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _15388_);
  nor (_15943_, _15932_, _15921_);
  nor (_15953_, _15943_, _15366_);
  not (_15964_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_15975_, _15366_, _15964_);
  nor (_15986_, _15975_, _15953_);
  and (_15997_, _15986_, _15344_);
  not (_16008_, _15997_);
  and (_16019_, _15486_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_16030_, _15518_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_16041_, _16030_, _16019_);
  and (_16051_, _16041_, _16008_);
  and (_16062_, _16051_, _15268_);
  nor (_16073_, _16062_, _15910_);
  not (_16084_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_16095_, _16084_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16106_, _16095_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16117_, _16106_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_16128_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16138_, _16128_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16149_, _16138_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_16160_, _16149_, _16117_);
  nor (_16171_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16182_, _16171_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_16193_, _16182_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_16204_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16215_, _16095_, _16204_);
  and (_16226_, _16215_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor (_16236_, _16226_, _16193_);
  and (_16247_, _16236_, _16160_);
  and (_16258_, _16128_, _16204_);
  and (_16269_, _16258_, _15986_);
  and (_16280_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_16291_, _16280_, _16204_);
  and (_16302_, _16291_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_16313_, _16280_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_16323_, _16313_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor (_16334_, _16323_, _16302_);
  not (_16345_, _16334_);
  nor (_16356_, _16345_, _16269_);
  and (_16367_, _16356_, _16247_);
  not (_16388_, _16367_);
  and (_16389_, _16388_, _16073_);
  not (_16400_, _16389_);
  nor (_16411_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor (_16421_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _15388_);
  nor (_16432_, _16421_, _16411_);
  nor (_16443_, _16432_, _15366_);
  not (_16454_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_16465_, _15366_, _16454_);
  nor (_16476_, _16465_, _16443_);
  and (_16487_, _16476_, _15344_);
  not (_16498_, _16487_);
  and (_16508_, _15486_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and (_16519_, _15518_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_16530_, _16519_, _16508_);
  and (_16541_, _16530_, _16498_);
  nor (_16552_, _16541_, _15333_);
  nor (_16563_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor (_16574_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _15388_);
  nor (_16585_, _16574_, _16563_);
  nor (_16596_, _16585_, _15366_);
  not (_16597_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_16603_, _15366_, _16597_);
  nor (_16614_, _16603_, _16596_);
  and (_16625_, _16614_, _15344_);
  not (_16636_, _16625_);
  and (_16647_, _15486_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_16658_, _15518_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_16669_, _16658_, _16647_);
  and (_16680_, _16669_, _16636_);
  nor (_16691_, _16680_, _15573_);
  nor (_16702_, _16691_, _16552_);
  nor (_16712_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor (_16723_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _15388_);
  nor (_16734_, _16723_, _16712_);
  nor (_16745_, _16734_, _15366_);
  not (_16756_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_16767_, _15366_, _16756_);
  nor (_16778_, _16767_, _16745_);
  and (_16789_, _16778_, _15344_);
  not (_16800_, _16789_);
  and (_16811_, _15486_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and (_16821_, _15518_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_16832_, _16821_, _16811_);
  and (_16843_, _16832_, _16800_);
  nor (_16854_, _16843_, _15225_);
  nor (_16865_, _16854_, _15268_);
  and (_16876_, _16865_, _16702_);
  nor (_16887_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_16898_, _15388_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_16909_, _16898_, _16887_);
  nor (_16920_, _16909_, _15366_);
  not (_16930_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_16941_, _15366_, _16930_);
  nor (_16952_, _16941_, _16920_);
  and (_16963_, _16952_, _15344_);
  not (_16974_, _16963_);
  and (_16985_, _15486_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_16996_, _15518_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_17007_, _16996_, _16985_);
  and (_17018_, _17007_, _16974_);
  and (_17029_, _17018_, _15268_);
  nor (_17039_, _17029_, _16876_);
  and (_17050_, _16138_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_17061_, _16106_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_17072_, _17061_, _17050_);
  and (_17093_, _16291_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_17094_, _16182_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_17115_, _17094_, _17093_);
  and (_17116_, _17115_, _17072_);
  and (_17127_, _16952_, _16258_);
  and (_17138_, _16215_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_17148_, _16313_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_17159_, _17148_, _17138_);
  not (_17170_, _17159_);
  nor (_17181_, _17170_, _17127_);
  and (_17192_, _17181_, _17116_);
  not (_17203_, _17192_);
  and (_17214_, _17203_, _17039_);
  and (_17225_, _17214_, _16400_);
  not (_17236_, _17225_);
  and (_17247_, _16106_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_17257_, _16138_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_17268_, _17257_, _17247_);
  and (_17279_, _16182_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and (_17290_, _16215_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_17301_, _17290_, _17279_);
  and (_17312_, _17301_, _17268_);
  and (_17323_, _16614_, _16258_);
  and (_17334_, _16313_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_17345_, _16291_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_17356_, _17345_, _17334_);
  not (_17366_, _17356_);
  nor (_17377_, _17366_, _17323_);
  and (_17388_, _17377_, _17312_);
  not (_17399_, _17388_);
  and (_17410_, _17399_, _17039_);
  and (_17421_, _16106_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_17432_, _16138_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_17443_, _17432_, _17421_);
  and (_17454_, _16215_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_17465_, _16182_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor (_17475_, _17465_, _17454_);
  and (_17486_, _17475_, _17443_);
  and (_17497_, _16258_, _15649_);
  and (_17508_, _16291_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_17519_, _16313_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_17530_, _17519_, _17508_);
  not (_17541_, _17530_);
  nor (_17552_, _17541_, _17497_);
  and (_17563_, _17552_, _17486_);
  not (_17574_, _17563_);
  and (_17584_, _17574_, _16073_);
  and (_17595_, _17410_, _17584_);
  and (_17606_, _16388_, _17595_);
  nor (_17617_, _16389_, _17595_);
  nor (_17628_, _17617_, _17606_);
  and (_17639_, _17628_, _17410_);
  and (_17650_, _17214_, _16389_);
  and (_17661_, _16388_, _17039_);
  and (_17672_, _17203_, _16073_);
  nor (_17683_, _17672_, _17661_);
  nor (_17693_, _17683_, _17650_);
  and (_17704_, _17693_, _17639_);
  nor (_17715_, _17693_, _17639_);
  nor (_17726_, _17715_, _17704_);
  and (_17737_, _17726_, _17606_);
  nor (_17748_, _17737_, _17704_);
  nor (_17759_, _17748_, _17236_);
  and (_17770_, _17039_, _17574_);
  and (_17781_, _16106_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_17792_, _16138_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_17802_, _17792_, _17781_);
  and (_17813_, _16182_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_17824_, _16215_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor (_17835_, _17824_, _17813_);
  and (_17846_, _17835_, _17802_);
  and (_17857_, _16476_, _16258_);
  and (_17868_, _16291_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_17879_, _16313_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor (_17890_, _17879_, _17868_);
  not (_17901_, _17890_);
  nor (_17911_, _17901_, _17857_);
  and (_17922_, _17911_, _17846_);
  not (_17933_, _17922_);
  and (_17944_, _17933_, _16073_);
  and (_17955_, _17944_, _17770_);
  and (_17966_, _17399_, _16073_);
  nor (_17977_, _17966_, _17770_);
  nor (_17988_, _17977_, _17595_);
  and (_17999_, _17988_, _17955_);
  nor (_18010_, _16389_, _17410_);
  nor (_18020_, _18010_, _17639_);
  and (_18031_, _18020_, _17999_);
  nor (_18042_, _17726_, _17606_);
  nor (_18053_, _18042_, _17737_);
  and (_18064_, _18053_, _18031_);
  nor (_18075_, _18053_, _18031_);
  nor (_18086_, _18075_, _18064_);
  not (_18097_, _18086_);
  and (_18108_, _16106_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_18119_, _16138_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_18129_, _18119_, _18108_);
  and (_18140_, _16182_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and (_18151_, _16215_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor (_18162_, _18151_, _18140_);
  and (_18173_, _18162_, _18129_);
  and (_18184_, _16778_, _16258_);
  and (_18195_, _16313_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and (_18206_, _16291_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_18217_, _18206_, _18195_);
  not (_18227_, _18217_);
  nor (_18238_, _18227_, _18184_);
  and (_18249_, _18238_, _18173_);
  not (_18260_, _18249_);
  and (_18271_, _18260_, _17039_);
  and (_18282_, _16106_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_18293_, _16138_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_18304_, _18293_, _18282_);
  and (_18315_, _16182_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and (_18326_, _16215_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor (_18336_, _18326_, _18315_);
  and (_18347_, _18336_, _18304_);
  and (_18358_, _16258_, _15453_);
  and (_18369_, _16291_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_18380_, _16313_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor (_18391_, _18380_, _18369_);
  not (_18402_, _18391_);
  nor (_18413_, _18402_, _18358_);
  and (_18424_, _18413_, _18347_);
  not (_18435_, _18424_);
  and (_18445_, _18435_, _16073_);
  and (_18456_, _18445_, _18271_);
  and (_18467_, _18260_, _16073_);
  not (_18478_, _18467_);
  and (_18489_, _18435_, _17039_);
  and (_18500_, _18489_, _18478_);
  and (_18511_, _18500_, _17944_);
  nor (_18522_, _18511_, _18456_);
  and (_18533_, _17933_, _17039_);
  nor (_18544_, _18533_, _17584_);
  nor (_18554_, _18544_, _17955_);
  not (_18565_, _18554_);
  nor (_18576_, _18565_, _18522_);
  nor (_18587_, _17988_, _17955_);
  nor (_18598_, _18587_, _17999_);
  and (_18609_, _18598_, _18576_);
  nor (_18620_, _18020_, _17999_);
  nor (_18631_, _18620_, _18031_);
  and (_18642_, _18631_, _18609_);
  and (_18653_, _16106_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_18663_, _16138_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_18674_, _18663_, _18653_);
  and (_18685_, _16215_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and (_18696_, _16182_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor (_18707_, _18696_, _18685_);
  and (_18718_, _18707_, _18674_);
  and (_18729_, _16258_, _15812_);
  and (_18740_, _16291_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_18751_, _16313_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_18762_, _18751_, _18740_);
  not (_18772_, _18762_);
  nor (_18783_, _18772_, _18729_);
  and (_18794_, _18783_, _18718_);
  not (_18805_, _18794_);
  and (_18816_, _18805_, _17039_);
  and (_18827_, _18816_, _18467_);
  nor (_18838_, _18445_, _18271_);
  nor (_18849_, _18838_, _18456_);
  and (_18860_, _18849_, _18827_);
  nor (_18871_, _18500_, _17944_);
  nor (_18881_, _18871_, _18511_);
  and (_18892_, _18881_, _18860_);
  and (_18903_, _18565_, _18522_);
  nor (_18914_, _18903_, _18576_);
  and (_18925_, _18914_, _18892_);
  nor (_18936_, _18598_, _18576_);
  nor (_18947_, _18936_, _18609_);
  and (_18958_, _18947_, _18925_);
  nor (_18969_, _18631_, _18609_);
  nor (_18980_, _18969_, _18642_);
  and (_18990_, _18980_, _18958_);
  nor (_19001_, _18990_, _18642_);
  nor (_19012_, _19001_, _18097_);
  nor (_19023_, _19012_, _18064_);
  and (_19034_, _17748_, _17236_);
  nor (_19045_, _19034_, _17759_);
  not (_19056_, _19045_);
  nor (_19067_, _19056_, _19023_);
  or (_19078_, _19067_, _17650_);
  nor (_19089_, _19078_, _17759_);
  nor (_19099_, _19089_, _15322_);
  and (_19110_, _19089_, _15322_);
  nor (_19121_, _19110_, _19099_);
  not (_19132_, _19121_);
  and (_19143_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_19154_, _19056_, _19023_);
  nor (_19165_, _19154_, _19067_);
  and (_19176_, _19165_, _19143_);
  and (_19187_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and (_19198_, _19001_, _18097_);
  nor (_19208_, _19198_, _19012_);
  and (_19219_, _19208_, _19187_);
  nor (_19230_, _19208_, _19187_);
  nor (_19241_, _19230_, _19219_);
  not (_19252_, _19241_);
  and (_19263_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor (_19274_, _18980_, _18958_);
  nor (_19285_, _19274_, _18990_);
  and (_19296_, _19285_, _19263_);
  nor (_19307_, _19285_, _19263_);
  nor (_19317_, _19307_, _19296_);
  not (_19328_, _19317_);
  and (_19339_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor (_19350_, _18947_, _18925_);
  nor (_19361_, _19350_, _18958_);
  and (_19372_, _19361_, _19339_);
  nor (_19383_, _19361_, _19339_);
  nor (_19394_, _19383_, _19372_);
  not (_19405_, _19394_);
  and (_19416_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor (_19426_, _18914_, _18892_);
  nor (_19437_, _19426_, _18925_);
  and (_19448_, _19437_, _19416_);
  and (_19459_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor (_19470_, _18881_, _18860_);
  nor (_19481_, _19470_, _18892_);
  and (_19492_, _19481_, _19459_);
  and (_19503_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor (_19514_, _18849_, _18827_);
  nor (_19524_, _19514_, _18860_);
  and (_19535_, _19524_, _19503_);
  nor (_19546_, _19481_, _19459_);
  nor (_19557_, _19546_, _19492_);
  and (_19568_, _19557_, _19535_);
  nor (_19579_, _19568_, _19492_);
  not (_19590_, _19579_);
  nor (_19601_, _19437_, _19416_);
  nor (_19612_, _19601_, _19448_);
  and (_19623_, _19612_, _19590_);
  nor (_19633_, _19623_, _19448_);
  nor (_19644_, _19633_, _19405_);
  nor (_19655_, _19644_, _19372_);
  nor (_19666_, _19655_, _19328_);
  nor (_19677_, _19666_, _19296_);
  nor (_19688_, _19677_, _19252_);
  nor (_19699_, _19688_, _19219_);
  nor (_19710_, _19165_, _19143_);
  nor (_19721_, _19710_, _19176_);
  not (_19732_, _19721_);
  nor (_19743_, _19732_, _19699_);
  nor (_19754_, _19743_, _19176_);
  nor (_19765_, _19754_, _19132_);
  nor (_19776_, _19765_, _19099_);
  not (_19787_, _19776_);
  and (_19798_, _19787_, _15301_);
  and (_19809_, _19798_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_19820_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_19831_, _19820_, _19809_);
  and (_19842_, _19831_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_19853_, _19842_, _15290_);
  and (_19864_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_19875_, _19864_, _19853_);
  and (_19886_, _19853_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor (_19897_, _19886_, _19875_);
  and (_35775_[15], _19897_, _35583_);
  nor (_19917_, _15159_, _15192_);
  and (_19928_, _15159_, _15192_);
  or (_19939_, _19928_, _19917_);
  and (_35774_[0], _19939_, _35583_);
  and (_19960_, _18805_, _16073_);
  and (_35775_[0], _19960_, _35583_);
  nor (_19981_, _18816_, _18467_);
  nor (_19992_, _19981_, _18827_);
  and (_35775_[1], _19992_, _35583_);
  nor (_20013_, _19524_, _19503_);
  nor (_20024_, _20013_, _19535_);
  and (_35775_[2], _20024_, _35583_);
  nor (_20045_, _19557_, _19535_);
  nor (_20056_, _20045_, _19568_);
  and (_35775_[3], _20056_, _35583_);
  nor (_20077_, _19612_, _19590_);
  nor (_20088_, _20077_, _19623_);
  and (_35775_[4], _20088_, _35583_);
  and (_20109_, _19633_, _19405_);
  nor (_20120_, _20109_, _19644_);
  and (_35775_[5], _20120_, _35583_);
  and (_20141_, _19655_, _19328_);
  nor (_20152_, _20141_, _19666_);
  and (_35775_[6], _20152_, _35583_);
  and (_20173_, _19677_, _19252_);
  nor (_20184_, _20173_, _19688_);
  and (_35775_[7], _20184_, _35583_);
  and (_20205_, _19732_, _19699_);
  nor (_20216_, _20205_, _19743_);
  and (_35775_[8], _20216_, _35583_);
  and (_20237_, _19754_, _19132_);
  nor (_20248_, _20237_, _19765_);
  and (_35775_[9], _20248_, _35583_);
  nor (_20269_, _19787_, _15301_);
  nor (_20280_, _20269_, _19798_);
  and (_35775_[10], _20280_, _35583_);
  and (_20300_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor (_20311_, _20300_, _19798_);
  nor (_20322_, _20311_, _19809_);
  and (_35775_[11], _20322_, _35583_);
  nor (_20343_, _19820_, _19809_);
  nor (_20354_, _20343_, _19831_);
  and (_35775_[12], _20354_, _35583_);
  and (_20375_, _15279_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor (_20386_, _20375_, _19831_);
  nor (_20397_, _20386_, _19842_);
  and (_35775_[13], _20397_, _35583_);
  nor (_20418_, _19842_, _15290_);
  nor (_20429_, _20418_, _19853_);
  and (_35775_[14], _20429_, _35583_);
  and (_20450_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _15093_);
  nor (_20461_, _20450_, _15104_);
  not (_20472_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_20483_, _15126_, _20472_);
  and (_20494_, _20483_, _20461_);
  and (_20505_, _20494_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_20516_, _20505_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_20527_, _20505_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20538_, _20527_, _20516_);
  and (_35771_[1], _20538_, _35583_);
  and (_35772_[5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _35583_);
  not (_20569_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_20580_, _16843_, _20569_);
  and (_20591_, _16541_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20602_, _20591_, _20580_);
  nor (_20613_, _20602_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20624_, _16680_, _20569_);
  and (_20635_, _17018_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_20646_, _20635_, _20624_);
  and (_20657_, _20646_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_20667_, _20657_, _20613_);
  nor (_20678_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20689_, _20678_, _17192_);
  nor (_20700_, _20678_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor (_20711_, _20700_, _20689_);
  not (_20722_, _20711_);
  and (_20733_, _15877_, _20569_);
  and (_20744_, _15551_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20755_, _20744_, _20733_);
  nor (_20766_, _20755_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_20777_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20788_, _15714_, _20569_);
  and (_20799_, _16051_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20810_, _20799_, _20788_);
  nor (_20821_, _20810_, _20777_);
  nor (_20832_, _20821_, _20766_);
  nor (_20843_, _20832_, _20722_);
  and (_20854_, _20832_, _20722_);
  nor (_20865_, _20854_, _20843_);
  nor (_20876_, _20678_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  and (_20887_, _20678_, _16367_);
  nor (_20898_, _20887_, _20876_);
  not (_20909_, _20898_);
  nor (_20920_, _16843_, _20569_);
  nor (_20931_, _20920_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_20942_, _16541_, _20569_);
  and (_20953_, _16680_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_20964_, _20953_, _20942_);
  nor (_20975_, _20964_, _20777_);
  nor (_20986_, _20975_, _20931_);
  nor (_20997_, _20986_, _20909_);
  and (_21008_, _20986_, _20909_);
  nor (_21019_, _21008_, _20997_);
  not (_21030_, _21019_);
  nor (_21040_, _20678_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  and (_21051_, _20678_, _17388_);
  nor (_21062_, _21051_, _21040_);
  not (_21073_, _21062_);
  nor (_21084_, _15877_, _20569_);
  nor (_21095_, _21084_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21106_, _15551_, _20569_);
  and (_21117_, _15714_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_21128_, _21117_, _21106_);
  nor (_21139_, _21128_, _20777_);
  nor (_21150_, _21139_, _21095_);
  nor (_21161_, _21150_, _21073_);
  and (_21172_, _21150_, _21073_);
  and (_21183_, _20602_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21194_, _21183_);
  nor (_21205_, _20678_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and (_21216_, _20678_, _17563_);
  nor (_21227_, _21216_, _21205_);
  and (_21238_, _21227_, _21194_);
  and (_21249_, _20755_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21260_, _21249_);
  and (_21271_, _20678_, _17922_);
  nor (_21282_, _20678_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor (_21293_, _21282_, _21271_);
  and (_21314_, _21293_, _21260_);
  nor (_21325_, _21293_, _21260_);
  nor (_21336_, _21325_, _21314_);
  not (_21347_, _21336_);
  and (_21358_, _20920_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21369_, _21358_);
  and (_21370_, _20678_, _18424_);
  nor (_21381_, _20678_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor (_21392_, _21381_, _21370_);
  and (_21402_, _21392_, _21369_);
  and (_21413_, _21084_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_21424_, _21413_);
  nor (_21435_, _20678_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and (_21446_, _20678_, _18249_);
  nor (_21457_, _21446_, _21435_);
  nor (_21468_, _21457_, _21424_);
  not (_21479_, _21468_);
  nor (_21490_, _21392_, _21369_);
  nor (_21501_, _21490_, _21402_);
  and (_21512_, _21501_, _21479_);
  nor (_21523_, _21512_, _21402_);
  nor (_21534_, _21523_, _21347_);
  nor (_21545_, _21534_, _21314_);
  nor (_21556_, _21227_, _21194_);
  nor (_21567_, _21556_, _21238_);
  not (_21578_, _21567_);
  nor (_21589_, _21578_, _21545_);
  nor (_21600_, _21589_, _21238_);
  nor (_21611_, _21600_, _21172_);
  nor (_21622_, _21611_, _21161_);
  nor (_21633_, _21622_, _21030_);
  nor (_21644_, _21633_, _20997_);
  not (_21655_, _21644_);
  and (_21666_, _21655_, _20865_);
  or (_21677_, _21666_, _20843_);
  and (_21688_, _17018_, _16051_);
  or (_21699_, _21688_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_21710_, _20964_);
  and (_21721_, _20646_, _21710_);
  nor (_21732_, _21128_, _20810_);
  and (_21743_, _21732_, _21721_);
  or (_21754_, _21743_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_21765_, _21754_, _21699_);
  and (_21775_, _21765_, _21677_);
  and (_21786_, _21775_, _20667_);
  nor (_21797_, _21655_, _20865_);
  or (_21808_, _21797_, _21666_);
  and (_21819_, _21808_, _21786_);
  nor (_21830_, _21786_, _20711_);
  nor (_21841_, _21830_, _21819_);
  not (_21852_, _21841_);
  and (_21863_, _21841_, _20667_);
  not (_21884_, _20832_);
  nor (_21885_, _21786_, _20909_);
  and (_21896_, _21622_, _21030_);
  nor (_21907_, _21896_, _21633_);
  and (_21918_, _21907_, _21786_);
  or (_21929_, _21918_, _21885_);
  and (_21940_, _21929_, _21884_);
  nor (_21951_, _21929_, _21884_);
  nor (_21962_, _21951_, _21940_);
  not (_21973_, _21962_);
  not (_21984_, _20986_);
  nor (_21995_, _21786_, _21073_);
  nor (_22006_, _21172_, _21161_);
  nor (_22017_, _22006_, _21600_);
  and (_22028_, _22006_, _21600_);
  or (_22039_, _22028_, _22017_);
  and (_22050_, _22039_, _21786_);
  or (_22061_, _22050_, _21995_);
  and (_22072_, _22061_, _21984_);
  nor (_22083_, _22061_, _21984_);
  nor (_22094_, _22083_, _22072_);
  not (_22105_, _22094_);
  not (_22116_, _21150_);
  and (_22126_, _21578_, _21545_);
  or (_22147_, _22126_, _21589_);
  and (_22148_, _22147_, _21786_);
  nor (_22159_, _21786_, _21227_);
  nor (_22170_, _22159_, _22148_);
  and (_22181_, _22170_, _22116_);
  and (_22192_, _21523_, _21347_);
  nor (_22203_, _22192_, _21534_);
  not (_22214_, _22203_);
  and (_22225_, _22214_, _21786_);
  nor (_22236_, _21786_, _21293_);
  nor (_22247_, _22236_, _22225_);
  and (_22258_, _22247_, _21194_);
  nor (_22269_, _22247_, _21194_);
  nor (_22280_, _22269_, _22258_);
  not (_22291_, _22280_);
  nor (_22302_, _21501_, _21479_);
  nor (_22313_, _22302_, _21512_);
  not (_22324_, _22313_);
  and (_22335_, _22324_, _21786_);
  nor (_22346_, _21786_, _21392_);
  nor (_22357_, _22346_, _22335_);
  and (_22368_, _22357_, _21260_);
  and (_22379_, _21786_, _21413_);
  nor (_22390_, _22379_, _21457_);
  and (_22401_, _22379_, _21457_);
  nor (_22412_, _22401_, _22390_);
  and (_22423_, _22412_, _21369_);
  nor (_22434_, _22412_, _21369_);
  nor (_22445_, _22434_, _22423_);
  and (_22456_, _20678_, _18794_);
  nor (_22467_, _20678_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_22478_, _22467_, _22456_);
  nor (_22489_, _22478_, _21424_);
  not (_22499_, _22489_);
  and (_22510_, _22499_, _22445_);
  nor (_22521_, _22510_, _22423_);
  nor (_22532_, _22357_, _21260_);
  nor (_22543_, _22532_, _22368_);
  not (_22554_, _22543_);
  nor (_22565_, _22554_, _22521_);
  nor (_22576_, _22565_, _22368_);
  nor (_22587_, _22576_, _22291_);
  nor (_22598_, _22587_, _22258_);
  nor (_22609_, _22170_, _22116_);
  nor (_22620_, _22609_, _22181_);
  not (_22631_, _22620_);
  nor (_22642_, _22631_, _22598_);
  nor (_22653_, _22642_, _22181_);
  nor (_22664_, _22653_, _22105_);
  nor (_22675_, _22664_, _22072_);
  nor (_22686_, _22675_, _21973_);
  or (_22697_, _22686_, _21940_);
  or (_22708_, _22697_, _21863_);
  and (_22719_, _22708_, _21765_);
  nor (_22730_, _22719_, _21852_);
  and (_22741_, _21863_, _21765_);
  and (_22752_, _22741_, _22697_);
  or (_22763_, _22752_, _22730_);
  and (_35773_[7], _22763_, _35583_);
  or (_22784_, _21841_, _20667_);
  and (_22795_, _22784_, _22719_);
  and (_35772_[0], _22795_, _35583_);
  and (_35772_[1], _21786_, _35583_);
  and (_35772_[2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _35583_);
  and (_35772_[3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _35583_);
  and (_35772_[4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _35583_);
  or (_22855_, _20494_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_22866_, _20505_, rst);
  and (_35771_[0], _22866_, _22855_);
  and (_22887_, _22795_, _21413_);
  or (_22898_, _22887_, _22478_);
  nand (_22919_, _22887_, _22478_);
  and (_22920_, _22919_, _22898_);
  and (_35773_[0], _22920_, _35583_);
  nor (_22951_, _22499_, _22445_);
  or (_22952_, _22951_, _22510_);
  nand (_22963_, _22952_, _22795_);
  or (_22984_, _22795_, _22412_);
  and (_22985_, _22984_, _22963_);
  and (_35773_[1], _22985_, _35583_);
  and (_23016_, _22554_, _22521_);
  or (_23017_, _23016_, _22565_);
  nand (_23028_, _23017_, _22795_);
  or (_23039_, _22795_, _22357_);
  and (_23050_, _23039_, _23028_);
  and (_35773_[2], _23050_, _35583_);
  and (_23071_, _22576_, _22291_);
  or (_23082_, _23071_, _22587_);
  nand (_23093_, _23082_, _22795_);
  or (_23104_, _22795_, _22247_);
  and (_23115_, _23104_, _23093_);
  and (_35773_[3], _23115_, _35583_);
  and (_23136_, _22631_, _22598_);
  or (_23147_, _23136_, _22642_);
  nand (_23158_, _23147_, _22795_);
  or (_23168_, _22795_, _22170_);
  and (_23179_, _23168_, _23158_);
  and (_35773_[4], _23179_, _35583_);
  and (_23200_, _22653_, _22105_);
  or (_23211_, _23200_, _22664_);
  nand (_23222_, _23211_, _22795_);
  or (_23233_, _22795_, _22061_);
  and (_23244_, _23233_, _23222_);
  and (_35773_[5], _23244_, _35583_);
  and (_23265_, _22675_, _21973_);
  or (_23276_, _23265_, _22686_);
  nand (_23287_, _23276_, _22795_);
  or (_23298_, _22795_, _21929_);
  and (_23309_, _23298_, _23287_);
  and (_35773_[6], _23309_, _35583_);
  and (_23330_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_23341_, _23330_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_23352_, _23341_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_23363_, _23352_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_23374_, _23363_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_23385_, _23374_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_23396_, _23385_);
  not (_23407_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23418_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _15093_);
  and (_23429_, _23418_, _23407_);
  and (_23440_, _23429_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  not (_23451_, _23440_);
  nor (_23462_, _23374_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_23473_, _23462_, _23451_);
  and (_23483_, _23473_, _23396_);
  not (_23494_, _23483_);
  and (_23505_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23516_, _23505_, _23418_);
  not (_23527_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_23538_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _15093_);
  and (_23549_, _23538_, _23527_);
  and (_23560_, _23549_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23571_, _23560_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor (_23582_, _23571_, _23516_);
  not (_23593_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_23604_, _23429_, _23593_);
  and (_23615_, _23604_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_23626_, _23549_, _23407_);
  and (_23637_, _23626_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor (_23648_, _23637_, _23615_);
  and (_23659_, _23648_, _23582_);
  and (_23670_, _23659_, _23494_);
  not (_23681_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_23692_, _23385_, _23681_);
  and (_23703_, _23385_, _23681_);
  nor (_23714_, _23703_, _23692_);
  nor (_23725_, _23714_, _23451_);
  not (_23736_, _23725_);
  and (_23747_, _23626_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_23758_, _23747_, _23516_);
  and (_23769_, _23604_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_23780_, _23560_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor (_23790_, _23780_, _23769_);
  and (_23801_, _23790_, _23758_);
  and (_23812_, _23801_, _23736_);
  nor (_23823_, _23812_, _23670_);
  and (_23834_, _23560_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_23845_, _23626_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_23856_, _23845_, _23834_);
  not (_23867_, _23352_);
  nor (_23878_, _23341_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_23889_, _23878_, _23451_);
  and (_23900_, _23889_, _23867_);
  or (_23911_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_23922_, _23911_, _15093_);
  nor (_23933_, _23922_, _23538_);
  and (_23944_, _23933_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_23955_, _23604_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_23966_, _23955_, _23944_);
  not (_23977_, _23966_);
  nor (_23988_, _23977_, _23900_);
  and (_24009_, _23988_, _23856_);
  not (_24020_, _24009_);
  and (_24031_, _23560_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor (_24042_, _24031_, _23516_);
  nor (_24053_, _23352_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or (_24064_, _24053_, _23451_);
  nor (_24075_, _24064_, _23363_);
  and (_24076_, _23626_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_24087_, _24076_, _24075_);
  and (_24098_, _24087_, _24042_);
  and (_24108_, _23933_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and (_24119_, _23604_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_24130_, _24119_, _24108_);
  and (_24141_, _24130_, _24098_);
  nor (_24152_, _24141_, _24020_);
  nor (_24163_, _23363_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_24174_, _24163_);
  nor (_24185_, _23451_, _23374_);
  and (_24196_, _24185_, _24174_);
  not (_24207_, _24196_);
  and (_24218_, _23626_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor (_24229_, _24218_, _23516_);
  and (_24240_, _23604_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_24251_, _23560_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_24262_, _24251_, _24240_);
  and (_24273_, _24262_, _24229_);
  and (_24284_, _24273_, _24207_);
  not (_24295_, _24284_);
  and (_24306_, _23560_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  and (_24317_, _23626_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_24328_, _24317_, _24306_);
  and (_24339_, _23604_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  not (_24350_, _24339_);
  not (_24361_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_24372_, _23440_, _24361_);
  and (_24383_, _23933_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_24394_, _24383_, _24372_);
  and (_24405_, _24394_, _24350_);
  and (_24416_, _24405_, _24328_);
  nor (_24426_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_24437_, _24426_, _23330_);
  and (_24448_, _24437_, _23440_);
  and (_24459_, _23626_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  nor (_24470_, _24459_, _24448_);
  and (_24481_, _23933_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  not (_24492_, _24481_);
  and (_24503_, _23560_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_24514_, _23604_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_24525_, _24514_, _24503_);
  and (_24536_, _24525_, _24492_);
  and (_24547_, _24536_, _24470_);
  nor (_24558_, _23330_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_24569_, _24558_, _23341_);
  and (_24580_, _24569_, _23440_);
  and (_24591_, _23604_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_24602_, _24591_, _24580_);
  and (_24613_, _23560_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_24624_, _23626_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  and (_24635_, _23933_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_24646_, _24635_, _24624_);
  nor (_24657_, _24646_, _24613_);
  and (_24668_, _24657_, _24602_);
  and (_24679_, _24668_, _24547_);
  and (_24690_, _24679_, _24416_);
  and (_24701_, _24690_, _24295_);
  and (_24712_, _24701_, _24152_);
  nand (_24723_, _24712_, _23823_);
  and (_24733_, _22763_, _20494_);
  not (_24744_, _24733_);
  and (_24755_, _19897_, _15159_);
  not (_24766_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_24777_, _15104_, _24766_);
  and (_24788_, _24777_, _15148_);
  not (_24799_, _24788_);
  nor (_24810_, _17192_, _17018_);
  and (_24821_, _17192_, _17018_);
  nor (_24832_, _24821_, _24810_);
  not (_24843_, _16051_);
  nor (_24854_, _16367_, _24843_);
  nor (_24865_, _16367_, _16051_);
  and (_24876_, _16367_, _16051_);
  nor (_24887_, _24876_, _24865_);
  not (_24898_, _16680_);
  nor (_24909_, _17388_, _24898_);
  nor (_24930_, _17388_, _16680_);
  and (_24931_, _17388_, _16680_);
  nor (_24942_, _24931_, _24930_);
  not (_24953_, _15714_);
  and (_24974_, _17563_, _24953_);
  nor (_24975_, _24974_, _24942_);
  nor (_24986_, _24975_, _24909_);
  nor (_25007_, _24986_, _24887_);
  nor (_25008_, _25007_, _24854_);
  and (_25019_, _24986_, _24887_);
  nor (_25030_, _25019_, _25007_);
  not (_25041_, _25030_);
  and (_25062_, _24974_, _24942_);
  nor (_25063_, _25062_, _24975_);
  not (_25074_, _25063_);
  nor (_25085_, _17563_, _15714_);
  and (_25096_, _17563_, _15714_);
  nor (_25107_, _25096_, _25085_);
  not (_25118_, _25107_);
  and (_25129_, _17922_, _16541_);
  nor (_25140_, _17922_, _16541_);
  nor (_25151_, _25140_, _25129_);
  nor (_25162_, _18424_, _15551_);
  and (_25173_, _18424_, _15551_);
  nor (_25194_, _25173_, _25162_);
  nor (_25195_, _18249_, _16843_);
  and (_25206_, _18249_, _16843_);
  nor (_25217_, _25206_, _25195_);
  not (_25228_, _15877_);
  and (_25239_, _18794_, _25228_);
  nor (_25250_, _25239_, _25217_);
  not (_25261_, _16843_);
  nor (_25272_, _18249_, _25261_);
  nor (_25283_, _25272_, _25250_);
  nor (_25294_, _25283_, _25194_);
  not (_25305_, _15551_);
  nor (_25316_, _18424_, _25305_);
  nor (_25327_, _25316_, _25294_);
  nor (_25338_, _25327_, _25151_);
  and (_25349_, _25327_, _25151_);
  nor (_25370_, _25349_, _25338_);
  not (_25371_, _25370_);
  and (_25382_, _25283_, _25194_);
  nor (_25393_, _25382_, _25294_);
  not (_25404_, _25393_);
  and (_25415_, _25239_, _25217_);
  nor (_25426_, _25415_, _25250_);
  not (_25437_, _25426_);
  nor (_25448_, _18794_, _15877_);
  and (_25459_, _18794_, _15877_);
  nor (_25470_, _25459_, _25448_);
  not (_25481_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and (_25492_, _15366_, _25481_);
  not (_25503_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_25514_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and (_25525_, _25514_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25536_, _25525_, _15943_);
  nor (_25547_, _25536_, _25503_);
  nor (_25568_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25569_, _25568_, _15605_);
  not (_25580_, _25569_);
  and (_25591_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25602_, _25591_, _16909_);
  not (_25613_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and (_25624_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _25613_);
  and (_25635_, _25624_, _16585_);
  nor (_25646_, _25635_, _25602_);
  and (_25657_, _25646_, _25580_);
  and (_25668_, _25657_, _25547_);
  and (_25679_, _25525_, _15409_);
  nor (_25690_, _25679_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_25701_, _25624_, _16734_);
  not (_25712_, _25701_);
  and (_25723_, _25591_, _16432_);
  and (_25734_, _25568_, _15769_);
  nor (_25745_, _25734_, _25723_);
  and (_25756_, _25745_, _25712_);
  and (_25767_, _25756_, _25690_);
  nor (_25778_, _25767_, _25668_);
  nor (_25789_, _25778_, _15366_);
  nor (_25800_, _25789_, _25492_);
  and (_25811_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_25822_, _25811_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_25833_, _25822_);
  and (_25844_, _25833_, _25800_);
  and (_25855_, _25833_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_25866_, _25855_, _25844_);
  nor (_25877_, _25866_, _25470_);
  and (_25888_, _25877_, _25437_);
  and (_25899_, _25888_, _25404_);
  and (_25920_, _25899_, _25371_);
  not (_25921_, _16541_);
  or (_25932_, _17922_, _25921_);
  and (_25943_, _17922_, _25921_);
  or (_25954_, _25327_, _25943_);
  and (_25965_, _25954_, _25932_);
  or (_25976_, _25965_, _25920_);
  and (_25987_, _25976_, _25118_);
  and (_25998_, _25987_, _25074_);
  and (_26009_, _25998_, _25041_);
  nor (_26030_, _26009_, _25008_);
  nor (_26031_, _26030_, _24832_);
  and (_26042_, _26030_, _24832_);
  nor (_26053_, _26042_, _26031_);
  nor (_26064_, _26053_, _24799_);
  not (_26075_, _26064_);
  not (_26086_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_26097_, _20450_, _26086_);
  and (_26108_, _26097_, _15148_);
  not (_26119_, _24832_);
  not (_26130_, _24887_);
  and (_26141_, _25085_, _24942_);
  nor (_26152_, _26141_, _24930_);
  nor (_26163_, _26152_, _26130_);
  not (_26174_, _25194_);
  and (_26185_, _25448_, _25217_);
  nor (_26196_, _26185_, _25195_);
  nor (_26207_, _26196_, _26174_);
  nor (_26217_, _26207_, _25162_);
  nor (_26228_, _26217_, _25151_);
  and (_26239_, _26217_, _25151_);
  nor (_26250_, _26239_, _26228_);
  not (_26261_, _25470_);
  nor (_26272_, _25866_, _26261_);
  and (_26283_, _26272_, _25217_);
  and (_26294_, _26196_, _26174_);
  nor (_26305_, _26294_, _26207_);
  and (_26316_, _26305_, _26283_);
  not (_26326_, _26316_);
  nor (_26337_, _26326_, _26250_);
  nor (_26348_, _26217_, _25129_);
  or (_26359_, _26348_, _25140_);
  or (_26370_, _26359_, _26337_);
  and (_26381_, _26370_, _25107_);
  nor (_26392_, _25085_, _24942_);
  nor (_26403_, _26392_, _26141_);
  and (_26414_, _26403_, _26381_);
  and (_26425_, _26152_, _26130_);
  nor (_26436_, _26425_, _26163_);
  and (_26447_, _26436_, _26414_);
  or (_26458_, _26447_, _26163_);
  nor (_26479_, _26458_, _24865_);
  nor (_26480_, _26479_, _26119_);
  and (_26491_, _26479_, _26119_);
  nor (_26502_, _26491_, _26480_);
  and (_26513_, _26502_, _26108_);
  not (_26524_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_26535_, _15137_, _26524_);
  and (_26546_, _26535_, _26097_);
  not (_26557_, _26546_);
  nor (_26568_, _26557_, _24821_);
  and (_26578_, _26535_, _20461_);
  and (_26589_, _26578_, _24832_);
  nor (_26600_, _26589_, _26568_);
  and (_26611_, _26535_, _15104_);
  not (_26622_, _26611_);
  nor (_26633_, _26622_, _16367_);
  and (_26644_, _15137_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_26655_, _26644_, _20461_);
  not (_26666_, _26655_);
  nor (_26677_, _26666_, _18794_);
  nor (_26687_, _26677_, _26633_);
  and (_26698_, _26644_, _26097_);
  not (_26709_, _26698_);
  nor (_26720_, _26709_, _25866_);
  and (_26731_, _20483_, _15115_);
  and (_26742_, _26731_, _24810_);
  and (_26753_, _24777_, _20483_);
  and (_26774_, _26753_, _17192_);
  nor (_26775_, _26774_, _26742_);
  and (_26786_, _20461_, _15148_);
  not (_26796_, _26786_);
  nor (_26807_, _26796_, _17192_);
  not (_26818_, _26807_);
  nand (_26829_, _26818_, _26775_);
  nor (_26840_, _26829_, _26720_);
  and (_26851_, _26840_, _26687_);
  and (_26862_, _26644_, _24777_);
  nor (_26883_, _18794_, _18249_);
  and (_26884_, _26883_, _18435_);
  and (_26895_, _26884_, _17933_);
  and (_26906_, _26895_, _17574_);
  and (_26916_, _26906_, _17399_);
  and (_26927_, _26916_, _16388_);
  and (_26938_, _26927_, _25866_);
  not (_26949_, _25866_);
  and (_26960_, _16367_, _17388_);
  and (_26971_, _18794_, _18249_);
  and (_26982_, _26971_, _18424_);
  and (_26993_, _26982_, _17922_);
  and (_27004_, _26993_, _17563_);
  and (_27015_, _27004_, _26960_);
  and (_27026_, _27015_, _26949_);
  nor (_27037_, _27026_, _26938_);
  and (_27048_, _27037_, _17192_);
  nor (_27059_, _27037_, _17192_);
  nor (_27070_, _27059_, _27048_);
  and (_27081_, _27070_, _26862_);
  not (_27095_, _17018_);
  nor (_27096_, _25866_, _27095_);
  not (_27097_, _27096_);
  and (_27103_, _25866_, _17192_);
  and (_27114_, _26644_, _15115_);
  not (_27125_, _27114_);
  nor (_27136_, _27125_, _27103_);
  and (_27147_, _27136_, _27097_);
  nor (_27158_, _27147_, _27081_);
  and (_27169_, _26097_, _20483_);
  not (_27179_, _27169_);
  and (_27190_, _18424_, _18249_);
  nor (_27201_, _27190_, _17922_);
  and (_27212_, _27201_, _27169_);
  and (_27223_, _27212_, _17574_);
  not (_27234_, _27223_);
  and (_27245_, _27234_, _26960_);
  nor (_27256_, _26960_, _17192_);
  nor (_27267_, _27256_, _27212_);
  and (_27278_, _27267_, _25866_);
  nor (_27289_, _27278_, _27245_);
  and (_27299_, _27289_, _17192_);
  nor (_27310_, _27289_, _17192_);
  nor (_27321_, _27310_, _27299_);
  nor (_27342_, _27321_, _27179_);
  not (_27343_, _27342_);
  and (_27354_, _27343_, _27158_);
  and (_27365_, _27354_, _26851_);
  and (_27376_, _27365_, _26600_);
  not (_27387_, _27376_);
  nor (_27398_, _27387_, _26513_);
  and (_27409_, _27398_, _26075_);
  not (_27419_, _27409_);
  nor (_27430_, _27419_, _24755_);
  and (_27441_, _27430_, _24744_);
  not (_27452_, _27441_);
  or (_27463_, _27452_, _24723_);
  not (_27474_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_27485_, \oc8051_top_1.oc8051_decoder1.wr , _15093_);
  not (_27496_, _27485_);
  nor (_27507_, _27496_, _23429_);
  and (_27518_, _27507_, _27474_);
  not (_27529_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_27539_, _24723_, _27529_);
  and (_27550_, _27539_, _27518_);
  and (_27561_, _27550_, _27463_);
  nor (_27572_, _27507_, _27529_);
  not (_27583_, _26108_);
  nor (_27594_, _26480_, _24810_);
  nor (_27605_, _27594_, _27583_);
  not (_27626_, _27605_);
  and (_27627_, _17192_, _27095_);
  nor (_27638_, _27627_, _26031_);
  nor (_27649_, _27638_, _24799_);
  nor (_27660_, _27223_, _17399_);
  and (_27671_, _25866_, _16367_);
  and (_27681_, _27671_, _27660_);
  nor (_27692_, _27681_, _27103_);
  nor (_27703_, _25866_, _17192_);
  not (_27714_, _27703_);
  nor (_27725_, _27714_, _27245_);
  nor (_27736_, _27725_, _27179_);
  and (_27747_, _27736_, _27692_);
  or (_27758_, _27747_, _27212_);
  and (_27769_, _25822_, _25800_);
  and (_27780_, _26535_, _24777_);
  and (_27791_, _26731_, _25800_);
  nor (_27802_, _27791_, _27780_);
  nor (_27812_, _27802_, _27769_);
  not (_27823_, _27812_);
  nor (_27834_, _26796_, _25866_);
  nor (_27845_, _26709_, _18794_);
  and (_27856_, _26535_, _15115_);
  not (_27867_, _27856_);
  nor (_27878_, _27867_, _17192_);
  nor (_27889_, _27878_, _27845_);
  not (_27900_, _27889_);
  nor (_27911_, _27900_, _27834_);
  and (_27922_, _27911_, _27823_);
  nor (_27933_, _25855_, _25800_);
  not (_27938_, _26578_);
  nor (_27939_, _27938_, _25844_);
  nor (_27940_, _27939_, _26546_);
  nor (_27941_, _27940_, _27933_);
  nor (_27945_, _26753_, _26949_);
  and (_27956_, _26666_, _25855_);
  nor (_27967_, _27956_, _25844_);
  not (_27978_, _27967_);
  nor (_27989_, _27978_, _27945_);
  nor (_28000_, _27989_, _27941_);
  and (_28020_, _28000_, _27922_);
  not (_28021_, _28020_);
  nor (_28031_, _28021_, _27758_);
  not (_28041_, _28031_);
  nor (_28051_, _28041_, _27649_);
  and (_28062_, _28051_, _27626_);
  nor (_28072_, _24284_, _23670_);
  not (_28082_, _23812_);
  and (_28093_, _24152_, _28082_);
  and (_28103_, _28093_, _28072_);
  not (_28113_, _24416_);
  nor (_28123_, _24668_, _24547_);
  and (_28134_, _28123_, _28113_);
  and (_28145_, _28134_, _28103_);
  nand (_28155_, _28145_, _28062_);
  and (_28166_, _27507_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_28176_, _28145_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_28194_, _28176_, _28166_);
  and (_28195_, _28194_, _28155_);
  or (_28205_, _28195_, _27572_);
  or (_28216_, _28205_, _27561_);
  and (_35966_[7], _28216_, _35583_);
  and (_28236_, _22920_, _20494_);
  not (_28247_, _28236_);
  and (_28258_, _20216_, _15159_);
  and (_28268_, _25866_, _26261_);
  nor (_28278_, _28268_, _26272_);
  nor (_28289_, _26108_, _24788_);
  not (_28300_, _28289_);
  and (_28310_, _28300_, _28278_);
  not (_28321_, _28310_);
  nor (_28332_, _27867_, _25866_);
  not (_28342_, _28332_);
  nor (_28352_, _27938_, _25448_);
  nor (_28363_, _28352_, _26546_);
  or (_28372_, _28363_, _25459_);
  and (_28380_, _26644_, _26086_);
  not (_28387_, _28380_);
  nor (_28395_, _28387_, _18249_);
  and (_28403_, _27780_, _17203_);
  nor (_28410_, _28403_, _28395_);
  and (_28418_, _26731_, _25448_);
  and (_28426_, _26753_, _18794_);
  nor (_28433_, _28426_, _28418_);
  nor (_28434_, _27125_, _15877_);
  and (_28435_, _26862_, _18794_);
  nor (_28436_, _28435_, _28434_);
  nor (_28442_, _26786_, _27169_);
  nor (_28453_, _28442_, _18794_);
  not (_28464_, _28453_);
  and (_28475_, _28464_, _28436_);
  and (_28485_, _28475_, _28433_);
  and (_28496_, _28485_, _28410_);
  and (_28507_, _28496_, _28372_);
  and (_28516_, _28507_, _28342_);
  and (_28523_, _28516_, _28321_);
  not (_28534_, _28523_);
  nor (_28545_, _28534_, _28258_);
  and (_28556_, _28545_, _28247_);
  not (_28567_, _28556_);
  or (_28578_, _28567_, _24723_);
  not (_28589_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_28600_, _24723_, _28589_);
  and (_28611_, _28600_, _27518_);
  and (_28622_, _28611_, _28578_);
  nor (_28633_, _27507_, _28589_);
  not (_28654_, _28062_);
  or (_28655_, _28654_, _24723_);
  and (_28666_, _28600_, _28166_);
  and (_28677_, _28666_, _28655_);
  or (_28688_, _28677_, _28633_);
  or (_28699_, _28688_, _28622_);
  and (_35966_[0], _28699_, _35583_);
  and (_28720_, _20248_, _15159_);
  not (_28731_, _28720_);
  and (_28742_, _22985_, _20494_);
  nor (_28753_, _25448_, _25217_);
  or (_28764_, _28753_, _26185_);
  and (_28775_, _28764_, _26272_);
  nor (_28786_, _28764_, _26272_);
  or (_28797_, _28786_, _28775_);
  and (_28808_, _28797_, _26108_);
  nor (_28819_, _25877_, _25437_);
  nor (_28830_, _28819_, _25888_);
  nor (_28841_, _28830_, _24799_);
  not (_28852_, _28841_);
  nor (_28863_, _27201_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_28874_, _28863_, _18260_);
  nor (_28885_, _28863_, _18260_);
  nor (_28896_, _28885_, _28874_);
  nor (_28907_, _28896_, _27179_);
  not (_28918_, _28907_);
  and (_28929_, _26578_, _25217_);
  nor (_28940_, _26557_, _25206_);
  not (_28951_, _28940_);
  and (_28962_, _26731_, _25195_);
  and (_28973_, _26753_, _18249_);
  nor (_28984_, _28973_, _28962_);
  nand (_28995_, _28984_, _28951_);
  nor (_29006_, _28995_, _28929_);
  nor (_29017_, _26622_, _18794_);
  not (_29028_, _29017_);
  nor (_29039_, _26796_, _18249_);
  nor (_29050_, _28387_, _18424_);
  nor (_29061_, _29050_, _29039_);
  and (_29071_, _29061_, _29028_);
  and (_29082_, _29071_, _29006_);
  and (_29093_, _29082_, _28918_);
  and (_29103_, _29093_, _28852_);
  nor (_29114_, _27125_, _16843_);
  nor (_29125_, _26971_, _26883_);
  not (_29135_, _29125_);
  nor (_29146_, _29135_, _25866_);
  and (_29157_, _29135_, _25866_);
  nor (_29168_, _29157_, _29146_);
  and (_29178_, _29168_, _26862_);
  nor (_29199_, _29178_, _29114_);
  nand (_29200_, _29199_, _29103_);
  nor (_29210_, _29200_, _28808_);
  not (_29221_, _29210_);
  nor (_29232_, _29221_, _28742_);
  and (_29242_, _29232_, _28731_);
  not (_29253_, _29242_);
  or (_29264_, _29253_, _24723_);
  not (_29274_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_29285_, _24723_, _29274_);
  and (_29296_, _29285_, _27518_);
  and (_29307_, _29296_, _29264_);
  nor (_29318_, _27507_, _29274_);
  and (_29329_, _24679_, _28113_);
  and (_29340_, _29329_, _28103_);
  or (_29351_, _29340_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_29362_, _29351_, _28166_);
  nand (_29373_, _29340_, _28062_);
  and (_29384_, _29373_, _29362_);
  or (_29395_, _29384_, _29318_);
  or (_29406_, _29395_, _29307_);
  and (_35966_[1], _29406_, _35583_);
  and (_29427_, _20280_, _15159_);
  not (_29438_, _29427_);
  and (_29459_, _23050_, _20494_);
  nor (_29460_, _27125_, _15551_);
  and (_29471_, _26883_, _25866_);
  and (_29482_, _26971_, _26949_);
  nor (_29493_, _29482_, _29471_);
  and (_29504_, _29493_, _18424_);
  nor (_29515_, _29493_, _18424_);
  nor (_29526_, _29515_, _29504_);
  and (_29537_, _29526_, _26862_);
  nor (_29548_, _29537_, _29460_);
  nor (_29559_, _25888_, _25404_);
  nor (_29570_, _29559_, _25899_);
  nor (_29581_, _29570_, _24799_);
  not (_29592_, _29581_);
  nor (_29603_, _28387_, _17922_);
  and (_29614_, _26731_, _25162_);
  and (_29625_, _26753_, _18424_);
  nor (_29636_, _29625_, _29614_);
  nor (_29647_, _26557_, _25173_);
  and (_29658_, _26578_, _25194_);
  nor (_29669_, _29658_, _29647_);
  nor (_29680_, _26622_, _18249_);
  nor (_29691_, _26796_, _18424_);
  nor (_29702_, _29691_, _29680_);
  and (_29713_, _29702_, _29669_);
  nand (_29724_, _29713_, _29636_);
  nor (_29735_, _29724_, _29603_);
  and (_29746_, _29735_, _29592_);
  nor (_29767_, _26305_, _26283_);
  nor (_29768_, _29767_, _27583_);
  and (_29779_, _29768_, _26326_);
  nor (_29790_, _28885_, _18424_);
  and (_29801_, _27190_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_29812_, _29801_, _29790_);
  nor (_29823_, _29812_, _27179_);
  nor (_29833_, _29823_, _29779_);
  and (_29844_, _29833_, _29746_);
  and (_29855_, _29844_, _29548_);
  not (_29866_, _29855_);
  nor (_29876_, _29866_, _29459_);
  and (_29887_, _29876_, _29438_);
  not (_29898_, _29887_);
  or (_29908_, _29898_, _24723_);
  not (_29919_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_29930_, _24723_, _29919_);
  and (_29940_, _29930_, _27518_);
  and (_29951_, _29940_, _29908_);
  nor (_29962_, _27507_, _29919_);
  nor (_29972_, _24547_, _24416_);
  nand (_29983_, _24668_, _28103_);
  or (_29994_, _29983_, _29972_);
  and (_30005_, _29994_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_30016_, _24547_);
  and (_30027_, _24668_, _30016_);
  and (_30038_, _30027_, _24416_);
  and (_30039_, _30038_, _28654_);
  and (_30040_, _24679_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_30041_, _30040_, _30039_);
  and (_30042_, _30041_, _28103_);
  or (_30043_, _30042_, _30005_);
  and (_30044_, _30043_, _28166_);
  or (_30045_, _30044_, _29962_);
  or (_30046_, _30045_, _29951_);
  and (_35966_[2], _30046_, _35583_);
  and (_30047_, _20322_, _15159_);
  not (_30048_, _30047_);
  and (_30049_, _23115_, _20494_);
  nor (_30050_, _25899_, _25371_);
  nor (_30051_, _30050_, _25920_);
  nor (_30052_, _30051_, _24799_);
  not (_30053_, _30052_);
  not (_30054_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_30055_, _27190_, _30054_);
  nor (_30056_, _30055_, _17933_);
  or (_30057_, _30056_, _27179_);
  or (_30058_, _30057_, _27201_);
  and (_30059_, _26731_, _25140_);
  and (_30060_, _26753_, _17922_);
  nor (_30061_, _30060_, _30059_);
  nor (_30062_, _28387_, _17563_);
  nor (_30063_, _26796_, _17922_);
  nor (_30064_, _26622_, _18424_);
  or (_30065_, _30064_, _30063_);
  nor (_30066_, _30065_, _30062_);
  and (_30067_, _30066_, _30061_);
  and (_30068_, _30067_, _30058_);
  and (_30069_, _26326_, _26250_);
  or (_30070_, _30069_, _27583_);
  nor (_30071_, _30070_, _26337_);
  nor (_30072_, _27125_, _16541_);
  and (_30073_, _26884_, _25866_);
  and (_30074_, _26982_, _26949_);
  nor (_30075_, _30074_, _30073_);
  nor (_30076_, _30075_, _17922_);
  not (_30077_, _30076_);
  not (_30078_, _26862_);
  and (_30079_, _30075_, _17922_);
  nor (_30080_, _30079_, _30078_);
  and (_30081_, _30080_, _30077_);
  nor (_30082_, _30081_, _30072_);
  nor (_30083_, _26557_, _25129_);
  and (_30084_, _26578_, _25151_);
  nor (_30085_, _30084_, _30083_);
  nand (_30086_, _30085_, _30082_);
  nor (_30087_, _30086_, _30071_);
  and (_30088_, _30087_, _30068_);
  and (_30089_, _30088_, _30053_);
  not (_30090_, _30089_);
  nor (_30091_, _30090_, _30049_);
  and (_30092_, _30091_, _30048_);
  not (_30093_, _30092_);
  or (_30094_, _30093_, _24723_);
  not (_30095_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_30096_, _24723_, _30095_);
  and (_30097_, _30096_, _27518_);
  and (_30098_, _30097_, _30094_);
  nor (_30099_, _27507_, _30095_);
  and (_30100_, _29983_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_30101_, _29972_, _24668_);
  and (_30102_, _30101_, _28654_);
  not (_30103_, _24668_);
  or (_30104_, _29972_, _30103_);
  nor (_30105_, _30104_, _30095_);
  or (_30106_, _30105_, _30102_);
  and (_30107_, _30106_, _28103_);
  or (_30108_, _30107_, _30100_);
  and (_30109_, _30108_, _28166_);
  or (_30110_, _30109_, _30099_);
  or (_30111_, _30110_, _30098_);
  and (_35966_[3], _30111_, _35583_);
  and (_30112_, _23179_, _20494_);
  not (_30113_, _30112_);
  and (_30114_, _20354_, _15159_);
  nor (_30115_, _25976_, _25107_);
  and (_30116_, _25976_, _25107_);
  nor (_30117_, _30116_, _30115_);
  and (_30118_, _30117_, _24788_);
  not (_30119_, _30118_);
  nor (_30120_, _26370_, _25107_);
  not (_30121_, _30120_);
  nor (_30122_, _27583_, _26381_);
  and (_30123_, _30122_, _30121_);
  and (_30124_, _26895_, _25866_);
  and (_30125_, _26993_, _26949_);
  nor (_30126_, _30125_, _30124_);
  and (_30127_, _30126_, _17563_);
  nor (_30128_, _30126_, _17563_);
  nor (_30129_, _30128_, _30127_);
  and (_30130_, _30129_, _26862_);
  nor (_30131_, _25866_, _15714_);
  and (_30132_, _25866_, _17574_);
  nor (_30133_, _30132_, _30131_);
  nor (_30134_, _30133_, _27125_);
  and (_30135_, _26731_, _25085_);
  and (_30136_, _26753_, _17563_);
  nor (_30137_, _30136_, _30135_);
  and (_30138_, _26578_, _25107_);
  nor (_30139_, _26557_, _25096_);
  or (_30140_, _30139_, _30138_);
  not (_30141_, _30140_);
  and (_30142_, _30141_, _30137_);
  not (_30143_, _30142_);
  or (_30144_, _30143_, _30134_);
  nor (_30145_, _30144_, _30130_);
  nor (_30146_, _27212_, _17574_);
  nor (_30147_, _26796_, _17563_);
  nor (_30148_, _27223_, _27179_);
  nor (_30149_, _30148_, _30147_);
  or (_30150_, _30149_, _30146_);
  nor (_30151_, _28387_, _17388_);
  nor (_30152_, _26622_, _17922_);
  nor (_30153_, _30152_, _30151_);
  and (_30154_, _30153_, _30150_);
  and (_30155_, _30154_, _30145_);
  not (_30156_, _30155_);
  nor (_30157_, _30156_, _30123_);
  and (_30158_, _30157_, _30119_);
  not (_30159_, _30158_);
  nor (_30160_, _30159_, _30114_);
  and (_30161_, _30160_, _30113_);
  not (_30162_, _30161_);
  or (_30163_, _30162_, _24723_);
  not (_30164_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_30165_, _24723_, _30164_);
  and (_30166_, _30165_, _27518_);
  and (_30167_, _30166_, _30163_);
  nor (_30168_, _27507_, _30164_);
  not (_30169_, _28103_);
  and (_30170_, _24547_, _24416_);
  and (_30171_, _30170_, _30103_);
  nor (_30172_, _30170_, _30103_);
  nor (_30173_, _30172_, _30171_);
  or (_30174_, _30173_, _30169_);
  and (_30175_, _30174_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_30176_, _30171_, _28654_);
  and (_30177_, _30172_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_30178_, _30177_, _30176_);
  and (_30179_, _30178_, _28103_);
  or (_30180_, _30179_, _30175_);
  and (_30181_, _30180_, _28166_);
  or (_30182_, _30181_, _30168_);
  or (_30183_, _30182_, _30167_);
  and (_35966_[4], _30183_, _35583_);
  and (_30184_, _23244_, _20494_);
  not (_30185_, _30184_);
  and (_30186_, _20397_, _15159_);
  nor (_30187_, _26403_, _26381_);
  nor (_30188_, _30187_, _26414_);
  and (_30189_, _30188_, _26108_);
  not (_30190_, _30189_);
  nor (_30191_, _25987_, _25074_);
  nor (_30192_, _30191_, _25998_);
  nor (_30193_, _30192_, _24799_);
  nor (_30194_, _25866_, _16680_);
  and (_30195_, _25866_, _17399_);
  nor (_30196_, _30195_, _30194_);
  nor (_30197_, _30196_, _27125_);
  and (_30198_, _26906_, _25866_);
  and (_30199_, _27004_, _26949_);
  nor (_30200_, _30199_, _30198_);
  and (_30201_, _30200_, _17388_);
  nor (_30202_, _30200_, _17388_);
  or (_30203_, _30202_, _30078_);
  nor (_30204_, _30203_, _30201_);
  nor (_30205_, _30204_, _30197_);
  not (_30206_, _27278_);
  and (_30207_, _30206_, _27660_);
  nor (_30208_, _27278_, _27223_);
  nor (_30209_, _30208_, _17388_);
  nor (_30210_, _30209_, _30207_);
  nor (_30211_, _30210_, _27179_);
  and (_30212_, _26578_, _24942_);
  not (_30213_, _30212_);
  nor (_30214_, _26557_, _24931_);
  not (_30215_, _30214_);
  and (_30216_, _26731_, _24930_);
  and (_30217_, _26753_, _17388_);
  nor (_30218_, _30217_, _30216_);
  and (_30219_, _30218_, _30215_);
  and (_30220_, _30219_, _30213_);
  nor (_30221_, _28387_, _16367_);
  not (_30222_, _30221_);
  nor (_30223_, _26796_, _17388_);
  nor (_30224_, _26622_, _17563_);
  nor (_30225_, _30224_, _30223_);
  and (_30226_, _30225_, _30222_);
  and (_30227_, _30226_, _30220_);
  not (_30228_, _30227_);
  nor (_30229_, _30228_, _30211_);
  and (_30230_, _30229_, _30205_);
  not (_30231_, _30230_);
  nor (_30232_, _30231_, _30193_);
  and (_30233_, _30232_, _30190_);
  not (_30234_, _30233_);
  nor (_30235_, _30234_, _30186_);
  and (_30236_, _30235_, _30185_);
  not (_30237_, _30236_);
  or (_30238_, _30237_, _24723_);
  not (_30239_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_30240_, _24723_, _30239_);
  and (_30241_, _30240_, _27518_);
  and (_30242_, _30241_, _30238_);
  nor (_30243_, _27507_, _30239_);
  and (_30244_, _30103_, _24547_);
  nor (_30245_, _30244_, _30027_);
  or (_30246_, _30245_, _30169_);
  and (_30247_, _30246_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_30248_, _24547_, _28113_);
  and (_30249_, _30248_, _30103_);
  and (_30250_, _30249_, _28654_);
  or (_30251_, _30171_, _30027_);
  and (_30252_, _30251_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_30253_, _30252_, _30250_);
  and (_30254_, _30253_, _28103_);
  or (_30255_, _30254_, _30247_);
  and (_30256_, _30255_, _28166_);
  or (_30257_, _30256_, _30243_);
  or (_30258_, _30257_, _30242_);
  and (_35966_[5], _30258_, _35583_);
  and (_30259_, _23309_, _20494_);
  not (_30260_, _30259_);
  and (_30261_, _20429_, _15159_);
  nor (_30262_, _26436_, _26414_);
  not (_30263_, _30262_);
  nor (_30264_, _27583_, _26447_);
  and (_30265_, _30264_, _30263_);
  not (_30266_, _30265_);
  nor (_30267_, _25998_, _25041_);
  nor (_30268_, _30267_, _26009_);
  nor (_30269_, _30268_, _24799_);
  nor (_30270_, _25866_, _24843_);
  or (_30271_, _30270_, _27125_);
  nor (_30272_, _30271_, _27671_);
  or (_30273_, _25866_, _17388_);
  or (_30274_, _30199_, _26916_);
  and (_30275_, _30274_, _30273_);
  and (_30276_, _30275_, _16388_);
  nor (_30277_, _30275_, _16388_);
  or (_30278_, _30277_, _30078_);
  nor (_30279_, _30278_, _30276_);
  nor (_30280_, _30279_, _30272_);
  nor (_30281_, _30207_, _16367_);
  and (_30282_, _30207_, _16367_);
  nor (_30283_, _30282_, _30281_);
  nor (_30284_, _30283_, _27179_);
  and (_30285_, _26578_, _24887_);
  not (_30286_, _30285_);
  nor (_30287_, _26557_, _24876_);
  not (_30288_, _30287_);
  and (_30289_, _26731_, _24865_);
  and (_30290_, _26753_, _16367_);
  nor (_30291_, _30290_, _30289_);
  and (_30292_, _30291_, _30288_);
  and (_30293_, _30292_, _30286_);
  nor (_30294_, _28387_, _17192_);
  not (_30295_, _30294_);
  nor (_30296_, _26796_, _16367_);
  nor (_30297_, _26622_, _17388_);
  nor (_30298_, _30297_, _30296_);
  and (_30299_, _30298_, _30295_);
  and (_30300_, _30299_, _30293_);
  not (_30301_, _30300_);
  nor (_30302_, _30301_, _30284_);
  and (_30303_, _30302_, _30280_);
  not (_30304_, _30303_);
  nor (_30305_, _30304_, _30269_);
  and (_30306_, _30305_, _30266_);
  not (_30307_, _30306_);
  nor (_30308_, _30307_, _30261_);
  and (_30309_, _30308_, _30260_);
  not (_30310_, _30309_);
  or (_30311_, _30310_, _24723_);
  not (_30312_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_30313_, _24723_, _30312_);
  and (_30314_, _30313_, _27518_);
  and (_30315_, _30314_, _30311_);
  nor (_30316_, _27507_, _30312_);
  not (_30317_, _28134_);
  nand (_30318_, _30317_, _28103_);
  and (_30319_, _30318_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_30320_, _28123_, _24416_);
  and (_30321_, _30320_, _28654_);
  nor (_30322_, _28123_, _30312_);
  or (_30323_, _30322_, _30321_);
  and (_30324_, _30323_, _28103_);
  or (_30325_, _30324_, _30319_);
  and (_30326_, _30325_, _28166_);
  or (_30327_, _30326_, _30316_);
  or (_30328_, _30327_, _30315_);
  and (_35966_[6], _30328_, _35583_);
  and (_30329_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_30330_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_30331_, _30330_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_30332_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_30333_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_30334_, _30333_, _30332_);
  and (_30335_, _30330_, _15093_);
  and (_30336_, _30335_, _30334_);
  not (_30337_, _30336_);
  and (_30338_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30339_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_30340_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_30341_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_30342_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_30343_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30344_, _30343_, _30342_);
  and (_30345_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  not (_30346_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30347_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _30346_);
  and (_30348_, _30347_, _30342_);
  and (_30349_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_30350_, _30349_, _30345_);
  nor (_30351_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30352_, _30351_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_30353_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  not (_30354_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_30355_, _30354_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_30356_, _30355_, _30342_);
  and (_30357_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_30358_, _30357_, _30353_);
  and (_30359_, _30358_, _30350_);
  nor (_30360_, _30351_, _30342_);
  and (_30361_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_30362_, _30351_, _30342_);
  and (_30363_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_30364_, _30363_, _30361_);
  and (_30365_, _30364_, _30359_);
  nor (_30366_, _30365_, _30341_);
  and (_30367_, _30366_, _30340_);
  nor (_30368_, _30367_, _30339_);
  nor (_30369_, _30368_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_30370_, _30369_, _30338_);
  nor (_30371_, _30370_, _30337_);
  and (_30372_, _30334_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_30373_, _30372_, _30337_);
  nor (_30374_, _30373_, _30371_);
  not (_30375_, _30374_);
  and (_30376_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not (_30377_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30378_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_30379_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_30380_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_30381_, _30380_, _30379_);
  and (_30382_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_30383_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_30384_, _30383_, _30382_);
  and (_30385_, _30384_, _30381_);
  and (_30386_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_30387_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_30388_, _30387_, _30386_);
  and (_30389_, _30388_, _30385_);
  nor (_30390_, _30389_, _30341_);
  and (_30391_, _30390_, _30340_);
  or (_30392_, _30391_, _30378_);
  and (_30393_, _30392_, _30377_);
  nor (_30394_, _30393_, _30376_);
  nor (_30395_, _30394_, _30337_);
  and (_30396_, _30334_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_30397_, _30396_, _30337_);
  nor (_30398_, _30397_, _30395_);
  and (_30399_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and (_30400_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_30401_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_30402_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_30403_, _30402_, _30401_);
  and (_30404_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_30405_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_30406_, _30405_, _30404_);
  and (_30407_, _30406_, _30403_);
  and (_30408_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_30409_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_30410_, _30409_, _30408_);
  and (_30411_, _30410_, _30407_);
  nor (_30412_, _30411_, _30341_);
  and (_30413_, _30412_, _30340_);
  or (_30414_, _30413_, _30400_);
  and (_30415_, _30414_, _30377_);
  nor (_30416_, _30415_, _30399_);
  nor (_30417_, _30416_, _30337_);
  and (_30418_, _30334_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_30419_, _30418_, _30337_);
  nor (_30420_, _30419_, _30417_);
  not (_30421_, _30420_);
  and (_30422_, _30421_, _30398_);
  and (_30423_, _30422_, _30375_);
  and (_30424_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30425_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_30426_, _30341_);
  and (_30427_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_30428_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_30429_, _30428_, _30427_);
  and (_30430_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_30431_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_30432_, _30431_, _30430_);
  and (_30433_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_30434_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_30435_, _30434_, _30433_);
  and (_30436_, _30435_, _30432_);
  and (_30437_, _30436_, _30429_);
  and (_30438_, _30437_, _30426_);
  nor (_30439_, _30438_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  or (_30440_, _30439_, _30425_);
  and (_30441_, _30440_, _30377_);
  nor (_30442_, _30441_, _30424_);
  nor (_30443_, _30442_, _30337_);
  and (_30444_, _30334_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_30445_, _30444_, _30337_);
  nor (_30446_, _30445_, _30443_);
  and (_30447_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30448_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_30449_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_30450_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_30451_, _30450_, _30449_);
  and (_30452_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_30453_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_30454_, _30453_, _30452_);
  and (_30455_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_30456_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_30457_, _30456_, _30455_);
  and (_30458_, _30457_, _30454_);
  and (_30459_, _30458_, _30451_);
  or (_30460_, _30341_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_30461_, _30460_, _30459_);
  nor (_30462_, _30461_, _30448_);
  nor (_30463_, _30462_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_30464_, _30463_, _30447_);
  nor (_30465_, _30464_, _30337_);
  and (_30466_, _30334_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_30467_, _30466_, _30337_);
  nor (_30468_, _30467_, _30465_);
  nor (_30469_, _30468_, _30446_);
  and (_30470_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30471_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_30472_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and (_30473_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_30474_, _30473_, _30472_);
  and (_30475_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_30476_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_30477_, _30476_, _30475_);
  and (_30478_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_30479_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_30480_, _30479_, _30478_);
  and (_30481_, _30480_, _30477_);
  and (_30482_, _30481_, _30474_);
  nor (_30483_, _30482_, _30341_);
  and (_30484_, _30483_, _30340_);
  or (_30485_, _30484_, _30471_);
  and (_30486_, _30485_, _30377_);
  nor (_30487_, _30486_, _30470_);
  nor (_30488_, _30487_, _30337_);
  and (_30489_, _30334_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_30490_, _30489_, _30337_);
  nor (_30491_, _30490_, _30488_);
  and (_30492_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_30493_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_30494_, _30493_, _30492_);
  and (_30495_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_30496_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_30497_, _30496_, _30495_);
  and (_30498_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_30499_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_30500_, _30499_, _30498_);
  and (_30501_, _30500_, _30497_);
  and (_30502_, _30501_, _30494_);
  not (_30503_, _30502_);
  nor (_30504_, _30503_, _30460_);
  nor (_30505_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _30340_);
  or (_30506_, _30505_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_30507_, _30506_, _30504_);
  and (_30508_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  or (_30509_, _30508_, _30507_);
  and (_30510_, _30509_, _30336_);
  and (_30511_, _30334_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_30512_, _30511_, _30337_);
  nor (_30513_, _30512_, _30510_);
  not (_30514_, _30513_);
  and (_30515_, _30514_, _30491_);
  and (_30516_, _30515_, _30469_);
  and (_30517_, _30516_, _30423_);
  and (_30518_, _30469_, _30491_);
  and (_30519_, _30420_, _30398_);
  and (_30520_, _30519_, _30374_);
  and (_30521_, _30520_, _30518_);
  nor (_30522_, _30521_, _30517_);
  and (_30523_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and (_30524_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and (_30525_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_30526_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_30527_, _30526_, _30525_);
  and (_30528_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_30529_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_30530_, _30529_, _30528_);
  and (_30531_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_30532_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_30533_, _30532_, _30531_);
  and (_30534_, _30533_, _30530_);
  and (_30535_, _30534_, _30527_);
  nor (_30536_, _30535_, _30341_);
  and (_30537_, _30536_, _30340_);
  nor (_30538_, _30537_, _30524_);
  nor (_30539_, _30538_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor (_30540_, _30539_, _30523_);
  nor (_30541_, _30540_, _30337_);
  and (_30542_, _30334_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_30543_, _30542_, _30337_);
  nor (_30544_, _30543_, _30541_);
  not (_30545_, _30446_);
  and (_30546_, _30491_, _30468_);
  and (_30547_, _30546_, _30545_);
  and (_30548_, _30547_, _30544_);
  and (_30549_, _30519_, _30375_);
  and (_30550_, _30549_, _30548_);
  and (_30551_, _30513_, _30518_);
  not (_30552_, _30398_);
  and (_30553_, _30420_, _30552_);
  and (_30554_, _30553_, _30374_);
  nor (_30555_, _30420_, _30398_);
  and (_30556_, _30555_, _30375_);
  or (_30557_, _30556_, _30554_);
  and (_30558_, _30557_, _30551_);
  nor (_30559_, _30558_, _30550_);
  and (_30560_, _30559_, _30522_);
  and (_30561_, _30555_, _30374_);
  and (_30562_, _30561_, _30518_);
  and (_30563_, _30422_, _30374_);
  and (_30564_, _30563_, _30516_);
  nor (_30565_, _30564_, _30562_);
  not (_30566_, _30565_);
  not (_30567_, _30518_);
  and (_30568_, _30554_, _30514_);
  nor (_30569_, _30568_, _30549_);
  nor (_30570_, _30569_, _30567_);
  nor (_30571_, _30570_, _30566_);
  and (_30572_, _30571_, _30560_);
  and (_30573_, _30423_, _30513_);
  not (_30574_, _30544_);
  and (_30575_, _30547_, _30574_);
  and (_30576_, _30575_, _30573_);
  not (_30577_, _30576_);
  nor (_30578_, _30398_, _30374_);
  and (_30579_, _30578_, _30420_);
  and (_30580_, _30579_, _30514_);
  and (_30581_, _30580_, _30575_);
  and (_30582_, _30563_, _30514_);
  and (_30583_, _30575_, _30582_);
  nor (_30584_, _30583_, _30581_);
  and (_30585_, _30584_, _30577_);
  and (_30586_, _30561_, _30514_);
  and (_30587_, _30544_, _30446_);
  and (_30588_, _30587_, _30546_);
  and (_30589_, _30588_, _30586_);
  not (_30590_, _30589_);
  and (_30591_, _30579_, _30513_);
  and (_30592_, _30591_, _30518_);
  and (_30593_, _30374_, _30513_);
  and (_30594_, _30593_, _30422_);
  and (_30595_, _30594_, _30518_);
  nor (_30596_, _30595_, _30592_);
  and (_30597_, _30596_, _30590_);
  and (_30598_, _30597_, _30585_);
  and (_30599_, _30598_, _30572_);
  nor (_30600_, _30599_, _30331_);
  not (_30601_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_30602_, _15093_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_30603_, _30602_, _30601_);
  and (_30604_, _30603_, _30588_);
  and (_30605_, _30604_, _30579_);
  and (_30606_, _30550_, _30602_);
  and (_30607_, _30606_, \oc8051_top_1.oc8051_decoder1.state [0]);
  or (_30608_, _30607_, _30605_);
  nor (_30609_, _30608_, _30600_);
  nor (_30610_, _30609_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_30611_, _30610_, _30329_);
  and (_30612_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_30613_, _30468_);
  and (_30614_, _30491_, _30613_);
  and (_30615_, _30574_, _30446_);
  and (_30616_, _30615_, _30614_);
  and (_30617_, _30616_, _30586_);
  not (_30618_, _30617_);
  and (_30619_, _30580_, _30548_);
  and (_30620_, _30593_, _30553_);
  and (_30621_, _30620_, _30547_);
  nor (_30622_, _30621_, _30619_);
  and (_30623_, _30622_, _30618_);
  and (_30624_, _30423_, _30514_);
  and (_30625_, _30548_, _30624_);
  and (_30626_, _30561_, _30513_);
  and (_30627_, _30626_, _30548_);
  nor (_30628_, _30627_, _30625_);
  and (_30629_, _30620_, _30616_);
  and (_30630_, _30588_, _30573_);
  nor (_30631_, _30630_, _30629_);
  and (_30632_, _30520_, _30514_);
  and (_30633_, _30632_, _30616_);
  and (_30634_, _30588_, _30624_);
  nor (_30635_, _30634_, _30633_);
  and (_30636_, _30635_, _30631_);
  and (_30637_, _30636_, _30628_);
  and (_30638_, _30637_, _30623_);
  and (_30639_, _30588_, _30561_);
  and (_30640_, _30591_, _30547_);
  nor (_30641_, _30640_, _30639_);
  and (_30642_, _30582_, _30548_);
  and (_30643_, _30616_, _30594_);
  nor (_30644_, _30643_, _30642_);
  and (_30645_, _30644_, _30641_);
  and (_30646_, _30594_, _30548_);
  and (_30647_, _30568_, _30547_);
  nor (_30648_, _30647_, _30646_);
  not (_30649_, _30648_);
  and (_30650_, _30422_, _30514_);
  and (_30651_, _30650_, _30616_);
  nor (_30652_, _30651_, _30649_);
  and (_30653_, _30652_, _30645_);
  not (_30654_, _30616_);
  nor (_30655_, _30654_, _30569_);
  and (_30656_, _30556_, _30513_);
  and (_30657_, _30656_, _30616_);
  nor (_30658_, _30657_, _30550_);
  not (_30659_, _30658_);
  nor (_30660_, _30659_, _30655_);
  and (_30661_, _30586_, _30548_);
  and (_30662_, _30573_, _30548_);
  nor (_30663_, _30662_, _30661_);
  and (_30664_, _30616_, _30591_);
  and (_30665_, _30626_, _30616_);
  nor (_30666_, _30665_, _30664_);
  and (_30667_, _30666_, _30663_);
  and (_30668_, _30667_, _30660_);
  and (_30669_, _30588_, _30549_);
  and (_30670_, _30669_, _30513_);
  not (_30671_, _30588_);
  and (_30672_, _30549_, _30514_);
  nor (_30673_, _30632_, _30672_);
  nor (_30674_, _30673_, _30671_);
  nor (_30675_, _30674_, _30670_);
  and (_30676_, _30593_, _30519_);
  and (_30677_, _30676_, _30616_);
  not (_30678_, _30677_);
  and (_30679_, _30551_, _30423_);
  not (_30680_, _30491_);
  and (_30681_, _30573_, _30680_);
  nor (_30682_, _30681_, _30679_);
  and (_30683_, _30682_, _30678_);
  and (_30684_, _30683_, _30675_);
  and (_30685_, _30684_, _30668_);
  and (_30686_, _30685_, _30653_);
  and (_30687_, _30686_, _30638_);
  nor (_30688_, _30687_, _30331_);
  and (_30689_, _30602_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_30690_, _30689_, _30550_);
  not (_30691_, _30690_);
  and (_30692_, _30588_, _30553_);
  and (_30693_, _30692_, _30603_);
  not (_30694_, _30603_);
  nor (_30695_, _30374_, _30514_);
  and (_30696_, _30695_, _30519_);
  and (_30697_, _30588_, _30696_);
  and (_30698_, _30632_, _30588_);
  nor (_30699_, _30698_, _30697_);
  nor (_30700_, _30699_, _30694_);
  nor (_30701_, _30700_, _30693_);
  and (_30702_, _30701_, _30691_);
  not (_30703_, _30702_);
  nor (_30704_, _30703_, _30688_);
  nor (_30705_, _30704_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_30706_, _30705_, _30612_);
  nor (_30707_, _30706_, _30611_);
  and (_30708_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_30709_, _30587_, _30614_);
  and (_30710_, _30709_, _30594_);
  and (_30711_, _30709_, _30573_);
  nor (_30712_, _30711_, _30710_);
  and (_30713_, _30712_, _30585_);
  nor (_30714_, _30713_, _30331_);
  not (_30715_, _30714_);
  not (_30716_, _30330_);
  nor (_30717_, _30712_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_30718_, _30717_, _30716_);
  nor (_30719_, _30718_, _30693_);
  and (_30720_, _30719_, _30715_);
  nor (_30721_, _30720_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_30722_, _30721_, _30708_);
  and (_30723_, _30722_, _35583_);
  and (_35974_, _30723_, _30707_);
  and (_30724_, _24141_, _24284_);
  not (_30725_, _23670_);
  nor (_30726_, _23812_, _30725_);
  and (_30727_, _30726_, _30724_);
  and (_30728_, _30727_, _24009_);
  and (_30729_, _30728_, _29329_);
  and (_30730_, _30729_, _27518_);
  not (_30731_, _30730_);
  and (_30732_, _30731_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_30733_, _20494_, _15159_);
  and (_30734_, _26097_, _20472_);
  nor (_30735_, _26786_, _30734_);
  and (_30736_, _30735_, _26622_);
  and (_30737_, _30736_, _30733_);
  and (_30738_, _30737_, _28387_);
  nor (_30739_, _30738_, _16367_);
  not (_30740_, _30739_);
  and (_30741_, _30740_, _30293_);
  and (_30742_, _30741_, _30280_);
  nor (_30743_, _30742_, _30731_);
  nor (_30744_, _30743_, _30732_);
  and (_30745_, _30731_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_30746_, _30738_, _17388_);
  not (_30747_, _30746_);
  and (_30748_, _30747_, _30220_);
  and (_30749_, _30748_, _30205_);
  nor (_30750_, _30749_, _30731_);
  nor (_30751_, _30750_, _30745_);
  and (_30752_, _30731_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_30753_, _30738_, _17563_);
  not (_30754_, _30753_);
  and (_30755_, _30754_, _30145_);
  nor (_30756_, _30755_, _30731_);
  nor (_30757_, _30756_, _30752_);
  and (_30758_, _30731_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_30759_, _30738_, _17922_);
  not (_30760_, _30759_);
  and (_30761_, _30760_, _30061_);
  and (_30762_, _30761_, _30085_);
  and (_30763_, _30762_, _30082_);
  nor (_30764_, _30763_, _30731_);
  nor (_30765_, _30764_, _30758_);
  and (_30766_, _30731_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  or (_30767_, _30738_, _18424_);
  and (_30768_, _30767_, _29636_);
  and (_30769_, _30768_, _29669_);
  nand (_30770_, _30769_, _29548_);
  and (_30771_, _30770_, _30730_);
  nor (_30772_, _30771_, _30766_);
  and (_30773_, _30731_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_30774_, _30738_, _18249_);
  not (_30775_, _30774_);
  and (_30776_, _30775_, _29006_);
  and (_30777_, _30776_, _29199_);
  nor (_30778_, _30777_, _30731_);
  nor (_30779_, _30778_, _30773_);
  nor (_30780_, _30730_, _24361_);
  nor (_30781_, _30738_, _18794_);
  not (_30782_, _30781_);
  and (_30783_, _30782_, _28436_);
  and (_30784_, _30783_, _28433_);
  and (_30785_, _30784_, _28372_);
  not (_30786_, _30785_);
  and (_30787_, _30786_, _30730_);
  nor (_30788_, _30787_, _30780_);
  and (_30789_, _30788_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_30790_, _30789_, _30779_);
  and (_30791_, _30790_, _30772_);
  and (_30792_, _30791_, _30765_);
  and (_30793_, _30792_, _30757_);
  and (_30794_, _30793_, _30751_);
  and (_30795_, _30794_, _30744_);
  nor (_30796_, _30730_, _23681_);
  and (_30797_, _30796_, _30795_);
  nor (_30798_, _30796_, _30795_);
  nor (_30799_, _30798_, _30797_);
  and (_30800_, _30799_, _23451_);
  nor (_30801_, _30730_, _23725_);
  not (_30802_, _30801_);
  nor (_30803_, _30802_, _30800_);
  nor (_30804_, _30738_, _17192_);
  not (_30805_, _30804_);
  and (_30806_, _30805_, _26775_);
  and (_30807_, _30806_, _26600_);
  and (_30808_, _30807_, _27158_);
  and (_30809_, _30808_, _30730_);
  nor (_30810_, _30809_, _30803_);
  and (_35975_[7], _30810_, _35583_);
  not (_30811_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_30812_, _30788_, _30811_);
  nor (_30813_, _30788_, _30811_);
  nor (_30814_, _30813_, _30812_);
  and (_30815_, _30814_, _23451_);
  nor (_30816_, _30815_, _24372_);
  nor (_30817_, _30816_, _30730_);
  nor (_30818_, _30817_, _30787_);
  nand (_35975_[0], _30818_, _35583_);
  nor (_30819_, _30789_, _30779_);
  nor (_30820_, _30819_, _30790_);
  nor (_30821_, _30820_, _23440_);
  nor (_30822_, _30821_, _24448_);
  nor (_30823_, _30822_, _30730_);
  nor (_30824_, _30823_, _30778_);
  nand (_35975_[1], _30824_, _35583_);
  nor (_30825_, _30790_, _30772_);
  nor (_30826_, _30825_, _30791_);
  nor (_30827_, _30826_, _23440_);
  nor (_30828_, _30827_, _24580_);
  nor (_30829_, _30828_, _30730_);
  nor (_30830_, _30829_, _30771_);
  nand (_35975_[2], _30830_, _35583_);
  nor (_30831_, _30791_, _30765_);
  nor (_30832_, _30831_, _30792_);
  nor (_30833_, _30832_, _23440_);
  nor (_30834_, _30833_, _23900_);
  nor (_30835_, _30834_, _30730_);
  nor (_30836_, _30835_, _30764_);
  nor (_35975_[3], _30836_, rst);
  nor (_30837_, _30792_, _30757_);
  nor (_30838_, _30837_, _30793_);
  nor (_30839_, _30838_, _23440_);
  nor (_30840_, _30839_, _24075_);
  nor (_30841_, _30840_, _30730_);
  nor (_30842_, _30841_, _30756_);
  nor (_35975_[4], _30842_, rst);
  nor (_30843_, _30793_, _30751_);
  nor (_30844_, _30843_, _30794_);
  nor (_30845_, _30844_, _23440_);
  nor (_30846_, _30845_, _24196_);
  nor (_30847_, _30846_, _30730_);
  nor (_30848_, _30847_, _30750_);
  nor (_35975_[5], _30848_, rst);
  nor (_30849_, _30794_, _30744_);
  nor (_30850_, _30849_, _30795_);
  nor (_30851_, _30850_, _23440_);
  nor (_30852_, _30851_, _23483_);
  nor (_30853_, _30852_, _30730_);
  nor (_30854_, _30853_, _30743_);
  nor (_35975_[6], _30854_, rst);
  and (_30855_, _27518_, _24009_);
  and (_30856_, _30855_, _30101_);
  nand (_30857_, _30856_, _30727_);
  nor (_30858_, _30857_, _27441_);
  and (_30859_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _15093_);
  and (_30860_, _30859_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_30861_, _30857_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_30862_, _30861_, _30860_);
  or (_30863_, _30862_, _30858_);
  nor (_30864_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_30865_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_30866_, _30865_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30867_, _30866_, _30864_);
  nor (_30868_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not (_30869_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_30870_, _30869_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30871_, _30870_, _30868_);
  nor (_30872_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_30873_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_30874_, _30873_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30875_, _30874_, _30872_);
  not (_30876_, _30875_);
  nor (_30877_, _30876_, _27594_);
  nor (_30878_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not (_30879_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_30880_, _30879_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30881_, _30880_, _30878_);
  and (_30882_, _30881_, _30877_);
  nor (_30883_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not (_30884_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_30885_, _30884_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30886_, _30885_, _30883_);
  and (_30887_, _30886_, _30882_);
  and (_30888_, _30887_, _30871_);
  nor (_30889_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not (_30890_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_30891_, _30890_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30892_, _30891_, _30889_);
  and (_30893_, _30892_, _30888_);
  and (_30894_, _30893_, _30867_);
  nor (_30895_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_30896_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_30897_, _30896_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30898_, _30897_, _30895_);
  and (_30899_, _30898_, _30894_);
  nor (_30900_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_30901_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_30902_, _30901_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_30903_, _30902_, _30900_);
  nor (_30904_, _30903_, _30899_);
  and (_30905_, _30903_, _30899_);
  or (_30906_, _30905_, _30904_);
  nor (_30907_, _30906_, _27583_);
  not (_30908_, _30907_);
  and (_30909_, _20184_, _15159_);
  nor (_30910_, _17192_, _15877_);
  and (_30911_, _30910_, _26927_);
  and (_30912_, _30911_, _25261_);
  and (_30913_, _30912_, _25305_);
  and (_30914_, _30913_, _25921_);
  nor (_30915_, _30914_, _26949_);
  and (_30916_, _25866_, _15714_);
  nor (_30917_, _30916_, _30915_);
  and (_30918_, _27015_, _17192_);
  and (_30919_, _16541_, _15551_);
  and (_30920_, _16843_, _15877_);
  and (_30921_, _30920_, _30919_);
  and (_30922_, _30921_, _30918_);
  and (_30923_, _16680_, _15714_);
  and (_30924_, _30923_, _30922_);
  nor (_30925_, _30924_, _25866_);
  and (_30926_, _25866_, _16680_);
  nor (_30927_, _30926_, _30925_);
  and (_30928_, _30927_, _30917_);
  nor (_30929_, _25866_, _16051_);
  and (_30930_, _25866_, _16051_);
  nor (_30931_, _30930_, _30929_);
  and (_30932_, _30931_, _30928_);
  and (_30933_, _30932_, _27095_);
  nor (_30934_, _30932_, _27095_);
  nor (_30935_, _30934_, _30933_);
  and (_30936_, _30935_, _26862_);
  and (_30937_, _20494_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and (_30938_, _25866_, _27095_);
  nor (_30939_, _30938_, _27703_);
  nor (_30940_, _30939_, _27125_);
  nor (_30941_, _27867_, _17922_);
  nor (_30942_, _26796_, _17018_);
  or (_30943_, _30942_, _30941_);
  or (_30944_, _30943_, _30940_);
  nor (_30945_, _30944_, _30937_);
  not (_30946_, _30945_);
  nor (_30947_, _30946_, _30936_);
  not (_30948_, _30947_);
  nor (_30949_, _30948_, _30909_);
  and (_30950_, _30949_, _30908_);
  nand (_30951_, _30950_, _30860_);
  and (_30952_, _30951_, _35583_);
  and (_35967_[7], _30952_, _30863_);
  and (_30953_, _30855_, _30038_);
  and (_30954_, _30953_, _30727_);
  nor (_30955_, _30954_, _30860_);
  not (_30956_, _30955_);
  nand (_30957_, _30956_, _27441_);
  not (_30958_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand (_30959_, _30955_, _30958_);
  and (_30960_, _30959_, _35583_);
  and (_35968_[7], _30960_, _30957_);
  nor (_30961_, _30857_, _28556_);
  and (_30962_, _30857_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_30963_, _30962_, _30860_);
  or (_30964_, _30963_, _30961_);
  and (_30965_, _22795_, _20494_);
  not (_30966_, _30965_);
  and (_30967_, _30876_, _27594_);
  nor (_30968_, _30967_, _30877_);
  and (_30969_, _30968_, _26108_);
  nor (_30970_, _27703_, _27103_);
  not (_30971_, _30970_);
  nor (_30972_, _30971_, _27037_);
  nor (_30973_, _30972_, _25228_);
  and (_30974_, _30972_, _25228_);
  or (_30975_, _30974_, _30078_);
  nor (_30976_, _30975_, _30973_);
  nor (_30977_, _26796_, _15877_);
  and (_30978_, _19960_, _15159_);
  nor (_30979_, _27867_, _17563_);
  nor (_30980_, _27125_, _18794_);
  or (_30981_, _30980_, _30979_);
  or (_30982_, _30981_, _30978_);
  nor (_30983_, _30982_, _30977_);
  not (_30984_, _30983_);
  nor (_30985_, _30984_, _30976_);
  not (_30986_, _30985_);
  nor (_30987_, _30986_, _30969_);
  and (_30988_, _30987_, _30966_);
  nand (_30989_, _30988_, _30860_);
  and (_30990_, _30989_, _35583_);
  and (_35967_[0], _30990_, _30964_);
  nor (_30991_, _30857_, _29242_);
  and (_30992_, _30857_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_30993_, _30992_, _30860_);
  or (_30994_, _30993_, _30991_);
  nor (_30995_, _30881_, _30877_);
  nor (_30996_, _30995_, _30882_);
  and (_30997_, _30996_, _26108_);
  not (_30998_, _30997_);
  and (_30999_, _21786_, _20494_);
  and (_31000_, _30911_, _25866_);
  and (_31001_, _30918_, _15877_);
  and (_31002_, _31001_, _26949_);
  nor (_31003_, _31002_, _31000_);
  nor (_31004_, _31003_, _25261_);
  and (_31005_, _31003_, _25261_);
  nor (_31006_, _31005_, _31004_);
  nor (_31007_, _31006_, _30078_);
  nor (_31008_, _26796_, _16843_);
  and (_31009_, _19992_, _15159_);
  nor (_31010_, _27867_, _17388_);
  nor (_31011_, _27125_, _18249_);
  or (_31012_, _31011_, _31010_);
  or (_31013_, _31012_, _31009_);
  nor (_31014_, _31013_, _31008_);
  not (_31015_, _31014_);
  nor (_31016_, _31015_, _31007_);
  not (_31017_, _31016_);
  nor (_31018_, _31017_, _30999_);
  and (_31019_, _31018_, _30998_);
  nand (_31020_, _31019_, _30860_);
  and (_31021_, _31020_, _35583_);
  and (_35967_[1], _31021_, _30994_);
  nor (_31022_, _30857_, _29887_);
  and (_31023_, _30857_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_31024_, _31023_, _30860_);
  or (_31025_, _31024_, _31022_);
  nor (_31026_, _30886_, _30882_);
  nor (_31027_, _31026_, _30887_);
  and (_31028_, _31027_, _26108_);
  not (_31029_, _31028_);
  and (_31030_, _31001_, _16843_);
  and (_31031_, _31030_, _26949_);
  and (_31032_, _30912_, _25866_);
  nor (_31033_, _31032_, _31031_);
  and (_31034_, _31033_, _15551_);
  nor (_31035_, _31033_, _15551_);
  nor (_31036_, _31035_, _31034_);
  and (_31037_, _31036_, _26862_);
  not (_31038_, _31037_);
  nor (_31039_, _27125_, _18424_);
  and (_31040_, _20494_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_31041_, _31040_, _31039_);
  and (_31042_, _20024_, _15159_);
  nor (_31043_, _27867_, _16367_);
  nor (_31044_, _26796_, _15551_);
  or (_31045_, _31044_, _31043_);
  nor (_31046_, _31045_, _31042_);
  and (_31047_, _31046_, _31041_);
  and (_31048_, _31047_, _31038_);
  and (_31049_, _31048_, _31029_);
  nand (_31050_, _31049_, _30860_);
  and (_31051_, _31050_, _35583_);
  and (_35967_[2], _31051_, _31025_);
  nor (_31052_, _30857_, _30092_);
  and (_31053_, _30857_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_31054_, _31053_, _30860_);
  or (_31055_, _31054_, _31052_);
  nor (_31056_, _30887_, _30871_);
  nor (_31057_, _31056_, _30888_);
  and (_31058_, _31057_, _26108_);
  not (_31059_, _31058_);
  nor (_31060_, _30913_, _25921_);
  not (_31061_, _31060_);
  and (_31062_, _31061_, _30915_);
  and (_31063_, _31030_, _15551_);
  nor (_31064_, _31063_, _16541_);
  nor (_31065_, _31064_, _30922_);
  nor (_31066_, _31065_, _25866_);
  nor (_31067_, _31066_, _31062_);
  nor (_31068_, _31067_, _30078_);
  nor (_31069_, _26796_, _16541_);
  or (_31070_, _31069_, _27878_);
  nor (_31071_, _31070_, _31068_);
  and (_31072_, _20056_, _15159_);
  nor (_31073_, _27125_, _17922_);
  and (_31074_, _20494_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_31075_, _31074_, _31073_);
  nor (_31076_, _31075_, _31072_);
  and (_31077_, _31076_, _31071_);
  and (_31078_, _31077_, _31059_);
  nand (_31079_, _31078_, _30860_);
  and (_31080_, _31079_, _35583_);
  and (_35967_[3], _31080_, _31055_);
  nor (_31081_, _30857_, _30161_);
  and (_31082_, _30857_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_31083_, _31082_, _30860_);
  or (_31084_, _31083_, _31081_);
  nor (_31085_, _30892_, _30888_);
  not (_31086_, _31085_);
  nor (_31087_, _30893_, _27583_);
  and (_31088_, _31087_, _31086_);
  not (_31089_, _31088_);
  and (_31090_, _20088_, _15159_);
  nor (_31091_, _30922_, _25866_);
  nor (_31092_, _31091_, _30915_);
  nor (_31093_, _31092_, _24953_);
  and (_31094_, _31092_, _24953_);
  nor (_31095_, _31094_, _31093_);
  and (_31096_, _31095_, _26862_);
  and (_31097_, _20494_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_31098_, _25866_, _17574_);
  or (_31099_, _31098_, _27125_);
  nor (_31100_, _31099_, _30916_);
  nor (_31101_, _27867_, _18794_);
  nor (_31102_, _26796_, _15714_);
  or (_31103_, _31102_, _31101_);
  or (_31104_, _31103_, _31100_);
  nor (_31105_, _31104_, _31097_);
  not (_31106_, _31105_);
  nor (_31107_, _31106_, _31096_);
  not (_31108_, _31107_);
  nor (_31109_, _31108_, _31090_);
  and (_31110_, _31109_, _31089_);
  nand (_31111_, _31110_, _30860_);
  and (_31112_, _31111_, _35583_);
  and (_35967_[4], _31112_, _31084_);
  nor (_31113_, _30857_, _30236_);
  and (_31114_, _30857_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_31115_, _31114_, _30860_);
  or (_31116_, _31115_, _31113_);
  nor (_31117_, _30893_, _30867_);
  nor (_31118_, _31117_, _30894_);
  and (_31119_, _31118_, _26108_);
  not (_31120_, _31119_);
  and (_31121_, _20120_, _15159_);
  and (_31122_, _30922_, _15714_);
  nor (_31123_, _31122_, _25866_);
  not (_31124_, _31123_);
  and (_31125_, _31124_, _30917_);
  and (_31126_, _31125_, _16680_);
  nor (_31127_, _31125_, _16680_);
  nor (_31128_, _31127_, _31126_);
  nor (_31129_, _31128_, _30078_);
  and (_31130_, _20494_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_31131_, _25866_, _17399_);
  or (_31132_, _31131_, _27125_);
  nor (_31133_, _31132_, _30926_);
  nor (_31134_, _27867_, _18249_);
  nor (_31135_, _26796_, _16680_);
  or (_31136_, _31135_, _31134_);
  or (_31137_, _31136_, _31133_);
  nor (_31138_, _31137_, _31130_);
  not (_31139_, _31138_);
  nor (_31140_, _31139_, _31129_);
  not (_31141_, _31140_);
  nor (_31142_, _31141_, _31121_);
  and (_31143_, _31142_, _31120_);
  nand (_31144_, _31143_, _30860_);
  and (_31145_, _31144_, _35583_);
  and (_35967_[5], _31145_, _31116_);
  nor (_31146_, _30857_, _30309_);
  and (_31147_, _30857_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_31148_, _31147_, _30860_);
  or (_31149_, _31148_, _31146_);
  nor (_31150_, _30898_, _30894_);
  not (_31151_, _31150_);
  nor (_31152_, _30899_, _27583_);
  and (_31153_, _31152_, _31151_);
  not (_31154_, _31153_);
  and (_31155_, _20152_, _15159_);
  and (_31156_, _30928_, _16051_);
  nor (_31157_, _30928_, _16051_);
  nor (_31158_, _31157_, _31156_);
  nor (_31159_, _31158_, _30078_);
  nor (_31160_, _25866_, _16388_);
  not (_31161_, _31160_);
  nor (_31162_, _30930_, _27125_);
  and (_31163_, _31162_, _31161_);
  and (_31164_, _20494_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_31165_, _27867_, _18424_);
  nor (_31166_, _26796_, _16051_);
  or (_31167_, _31166_, _31165_);
  nor (_31168_, _31167_, _31164_);
  not (_31169_, _31168_);
  nor (_31170_, _31169_, _31163_);
  not (_31171_, _31170_);
  nor (_31172_, _31171_, _31159_);
  not (_31173_, _31172_);
  nor (_31174_, _31173_, _31155_);
  and (_31175_, _31174_, _31154_);
  nand (_31176_, _31175_, _30860_);
  and (_31177_, _31176_, _35583_);
  and (_35967_[6], _31177_, _31149_);
  nand (_31178_, _30956_, _28556_);
  not (_31179_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_31180_, _30955_, _31179_);
  and (_31181_, _31180_, _35583_);
  and (_35968_[0], _31181_, _31178_);
  nand (_31182_, _30956_, _29242_);
  not (_31183_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand (_31184_, _30955_, _31183_);
  and (_31185_, _31184_, _35583_);
  and (_35968_[1], _31185_, _31182_);
  nand (_31186_, _30956_, _29887_);
  not (_31187_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_31188_, _30955_, _31187_);
  and (_31189_, _31188_, _35583_);
  and (_35968_[2], _31189_, _31186_);
  nand (_31190_, _30956_, _30092_);
  or (_31191_, _30956_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_31192_, _31191_, _35583_);
  and (_35968_[3], _31192_, _31190_);
  nand (_31193_, _30956_, _30161_);
  or (_31194_, _30956_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_31195_, _31194_, _35583_);
  and (_35968_[4], _31195_, _31193_);
  nand (_31196_, _30956_, _30236_);
  or (_31197_, _30956_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_31198_, _31197_, _35583_);
  and (_35968_[5], _31198_, _31196_);
  nand (_31199_, _30956_, _30309_);
  or (_31200_, _30956_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_31201_, _31200_, _35583_);
  and (_35968_[6], _31201_, _31199_);
  and (_31202_, _24152_, _24284_);
  and (_31203_, _31202_, _23823_);
  and (_31204_, _31203_, _28166_);
  nor (_31205_, _30317_, _28062_);
  not (_31206_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_31207_, _28134_, _31206_);
  or (_31208_, _31207_, _31205_);
  and (_31209_, _31208_, _31204_);
  nor (_31210_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_31211_, _31210_);
  nand (_31212_, _31211_, _28062_);
  and (_31213_, _31210_, _31206_);
  nor (_31214_, _31213_, _31204_);
  and (_31215_, _31214_, _31212_);
  and (_31216_, _27518_, _24690_);
  and (_31217_, _31216_, _31203_);
  or (_31218_, _31217_, _31215_);
  or (_31219_, _31218_, _31209_);
  nand (_31220_, _31217_, _30808_);
  and (_31221_, _31220_, _31219_);
  and (_35973_[6], _31221_, _35583_);
  not (_31222_, _31217_);
  not (_31223_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand (_31224_, _31204_, _29329_);
  nand (_31225_, _31224_, _31223_);
  and (_31226_, _31225_, _31222_);
  or (_31227_, _31224_, _28654_);
  and (_31228_, _31227_, _31226_);
  nor (_31229_, _31222_, _30777_);
  or (_31230_, _31229_, _31228_);
  and (_35973_[0], _31230_, _35583_);
  not (_31231_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_31232_, _30038_, _31231_);
  or (_31233_, _31232_, _30039_);
  and (_31234_, _31233_, _31204_);
  or (_31235_, _20248_, _20216_);
  or (_31236_, _31235_, _20280_);
  or (_31237_, _31236_, _20322_);
  or (_31238_, _31237_, _20354_);
  or (_31239_, _31238_, _20397_);
  or (_31240_, _31239_, _20429_);
  or (_31241_, _31240_, _19897_);
  and (_31242_, _31241_, _15159_);
  or (_31243_, _27638_, _26030_);
  not (_31244_, _27627_);
  nand (_31245_, _31244_, _26030_);
  and (_31246_, _31245_, _24788_);
  and (_31247_, _31246_, _31243_);
  not (_31248_, _24810_);
  nand (_31249_, _26479_, _31248_);
  or (_31250_, _26479_, _24821_);
  and (_31251_, _26108_, _31250_);
  and (_31252_, _31251_, _31249_);
  and (_31253_, _30923_, _21688_);
  and (_31254_, _30921_, _20494_);
  nand (_31255_, _31254_, _31253_);
  nand (_31256_, _31255_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_31257_, _31256_, _31252_);
  or (_31258_, _31257_, _31247_);
  or (_31259_, _31258_, _31242_);
  nor (_31260_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor (_31261_, _31260_, _31204_);
  and (_31262_, _31261_, _31259_);
  or (_31263_, _31262_, _31234_);
  and (_31264_, _31263_, _31222_);
  and (_31265_, _31217_, _30770_);
  or (_31266_, _31265_, _31264_);
  and (_35973_[1], _31266_, _35583_);
  not (_31267_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand (_31268_, _31204_, _30101_);
  nand (_31269_, _31268_, _31267_);
  and (_31270_, _31269_, _31222_);
  or (_31271_, _31268_, _28654_);
  and (_31272_, _31271_, _31270_);
  nor (_31273_, _31222_, _30763_);
  or (_31274_, _31273_, _31272_);
  and (_35973_[2], _31274_, _35583_);
  and (_31275_, _30172_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_31276_, _31275_, _30176_);
  and (_31277_, _31276_, _31204_);
  nor (_31278_, _31222_, _30755_);
  not (_31279_, _31204_);
  or (_31280_, _31279_, _30173_);
  not (_31281_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_31282_, _31217_, _31281_);
  and (_31283_, _31282_, _31280_);
  or (_31284_, _31283_, _31278_);
  or (_31285_, _31284_, _31277_);
  and (_35973_[3], _31285_, _35583_);
  or (_31286_, _31279_, _30245_);
  and (_31287_, _31286_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_31288_, _31287_, _31217_);
  and (_31289_, _30251_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_31290_, _31289_, _30250_);
  and (_31291_, _31290_, _31204_);
  or (_31292_, _31291_, _31288_);
  nand (_31293_, _31217_, _30749_);
  and (_31294_, _31293_, _31292_);
  and (_35973_[4], _31294_, _35583_);
  or (_31295_, _30320_, _30054_);
  nand (_31296_, _31295_, _31204_);
  or (_31297_, _31296_, _30321_);
  and (_31298_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_31299_, _31298_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_31300_, _25976_, _24788_);
  and (_31301_, _26108_, _26370_);
  nand (_31302_, _26786_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_31303_, _31302_, _31298_);
  or (_31304_, _31303_, _31301_);
  or (_31305_, _31304_, _31300_);
  and (_31306_, _31305_, _31299_);
  or (_31307_, _31306_, _31204_);
  and (_31308_, _31307_, _31222_);
  and (_31309_, _31308_, _31297_);
  nor (_31310_, _31222_, _30742_);
  or (_31311_, _31310_, _31309_);
  and (_35973_[5], _31311_, _35583_);
  not (_31312_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_31313_, _30859_, _31312_);
  and (_31314_, _31313_, _30950_);
  nor (_31315_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_31316_, _31315_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_31317_, _24668_, _24009_);
  and (_31318_, _31317_, _30170_);
  and (_31319_, _24141_, _24295_);
  and (_31320_, _31319_, _23823_);
  and (_31321_, _31320_, _31318_);
  and (_31322_, _31321_, _27518_);
  nor (_31323_, _31322_, _31316_);
  nor (_31324_, _31323_, _27441_);
  not (_31325_, _31313_);
  and (_31326_, _28166_, _28082_);
  and (_31327_, _24141_, _24009_);
  and (_31328_, _31327_, _28072_);
  and (_31329_, _31328_, _31326_);
  and (_31330_, _31329_, _28134_);
  and (_31331_, _31330_, _28062_);
  not (_31332_, _31323_);
  nor (_31333_, _31330_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_31334_, _31333_, _31332_);
  or (_31335_, _31334_, _31331_);
  and (_31336_, _31335_, _31325_);
  not (_31337_, _31336_);
  nor (_31338_, _31337_, _31324_);
  nor (_31339_, _31338_, _31314_);
  and (_35965_[7], _31339_, _35583_);
  and (_31340_, _31313_, _30988_);
  nor (_31341_, _31323_, _28556_);
  and (_31342_, _31329_, _24690_);
  and (_31343_, _31342_, _28062_);
  nor (_31344_, _31342_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_31345_, _31344_, _31332_);
  or (_31346_, _31345_, _31343_);
  and (_31347_, _31346_, _31325_);
  not (_31348_, _31347_);
  nor (_31349_, _31348_, _31341_);
  nor (_31350_, _31349_, _31340_);
  and (_35965_[0], _31350_, _35583_);
  and (_31351_, _31313_, _31019_);
  nor (_31352_, _31323_, _29242_);
  and (_31353_, _31329_, _29329_);
  and (_31354_, _31353_, _28062_);
  nor (_31355_, _31353_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_31356_, _31355_, _31332_);
  or (_31357_, _31356_, _31354_);
  and (_31358_, _31357_, _31325_);
  not (_31359_, _31358_);
  nor (_31360_, _31359_, _31352_);
  nor (_31361_, _31360_, _31351_);
  and (_35965_[1], _31361_, _35583_);
  nor (_31362_, _31325_, _31049_);
  and (_31363_, _31332_, _29887_);
  not (_31364_, _31329_);
  not (_31365_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_31366_, _30038_, _31365_);
  nor (_31367_, _31366_, _30039_);
  nor (_31368_, _31367_, _31364_);
  nor (_31369_, _31329_, _31365_);
  nor (_31370_, _31369_, _31332_);
  not (_31371_, _31370_);
  nor (_31372_, _31371_, _31368_);
  nor (_31373_, _31372_, _31313_);
  not (_31374_, _31373_);
  nor (_31375_, _31374_, _31363_);
  nor (_31376_, _31375_, _31362_);
  nor (_35965_[2], _31376_, rst);
  nor (_31377_, _31325_, _31078_);
  and (_31378_, _31332_, _30092_);
  not (_31379_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_31380_, _30101_, _31379_);
  nor (_31381_, _31380_, _30102_);
  nor (_31382_, _31381_, _31364_);
  nor (_31383_, _31329_, _31379_);
  nor (_31384_, _31383_, _31332_);
  not (_31385_, _31384_);
  nor (_31386_, _31385_, _31382_);
  nor (_31387_, _31386_, _31313_);
  not (_31388_, _31387_);
  nor (_31389_, _31388_, _31378_);
  nor (_31390_, _31389_, _31377_);
  nor (_35965_[3], _31390_, rst);
  and (_31391_, _31313_, _31110_);
  nor (_31392_, _31323_, _30161_);
  and (_31393_, _31329_, _30171_);
  and (_31394_, _31393_, _28062_);
  nor (_31395_, _31393_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_31396_, _31395_, _31332_);
  or (_31397_, _31396_, _31394_);
  and (_31398_, _31397_, _31325_);
  not (_31399_, _31398_);
  nor (_31400_, _31399_, _31392_);
  nor (_31401_, _31400_, _31391_);
  and (_35965_[4], _31401_, _35583_);
  and (_31402_, _31313_, _31143_);
  nor (_31403_, _31323_, _30236_);
  and (_31404_, _31329_, _30249_);
  and (_31405_, _31404_, _28062_);
  nor (_31406_, _31404_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_31407_, _31406_, _31332_);
  or (_31408_, _31407_, _31405_);
  and (_31409_, _31408_, _31325_);
  not (_31410_, _31409_);
  nor (_31411_, _31410_, _31403_);
  nor (_31412_, _31411_, _31402_);
  and (_35965_[5], _31412_, _35583_);
  and (_31413_, _31313_, _31175_);
  nor (_31414_, _31323_, _30309_);
  and (_31415_, _31329_, _30320_);
  and (_31416_, _31415_, _28062_);
  nor (_31417_, _31415_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_31418_, _31417_, _31332_);
  or (_31419_, _31418_, _31416_);
  and (_31420_, _31419_, _31325_);
  not (_31421_, _31420_);
  nor (_31422_, _31421_, _31414_);
  nor (_31423_, _31422_, _31413_);
  and (_35965_[6], _31423_, _35583_);
  and (_31424_, _30728_, _28134_);
  nand (_31425_, _31424_, _28062_);
  or (_31426_, _31424_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_31427_, _31426_, _28166_);
  and (_31428_, _31427_, _31425_);
  and (_31429_, _30727_, _31318_);
  nand (_31430_, _31429_, _30808_);
  or (_31431_, _31429_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_31432_, _31431_, _27518_);
  and (_31433_, _31432_, _31430_);
  not (_31434_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_31435_, _27507_, _31434_);
  or (_31436_, _31435_, rst);
  or (_31437_, _31436_, _31433_);
  or (_35969_[7], _31437_, _31428_);
  and (_31438_, _31202_, _30726_);
  and (_31439_, _31438_, _28134_);
  nand (_31440_, _31439_, _28062_);
  or (_31441_, _31439_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_31442_, _31441_, _28166_);
  and (_31443_, _31442_, _31440_);
  and (_31444_, _31438_, _24690_);
  not (_31445_, _31444_);
  nor (_31446_, _31445_, _30808_);
  not (_31447_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_31448_, _31444_, _31447_);
  or (_31449_, _31448_, _31446_);
  and (_31450_, _31449_, _27518_);
  nor (_31451_, _27507_, _31447_);
  or (_31452_, _31451_, rst);
  or (_31453_, _31452_, _31450_);
  or (_35970_[7], _31453_, _31443_);
  and (_31454_, _24295_, _23670_);
  and (_31455_, _31454_, _31327_);
  and (_31456_, _31455_, _28082_);
  and (_31457_, _31456_, _28134_);
  nand (_31458_, _31457_, _28062_);
  or (_31459_, _31457_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_31460_, _31459_, _28166_);
  and (_31461_, _31460_, _31458_);
  and (_31462_, _31327_, _24701_);
  and (_31463_, _31462_, _30726_);
  not (_31464_, _31463_);
  nor (_31465_, _31464_, _30808_);
  not (_31466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_31467_, _31463_, _31466_);
  or (_31468_, _31467_, _31465_);
  and (_31469_, _31468_, _27518_);
  nor (_31470_, _27507_, _31466_);
  or (_31471_, _31470_, rst);
  or (_31472_, _31471_, _31469_);
  or (_35971_[7], _31472_, _31461_);
  and (_31473_, _31454_, _28093_);
  and (_31474_, _31473_, _28134_);
  nand (_31475_, _31474_, _28062_);
  or (_31476_, _31474_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_31477_, _31476_, _28166_);
  and (_31478_, _31477_, _31475_);
  and (_31479_, _30726_, _24712_);
  not (_31480_, _31479_);
  nor (_31481_, _31480_, _30808_);
  not (_31482_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_31483_, _31479_, _31482_);
  or (_31484_, _31483_, _31481_);
  and (_31485_, _31484_, _27518_);
  nor (_31486_, _27507_, _31482_);
  or (_31487_, _31486_, rst);
  or (_31488_, _31487_, _31485_);
  or (_35972_[7], _31488_, _31478_);
  not (_31489_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nor (_31490_, _31429_, _31489_);
  not (_31491_, _31429_);
  nor (_31492_, _31491_, _28062_);
  or (_31493_, _31492_, _31490_);
  and (_31494_, _31493_, _28166_);
  and (_31495_, _31429_, _30786_);
  or (_31496_, _31495_, _31490_);
  and (_31497_, _31496_, _27518_);
  nor (_31498_, _27507_, _31489_);
  or (_31499_, _31498_, rst);
  or (_31500_, _31499_, _31497_);
  or (_35969_[0], _31500_, _31494_);
  nand (_31501_, _30729_, _28062_);
  or (_31502_, _30729_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_31503_, _31502_, _28166_);
  and (_31504_, _31503_, _31501_);
  nand (_31505_, _31429_, _30777_);
  or (_31506_, _31429_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_31507_, _31506_, _27518_);
  and (_31508_, _31507_, _31505_);
  not (_31509_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_31510_, _27507_, _31509_);
  or (_31511_, _31510_, rst);
  or (_31512_, _31511_, _31508_);
  or (_35969_[1], _31512_, _31504_);
  not (_31513_, _30104_);
  nand (_31514_, _30728_, _31513_);
  and (_31515_, _31514_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_31516_, _24679_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_31517_, _31516_, _30039_);
  and (_31518_, _31517_, _30728_);
  or (_31519_, _31518_, _31515_);
  and (_31520_, _31519_, _28166_);
  or (_31521_, _31491_, _30770_);
  or (_31522_, _31429_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_31523_, _31522_, _27518_);
  and (_31524_, _31523_, _31521_);
  not (_31525_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_31526_, _27507_, _31525_);
  or (_31527_, _31526_, rst);
  or (_31528_, _31527_, _31524_);
  or (_35969_[2], _31528_, _31520_);
  nand (_31529_, _30728_, _24668_);
  and (_31530_, _31529_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_31531_, _31513_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_31532_, _31531_, _30102_);
  and (_31533_, _31532_, _30728_);
  or (_31534_, _31533_, _31530_);
  and (_31535_, _31534_, _28166_);
  nand (_31536_, _31429_, _30763_);
  or (_31537_, _31429_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_31538_, _31537_, _27518_);
  and (_31539_, _31538_, _31536_);
  not (_31540_, _27507_);
  and (_31541_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_31542_, _31541_, rst);
  or (_31543_, _31542_, _31539_);
  or (_35969_[3], _31543_, _31535_);
  and (_31544_, _30728_, _30171_);
  nand (_31545_, _31544_, _28062_);
  or (_31546_, _31544_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_31547_, _31546_, _28166_);
  and (_31548_, _31547_, _31545_);
  nand (_31549_, _31429_, _30755_);
  or (_31550_, _31429_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_31551_, _31550_, _27518_);
  and (_31552_, _31551_, _31549_);
  and (_31553_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_31554_, _31553_, rst);
  or (_31555_, _31554_, _31552_);
  or (_35969_[4], _31555_, _31548_);
  and (_31556_, _30728_, _30249_);
  nand (_31557_, _31556_, _28062_);
  or (_31558_, _31556_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_31559_, _31558_, _28166_);
  and (_31560_, _31559_, _31557_);
  nand (_31561_, _31429_, _30749_);
  or (_31562_, _31429_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_31563_, _31562_, _27518_);
  and (_31564_, _31563_, _31561_);
  and (_31565_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_31566_, _31565_, rst);
  or (_31567_, _31566_, _31564_);
  or (_35969_[5], _31567_, _31560_);
  nand (_31568_, _30728_, _30317_);
  and (_31569_, _31568_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  not (_31570_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_31571_, _28123_, _31570_);
  or (_31572_, _31571_, _30321_);
  and (_31573_, _31572_, _30728_);
  or (_31574_, _31573_, _31569_);
  and (_31575_, _31574_, _28166_);
  nand (_31576_, _31429_, _30742_);
  or (_31577_, _31429_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_31578_, _31577_, _27518_);
  and (_31579_, _31578_, _31576_);
  nor (_31580_, _27507_, _31570_);
  or (_31581_, _31580_, rst);
  or (_31582_, _31581_, _31579_);
  or (_35969_[6], _31582_, _31575_);
  nand (_31583_, _31444_, _28062_);
  or (_31584_, _31444_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_31585_, _31584_, _28166_);
  and (_31586_, _31585_, _31583_);
  and (_31587_, _31444_, _30786_);
  not (_31588_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nor (_31589_, _31444_, _31588_);
  or (_31590_, _31589_, _31587_);
  and (_31591_, _31590_, _27518_);
  nor (_31592_, _27507_, _31588_);
  or (_31593_, _31592_, rst);
  or (_31594_, _31593_, _31591_);
  or (_35970_[0], _31594_, _31586_);
  and (_31595_, _31438_, _29329_);
  nand (_31596_, _31595_, _28062_);
  or (_31597_, _31595_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_31598_, _31597_, _28166_);
  and (_31599_, _31598_, _31596_);
  nor (_31600_, _31445_, _30777_);
  not (_31601_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_31602_, _31444_, _31601_);
  or (_31603_, _31602_, _31600_);
  and (_31604_, _31603_, _27518_);
  nor (_31605_, _27507_, _31601_);
  or (_31606_, _31605_, rst);
  or (_31607_, _31606_, _31604_);
  or (_35970_[1], _31607_, _31599_);
  and (_31608_, _31438_, _30038_);
  nand (_31609_, _31608_, _28062_);
  or (_31610_, _31608_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_31611_, _31610_, _28166_);
  and (_31612_, _31611_, _31609_);
  and (_31613_, _31444_, _30770_);
  not (_31614_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_31615_, _31444_, _31614_);
  or (_31616_, _31615_, _31613_);
  and (_31617_, _31616_, _27518_);
  nor (_31618_, _27507_, _31614_);
  or (_31619_, _31618_, rst);
  or (_31620_, _31619_, _31617_);
  or (_35970_[2], _31620_, _31612_);
  and (_31621_, _31438_, _30101_);
  nand (_31622_, _31621_, _28062_);
  or (_31623_, _31621_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_31624_, _31623_, _28166_);
  and (_31625_, _31624_, _31622_);
  nor (_31626_, _31445_, _30763_);
  and (_31627_, _31445_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_31628_, _31627_, _31626_);
  and (_31629_, _31628_, _27518_);
  and (_31630_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_31631_, _31630_, rst);
  or (_31632_, _31631_, _31629_);
  or (_35970_[3], _31632_, _31625_);
  and (_31633_, _31438_, _30171_);
  nand (_31634_, _31633_, _28062_);
  or (_31635_, _31633_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_31636_, _31635_, _28166_);
  and (_31637_, _31636_, _31634_);
  nor (_31638_, _31445_, _30755_);
  and (_31639_, _31445_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_31640_, _31639_, _31638_);
  and (_31641_, _31640_, _27518_);
  and (_31642_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_31643_, _31642_, rst);
  or (_31644_, _31643_, _31641_);
  or (_35970_[4], _31644_, _31637_);
  and (_31645_, _31438_, _30249_);
  nand (_31646_, _31645_, _28062_);
  or (_31647_, _31645_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_31648_, _31647_, _28166_);
  and (_31649_, _31648_, _31646_);
  nor (_31650_, _31445_, _30749_);
  and (_31651_, _31445_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_31652_, _31651_, _31650_);
  and (_31653_, _31652_, _27518_);
  and (_31654_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_31655_, _31654_, rst);
  or (_31656_, _31655_, _31653_);
  or (_35970_[5], _31656_, _31649_);
  and (_31657_, _31438_, _30320_);
  nand (_31658_, _31657_, _28062_);
  or (_31659_, _31657_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_31660_, _31659_, _28166_);
  and (_31661_, _31660_, _31658_);
  nor (_31662_, _31445_, _30742_);
  not (_31663_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_31664_, _31444_, _31663_);
  or (_31665_, _31664_, _31662_);
  and (_31666_, _31665_, _27518_);
  nor (_31667_, _27507_, _31663_);
  or (_31668_, _31667_, rst);
  or (_31669_, _31668_, _31666_);
  or (_35970_[6], _31669_, _31661_);
  and (_31670_, _31456_, _24690_);
  nand (_31671_, _31670_, _28062_);
  or (_31672_, _31670_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_31673_, _31672_, _28166_);
  and (_31674_, _31673_, _31671_);
  nor (_31675_, _31464_, _30785_);
  not (_31676_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nor (_31677_, _31463_, _31676_);
  or (_31678_, _31677_, _31675_);
  and (_31679_, _31678_, _27518_);
  nor (_31680_, _27507_, _31676_);
  or (_31681_, _31680_, rst);
  or (_31682_, _31681_, _31679_);
  or (_35971_[0], _31682_, _31674_);
  and (_31683_, _31456_, _29329_);
  nand (_31684_, _31683_, _28062_);
  or (_31685_, _31683_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_31686_, _31685_, _28166_);
  and (_31687_, _31686_, _31684_);
  nor (_31688_, _31464_, _30777_);
  not (_31689_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_31690_, _31463_, _31689_);
  or (_31691_, _31690_, _31688_);
  and (_31692_, _31691_, _27518_);
  nor (_31693_, _27507_, _31689_);
  or (_31694_, _31693_, rst);
  or (_31695_, _31694_, _31692_);
  or (_35971_[1], _31695_, _31687_);
  and (_31696_, _31456_, _30038_);
  nand (_31697_, _31696_, _28062_);
  or (_31698_, _31696_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_31699_, _31698_, _28166_);
  and (_31700_, _31699_, _31697_);
  and (_31701_, _31463_, _30770_);
  not (_31702_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_31703_, _31463_, _31702_);
  or (_31704_, _31703_, _31701_);
  and (_31705_, _31704_, _27518_);
  nor (_31706_, _27507_, _31702_);
  or (_31707_, _31706_, rst);
  or (_31708_, _31707_, _31705_);
  or (_35971_[2], _31708_, _31700_);
  and (_31709_, _31456_, _30101_);
  nand (_31710_, _31709_, _28062_);
  or (_31711_, _31709_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_31712_, _31711_, _28166_);
  and (_31713_, _31712_, _31710_);
  nor (_31714_, _31464_, _30763_);
  and (_31715_, _31464_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_31716_, _31715_, _31714_);
  and (_31717_, _31716_, _27518_);
  and (_31718_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_31719_, _31718_, rst);
  or (_31720_, _31719_, _31717_);
  or (_35971_[3], _31720_, _31713_);
  and (_31721_, _31456_, _30171_);
  nand (_31722_, _31721_, _28062_);
  or (_31723_, _31721_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_31724_, _31723_, _28166_);
  and (_31725_, _31724_, _31722_);
  nor (_31726_, _31464_, _30755_);
  and (_31727_, _31464_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_31728_, _31727_, _31726_);
  and (_31729_, _31728_, _27518_);
  and (_31730_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_31731_, _31730_, rst);
  or (_31732_, _31731_, _31729_);
  or (_35971_[4], _31732_, _31725_);
  and (_31733_, _31456_, _30249_);
  nand (_31734_, _31733_, _28062_);
  or (_31735_, _31733_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_31736_, _31735_, _28166_);
  and (_31737_, _31736_, _31734_);
  nor (_31738_, _31464_, _30749_);
  and (_31739_, _31464_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_31740_, _31739_, _31738_);
  and (_31741_, _31740_, _27518_);
  and (_31742_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_31743_, _31742_, rst);
  or (_31744_, _31743_, _31741_);
  or (_35971_[5], _31744_, _31737_);
  and (_31745_, _31456_, _30320_);
  nand (_31746_, _31745_, _28062_);
  or (_31747_, _31745_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_31748_, _31747_, _28166_);
  and (_31749_, _31748_, _31746_);
  nor (_31750_, _31464_, _30742_);
  not (_31751_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_31752_, _31463_, _31751_);
  or (_31753_, _31752_, _31750_);
  and (_31754_, _31753_, _27518_);
  nor (_31755_, _27507_, _31751_);
  or (_31756_, _31755_, rst);
  or (_31757_, _31756_, _31754_);
  or (_35971_[6], _31757_, _31749_);
  and (_31758_, _31473_, _24690_);
  nand (_31759_, _31758_, _28062_);
  or (_31760_, _31758_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_31761_, _31760_, _28166_);
  and (_31762_, _31761_, _31759_);
  nor (_31763_, _31480_, _30785_);
  not (_31764_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_31765_, _31479_, _31764_);
  or (_31766_, _31765_, _31763_);
  and (_31767_, _31766_, _27518_);
  nor (_31768_, _27507_, _31764_);
  or (_31769_, _31768_, rst);
  or (_31770_, _31769_, _31767_);
  or (_35972_[0], _31770_, _31762_);
  and (_31771_, _31473_, _29329_);
  nand (_31772_, _31771_, _28062_);
  or (_31773_, _31771_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_31774_, _31773_, _28166_);
  and (_31775_, _31774_, _31772_);
  nor (_31776_, _31480_, _30777_);
  not (_31777_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_31778_, _31479_, _31777_);
  or (_31779_, _31778_, _31776_);
  and (_31780_, _31779_, _27518_);
  nor (_31781_, _27507_, _31777_);
  or (_31782_, _31781_, rst);
  or (_31783_, _31782_, _31780_);
  or (_35972_[1], _31783_, _31775_);
  and (_31784_, _31473_, _30038_);
  nand (_31785_, _31784_, _28062_);
  or (_31786_, _31784_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_31787_, _31786_, _28166_);
  and (_31788_, _31787_, _31785_);
  and (_31789_, _31479_, _30770_);
  not (_31790_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_31791_, _31479_, _31790_);
  or (_31792_, _31791_, _31789_);
  and (_31793_, _31792_, _27518_);
  nor (_31794_, _27507_, _31790_);
  or (_31795_, _31794_, rst);
  or (_31796_, _31795_, _31793_);
  or (_35972_[2], _31796_, _31788_);
  and (_31797_, _31473_, _30101_);
  nand (_31798_, _31797_, _28062_);
  or (_31799_, _31797_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_31800_, _31799_, _28166_);
  and (_31801_, _31800_, _31798_);
  nor (_31802_, _31480_, _30763_);
  and (_31803_, _31480_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31804_, _31803_, _31802_);
  and (_31805_, _31804_, _27518_);
  and (_31806_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_31807_, _31806_, rst);
  or (_31808_, _31807_, _31805_);
  or (_35972_[3], _31808_, _31801_);
  and (_31809_, _31473_, _30171_);
  nand (_31810_, _31809_, _28062_);
  or (_31811_, _31809_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_31812_, _31811_, _28166_);
  and (_31813_, _31812_, _31810_);
  nor (_31814_, _31480_, _30755_);
  and (_31815_, _31480_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31816_, _31815_, _31814_);
  and (_31817_, _31816_, _27518_);
  and (_31818_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_31819_, _31818_, rst);
  or (_31820_, _31819_, _31817_);
  or (_35972_[4], _31820_, _31813_);
  and (_31821_, _31473_, _30249_);
  nand (_31822_, _31821_, _28062_);
  or (_31823_, _31821_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_31824_, _31823_, _28166_);
  and (_31825_, _31824_, _31822_);
  nor (_31826_, _31480_, _30749_);
  and (_31827_, _31480_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_31828_, _31827_, _31826_);
  and (_31829_, _31828_, _27518_);
  and (_31830_, _31540_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_31831_, _31830_, rst);
  or (_31832_, _31831_, _31829_);
  or (_35972_[5], _31832_, _31825_);
  and (_31833_, _31473_, _30320_);
  nand (_31834_, _31833_, _28062_);
  or (_31835_, _31833_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_31836_, _31835_, _28166_);
  and (_31837_, _31836_, _31834_);
  nor (_31838_, _31480_, _30742_);
  not (_31839_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_31840_, _31479_, _31839_);
  or (_31841_, _31840_, _31838_);
  and (_31842_, _31841_, _27518_);
  nor (_31843_, _27507_, _31839_);
  or (_31844_, _31843_, rst);
  or (_31845_, _31844_, _31842_);
  or (_35972_[6], _31845_, _31837_);
  nor (_31846_, _23812_, _23429_);
  nor (_31847_, _31846_, _27496_);
  not (_31848_, _31847_);
  and (_31849_, _23812_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_31850_, _31849_, _24020_);
  nor (_31851_, _24416_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_31852_, _31851_, _31850_);
  not (_31853_, _31852_);
  and (_31854_, _30674_, _30603_);
  nor (_31855_, _30630_, _30619_);
  nor (_31856_, _30646_, _30634_);
  and (_31857_, _31856_, _30628_);
  and (_31858_, _31857_, _31855_);
  not (_31859_, _30642_);
  and (_31860_, _30663_, _31859_);
  and (_31861_, _31860_, _30675_);
  and (_31862_, _31861_, _31858_);
  nor (_31863_, _31862_, _30331_);
  nor (_31864_, _31863_, _31854_);
  not (_31865_, _31864_);
  not (_31866_, _30611_);
  and (_31867_, _30706_, _31866_);
  and (_31868_, _31867_, _30722_);
  nor (_31869_, _30544_, _24416_);
  and (_31870_, _30544_, _24416_);
  nor (_31871_, _31870_, _31869_);
  not (_31872_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_31873_, _24679_, _31872_);
  and (_31874_, _31873_, _31847_);
  not (_31875_, _31874_);
  nor (_31876_, _31875_, _31871_);
  nor (_31877_, _31217_, _31267_);
  nor (_31878_, _31877_, _31273_);
  nor (_31879_, _31878_, _24020_);
  and (_31880_, _31878_, _24020_);
  nor (_31881_, _31880_, _31879_);
  and (_31882_, _31881_, _31876_);
  and (_31883_, _31882_, _30786_);
  nor (_31884_, _31849_, _24020_);
  and (_31885_, _31849_, _23670_);
  nor (_31886_, _31885_, _31884_);
  and (_31887_, _31886_, _31878_);
  not (_31888_, _31887_);
  nor (_31889_, _31886_, _31878_);
  or (_31890_, _31852_, _30544_);
  nand (_31891_, _31852_, _30544_);
  and (_31892_, _31891_, _31890_);
  not (_31893_, _31892_);
  and (_31894_, _31849_, _24295_);
  nor (_31895_, _24668_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_31896_, _31895_, _31894_);
  not (_31897_, _24141_);
  and (_31898_, _31849_, _31897_);
  nor (_31899_, _24547_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_31900_, _31899_, _31898_);
  and (_31901_, _31900_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and (_31902_, _31901_, _31896_);
  and (_31903_, _31902_, _31893_);
  not (_31904_, _31903_);
  nor (_31905_, _31904_, _31889_);
  and (_31906_, _31905_, _31888_);
  not (_31907_, _31906_);
  and (_31908_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _25503_);
  and (_31909_, _31908_, _25568_);
  nand (_31910_, _31909_, _28062_);
  not (_31911_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand (_31912_, _30785_, _31911_);
  or (_31913_, _15769_, _31911_);
  and (_31914_, _31913_, _31912_);
  or (_31915_, _31914_, _31909_);
  and (_31916_, _31915_, _31910_);
  or (_31917_, _31916_, _31907_);
  not (_31918_, _31882_);
  and (_31919_, _31878_, _30544_);
  and (_31920_, _31919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_31921_, _31878_, _30574_);
  and (_31922_, _31921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  or (_31923_, _31922_, _31920_);
  nor (_31924_, _31878_, _30544_);
  and (_31925_, _31924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_31926_, _31878_, _30574_);
  and (_31927_, _31926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_31928_, _31927_, _31925_);
  or (_31929_, _31928_, _31923_);
  or (_31930_, _31929_, _31906_);
  and (_31931_, _31930_, _31918_);
  and (_31932_, _31931_, _31917_);
  or (_31933_, _31932_, _31883_);
  and (_31934_, _31933_, _31868_);
  not (_31935_, _31934_);
  and (_31936_, _30722_, _30707_);
  not (_31937_, _30818_);
  and (_31938_, _31937_, _31936_);
  not (_31939_, _31938_);
  and (_31940_, _30722_, _30611_);
  and (_31941_, _31940_, _30706_);
  and (_31942_, _31941_, _30574_);
  nor (_31943_, _30706_, _31866_);
  and (_31944_, _31943_, _30722_);
  not (_31945_, _30335_);
  and (_31946_, _31945_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and (_31947_, _30426_, _30335_);
  not (_31948_, _31947_);
  and (_31949_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_31950_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_31951_, _31950_, _31949_);
  and (_31952_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_31953_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_31954_, _31953_, _31952_);
  and (_31955_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_31956_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_31957_, _31956_, _31955_);
  and (_31958_, _31957_, _31954_);
  and (_31959_, _31958_, _31951_);
  nor (_31960_, _31959_, _31948_);
  nor (_31961_, _31960_, _31946_);
  not (_31962_, _31961_);
  and (_31963_, _31962_, _31944_);
  nor (_31964_, _31963_, _31942_);
  and (_31965_, _31964_, _31939_);
  and (_31966_, _31965_, _31935_);
  nor (_31967_, _31966_, _31865_);
  and (_31968_, _30588_, _30672_);
  nor (_31969_, _30698_, _31968_);
  nor (_31970_, _31969_, _30694_);
  not (_31971_, _30661_);
  and (_31972_, _30695_, _30422_);
  and (_31973_, _31972_, _30588_);
  nor (_31974_, _31973_, _30619_);
  and (_31975_, _31974_, _31971_);
  and (_31976_, _31975_, _31859_);
  and (_31977_, _31972_, _30548_);
  not (_31978_, _31977_);
  and (_31979_, _31978_, _31969_);
  not (_31980_, _30697_);
  and (_31981_, _30593_, _30555_);
  and (_31982_, _31981_, _30548_);
  nor (_31983_, _31982_, _30625_);
  and (_31984_, _31983_, _31980_);
  and (_31985_, _31984_, _31979_);
  and (_31986_, _31985_, _31976_);
  and (_31987_, _31986_, _31856_);
  nor (_31988_, _31987_, _30331_);
  nor (_31989_, _31988_, _31970_);
  not (_31990_, _16909_);
  not (_31991_, _25591_);
  and (_31992_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and (_31993_, _31992_, _31991_);
  nor (_31994_, _31993_, _31908_);
  nor (_31995_, _31994_, _31990_);
  and (_31996_, _31992_, _25591_);
  and (_31997_, _31996_, _28654_);
  nor (_31998_, _30808_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_31999_, _31998_, _31997_);
  nor (_32000_, _31999_, _31995_);
  and (_32001_, _32000_, _31906_);
  and (_32002_, _31926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_32003_, _31921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_32004_, _32003_, _32002_);
  and (_32005_, _31919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_32006_, _31924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor (_32007_, _32006_, _32005_);
  and (_32008_, _32007_, _32004_);
  and (_32009_, _32008_, _31907_);
  nor (_32010_, _32009_, _32001_);
  nor (_32011_, _32010_, _31882_);
  and (_32012_, _31882_, _30808_);
  nor (_32013_, _32012_, _32011_);
  and (_32014_, _32013_, _31868_);
  not (_32015_, _32014_);
  not (_32016_, _30722_);
  and (_32017_, _31945_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and (_32018_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_32019_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_32020_, _32019_, _32018_);
  and (_32021_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_32022_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_32023_, _32022_, _32021_);
  and (_32024_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_32025_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_32026_, _32025_, _32024_);
  and (_32027_, _32026_, _32023_);
  and (_32028_, _32027_, _32020_);
  nor (_32029_, _32028_, _31948_);
  nor (_32030_, _32029_, _32017_);
  not (_32031_, _32030_);
  and (_32032_, _32031_, _31943_);
  nor (_32033_, _32032_, _32016_);
  nand (_32034_, _30810_, _30707_);
  and (_32035_, _32034_, _32033_);
  and (_32036_, _32035_, _32015_);
  not (_32037_, _32036_);
  nor (_32038_, _32037_, _31989_);
  not (_32039_, _30763_);
  and (_32040_, _31882_, _32039_);
  and (_32041_, _31908_, _25591_);
  and (_32042_, _32041_, _28654_);
  nor (_32043_, _30763_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32044_, _31908_, _31991_);
  or (_32045_, _32044_, _31992_);
  and (_32046_, _32045_, _16432_);
  or (_32047_, _32046_, _32043_);
  or (_32048_, _32047_, _32042_);
  or (_32049_, _32048_, _31907_);
  and (_32050_, _31921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_32051_, _31926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_32052_, _32051_, _32050_);
  and (_32053_, _31924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_32054_, _31919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_32055_, _32054_, _32053_);
  or (_32056_, _32055_, _32052_);
  or (_32057_, _32056_, _31906_);
  and (_32058_, _32057_, _31918_);
  and (_32059_, _32058_, _32049_);
  or (_32060_, _32059_, _32040_);
  and (_32061_, _32060_, _31868_);
  not (_32062_, _32061_);
  not (_32063_, _30836_);
  and (_32064_, _32063_, _31936_);
  not (_32065_, _32064_);
  not (_32066_, _31878_);
  and (_32067_, _31941_, _32066_);
  and (_32068_, _31945_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and (_32069_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_32070_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_32071_, _32070_, _32069_);
  and (_32072_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_32073_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_32074_, _32073_, _32072_);
  and (_32075_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_32076_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_32077_, _32076_, _32075_);
  and (_32078_, _32077_, _32074_);
  and (_32079_, _32078_, _32071_);
  nor (_32080_, _32079_, _31948_);
  nor (_32081_, _32080_, _32068_);
  not (_32082_, _32081_);
  and (_32083_, _32082_, _31944_);
  nor (_32084_, _32083_, _32067_);
  and (_32085_, _32084_, _32065_);
  and (_32086_, _32085_, _32062_);
  not (_32087_, _32086_);
  and (_32088_, _32087_, _32038_);
  nor (_32089_, _32088_, _31967_);
  and (_32090_, _32089_, _31853_);
  nor (_32091_, _32090_, _31848_);
  not (_32092_, _31896_);
  and (_32093_, _31882_, _30770_);
  nand (_32094_, _31908_, _25525_);
  nor (_32095_, _32094_, _28062_);
  and (_32096_, _30770_, _31911_);
  nor (_32097_, _32041_, _31992_);
  nand (_32098_, _31908_, _25613_);
  nand (_32099_, _32098_, _32097_);
  and (_32100_, _32099_, _15409_);
  or (_32101_, _32100_, _32096_);
  or (_32102_, _32101_, _32095_);
  or (_32103_, _32102_, _31907_);
  and (_32104_, _31919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_32105_, _31921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_32106_, _32105_, _32104_);
  and (_32107_, _31924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_32108_, _31926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_32109_, _32108_, _32107_);
  or (_32110_, _32109_, _32106_);
  or (_32111_, _32110_, _31906_);
  and (_32112_, _32111_, _31918_);
  and (_32113_, _32112_, _32103_);
  or (_32114_, _32113_, _32093_);
  and (_32115_, _32114_, _31868_);
  not (_32116_, _32115_);
  not (_32117_, _30830_);
  and (_32118_, _32117_, _31936_);
  not (_32119_, _32118_);
  and (_32120_, _31941_, _30613_);
  and (_32121_, _31945_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and (_32122_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_32123_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_32124_, _32123_, _32122_);
  and (_32125_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_32126_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_32127_, _32126_, _32125_);
  and (_32128_, _32127_, _32124_);
  and (_32129_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_32130_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_32131_, _32130_, _32129_);
  and (_32132_, _32131_, _32128_);
  nor (_32133_, _32132_, _31948_);
  nor (_32134_, _32133_, _32121_);
  not (_32135_, _32134_);
  and (_32136_, _32135_, _31944_);
  nor (_32137_, _32136_, _32120_);
  and (_32138_, _32137_, _32119_);
  and (_32139_, _32138_, _32116_);
  nor (_32140_, _32139_, _31865_);
  not (_32141_, _31868_);
  nor (_32142_, _31918_, _30749_);
  and (_32143_, _25624_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_32144_, _32143_);
  and (_32145_, _16585_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32146_, _32145_, _32144_);
  and (_32147_, _31992_, _25624_);
  and (_32148_, _32147_, _28654_);
  nor (_32149_, _30749_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_32150_, _32149_, _32148_);
  nor (_32151_, _32150_, _32146_);
  and (_32152_, _32151_, _31906_);
  and (_32153_, _31919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_32154_, _31921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_32155_, _32154_, _32153_);
  and (_32156_, _31924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_32157_, _31926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_32158_, _32157_, _32156_);
  and (_32159_, _32158_, _32155_);
  and (_32160_, _32159_, _31907_);
  nor (_32161_, _32160_, _31882_);
  not (_32162_, _32161_);
  nor (_32163_, _32162_, _32152_);
  nor (_32164_, _32163_, _32142_);
  nor (_32165_, _32164_, _32141_);
  not (_32166_, _32165_);
  not (_32167_, _31943_);
  nor (_32168_, _31867_, _30722_);
  and (_32169_, _32168_, _32167_);
  not (_32170_, _32169_);
  not (_32171_, _30848_);
  and (_32172_, _32171_, _31936_);
  and (_32173_, _31945_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and (_32174_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_32175_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_32176_, _32175_, _32174_);
  and (_32177_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_32178_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_32179_, _32178_, _32177_);
  and (_32180_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_32181_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_32182_, _32181_, _32180_);
  and (_32183_, _32182_, _32179_);
  and (_32184_, _32183_, _32176_);
  nor (_32185_, _32184_, _31948_);
  nor (_32186_, _32185_, _32173_);
  not (_32187_, _32186_);
  and (_32188_, _32187_, _31944_);
  nor (_32189_, _32188_, _32172_);
  and (_32190_, _32189_, _32170_);
  and (_32191_, _32190_, _32166_);
  not (_32192_, _32191_);
  and (_32193_, _32038_, _32192_);
  nor (_32194_, _32193_, _32140_);
  and (_32195_, _32194_, _32092_);
  nor (_32196_, _32089_, _31853_);
  nor (_32197_, _32196_, _32195_);
  and (_32198_, _32197_, _32091_);
  and (_32199_, _31867_, _32016_);
  not (_32200_, _30824_);
  and (_32201_, _32200_, _31936_);
  nor (_32202_, _32201_, _32199_);
  and (_32203_, _31941_, _30545_);
  not (_32204_, _16734_);
  and (_32205_, _31908_, _25514_);
  not (_32206_, _32205_);
  and (_32207_, _32097_, _32206_);
  nor (_32208_, _32207_, _32204_);
  and (_32209_, _31908_, _25624_);
  and (_32210_, _32209_, _28654_);
  nor (_32211_, _30777_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_32212_, _32211_, _32210_);
  nor (_32213_, _32212_, _32208_);
  and (_32214_, _32213_, _31906_);
  and (_32215_, _31926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_32216_, _31921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_32217_, _32216_, _32215_);
  and (_32218_, _31924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_32219_, _31919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_32220_, _32219_, _32218_);
  and (_32221_, _32220_, _32217_);
  and (_32222_, _32221_, _31907_);
  nor (_32223_, _32222_, _32214_);
  nor (_32224_, _32223_, _31882_);
  and (_32225_, _31882_, _30777_);
  nor (_32226_, _32225_, _32224_);
  and (_32227_, _32226_, _31868_);
  and (_32228_, _31945_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and (_32229_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_32230_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_32231_, _32230_, _32229_);
  and (_32232_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_32233_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_32234_, _32233_, _32232_);
  and (_32235_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_32236_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_32237_, _32236_, _32235_);
  and (_32238_, _32237_, _32234_);
  and (_32239_, _32238_, _32231_);
  nor (_32240_, _32239_, _31948_);
  nor (_32241_, _32240_, _32228_);
  not (_32242_, _32241_);
  and (_32243_, _32242_, _31944_);
  or (_32244_, _32243_, _32227_);
  nor (_32245_, _32244_, _32203_);
  and (_32246_, _32245_, _32202_);
  nor (_32247_, _32246_, _31865_);
  not (_32248_, _30755_);
  and (_32249_, _31882_, _32248_);
  and (_32250_, _25568_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_32251_, _32250_);
  and (_32252_, _15605_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32253_, _32252_, _32251_);
  and (_32254_, _31992_, _25568_);
  and (_32255_, _32254_, _28654_);
  nor (_32256_, _30755_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or (_32257_, _32256_, _32255_);
  nor (_32258_, _32257_, _32253_);
  and (_32259_, _32258_, _31906_);
  and (_32260_, _31921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_32261_, _31926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_32262_, _32261_, _32260_);
  and (_32263_, _31924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_32264_, _31919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_32265_, _32264_, _32263_);
  and (_32266_, _32265_, _32262_);
  and (_32267_, _32266_, _31907_);
  nor (_32268_, _32267_, _31882_);
  not (_32269_, _32268_);
  nor (_32270_, _32269_, _32259_);
  nor (_32271_, _32270_, _32249_);
  nor (_32272_, _32271_, _32141_);
  not (_32273_, _32272_);
  not (_32274_, _30842_);
  and (_32275_, _32274_, _31936_);
  not (_32276_, _32275_);
  and (_32277_, _31945_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and (_32278_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_32279_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_32280_, _32279_, _32278_);
  and (_32281_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_32282_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_32283_, _32282_, _32281_);
  and (_32284_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_32285_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_32286_, _32285_, _32284_);
  and (_32287_, _32286_, _32283_);
  and (_32288_, _32287_, _32280_);
  nor (_32289_, _32288_, _31948_);
  nor (_32290_, _32289_, _32277_);
  not (_32291_, _32290_);
  and (_32292_, _32291_, _31944_);
  nor (_32293_, _31282_, _31278_);
  not (_32294_, _32293_);
  and (_32295_, _32294_, _31941_);
  and (_32296_, _32016_, _30611_);
  or (_32297_, _32296_, _32295_);
  nor (_32298_, _32297_, _32292_);
  and (_32299_, _32298_, _32276_);
  and (_32300_, _32299_, _32273_);
  not (_32301_, _32300_);
  and (_32302_, _32301_, _32038_);
  nor (_32303_, _32302_, _32247_);
  nand (_32304_, _32303_, _31900_);
  or (_32305_, _32303_, _31900_);
  and (_32306_, _32305_, _32304_);
  not (_32307_, _32306_);
  nor (_32308_, _32194_, _32092_);
  not (_32309_, _32308_);
  not (_32310_, _31886_);
  and (_32311_, _32036_, _31865_);
  nor (_32312_, _32087_, _32311_);
  not (_32313_, _30742_);
  and (_32314_, _31882_, _32313_);
  and (_32315_, _31926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_32316_, _31921_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_32317_, _32316_, _32315_);
  and (_32318_, _31924_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_32319_, _31919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_32320_, _32319_, _32318_);
  and (_32321_, _32320_, _32317_);
  and (_32322_, _32321_, _31907_);
  nor (_32323_, _30742_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32324_, _31992_, _25525_);
  and (_32325_, _32324_, _28654_);
  and (_32326_, _25525_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_32327_, _32326_);
  and (_32328_, _15943_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and (_32329_, _32328_, _32327_);
  or (_32330_, _32329_, _32325_);
  nor (_32331_, _32330_, _32323_);
  and (_32332_, _32331_, _31906_);
  or (_32333_, _32332_, _31882_);
  nor (_32334_, _32333_, _32322_);
  nor (_32335_, _32334_, _32314_);
  nor (_32336_, _32335_, _32141_);
  not (_32337_, _30854_);
  and (_32338_, _32337_, _31936_);
  and (_32339_, _31945_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and (_32340_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_32341_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_32342_, _32341_, _32340_);
  and (_32343_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_32344_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_32345_, _32344_, _32343_);
  and (_32346_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_32347_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_32348_, _32347_, _32346_);
  and (_32349_, _32348_, _32345_);
  and (_32350_, _32349_, _32342_);
  nor (_32351_, _32350_, _31948_);
  nor (_32352_, _32351_, _32339_);
  not (_32353_, _32352_);
  and (_32354_, _32353_, _31943_);
  nor (_32355_, _32354_, _32168_);
  not (_32356_, _32355_);
  nor (_32357_, _32356_, _32338_);
  not (_32358_, _32357_);
  nor (_32359_, _32358_, _32336_);
  and (_32360_, _32359_, _32311_);
  nor (_32361_, _32360_, _32312_);
  nor (_32362_, _32361_, _32310_);
  and (_32363_, _32361_, _32310_);
  nor (_32364_, _32363_, _32362_);
  and (_32365_, _32364_, _32309_);
  and (_32366_, _32365_, _32307_);
  and (_32367_, _32366_, _32198_);
  not (_32368_, _32194_);
  and (_32369_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not (_32370_, _32089_);
  and (_32371_, _32370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_32372_, _32371_, _32369_);
  and (_32373_, _32372_, _32303_);
  not (_32374_, _32303_);
  not (_32375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_32376_, _32089_, _32375_);
  and (_32377_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_32378_, _32377_, _32376_);
  and (_32379_, _32378_, _32374_);
  or (_32380_, _32379_, _32373_);
  or (_32381_, _32380_, _32368_);
  not (_32382_, _32361_);
  and (_32383_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_32384_, _32370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_32385_, _32384_, _32383_);
  and (_32386_, _32385_, _32303_);
  not (_32387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_32388_, _32089_, _32387_);
  and (_32389_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or (_32390_, _32389_, _32388_);
  and (_32391_, _32390_, _32374_);
  or (_32392_, _32391_, _32386_);
  or (_32393_, _32392_, _32194_);
  and (_32394_, _32393_, _32382_);
  and (_32395_, _32394_, _32381_);
  or (_32396_, _32370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_32397_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_32398_, _32397_, _32396_);
  and (_32399_, _32398_, _32303_);
  or (_32400_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not (_32401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand (_32402_, _32089_, _32401_);
  and (_32403_, _32402_, _32400_);
  and (_32404_, _32403_, _32374_);
  or (_32405_, _32404_, _32399_);
  or (_32406_, _32405_, _32368_);
  or (_32407_, _32370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_32408_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_32409_, _32408_, _32407_);
  and (_32410_, _32409_, _32303_);
  or (_32411_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not (_32412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand (_32413_, _32089_, _32412_);
  and (_32414_, _32413_, _32411_);
  and (_32415_, _32414_, _32374_);
  or (_32416_, _32415_, _32410_);
  or (_32417_, _32416_, _32194_);
  and (_32418_, _32417_, _32361_);
  and (_32419_, _32418_, _32406_);
  or (_32420_, _32419_, _32395_);
  or (_32421_, _32420_, _32367_);
  not (_32422_, _32367_);
  or (_32423_, _32422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  and (_32424_, _32423_, _35583_);
  and (_35960_[7], _32424_, _32421_);
  nor (_32425_, _31852_, _31848_);
  nor (_32426_, _31900_, _31848_);
  and (_32427_, _32426_, _32425_);
  nor (_32428_, _31896_, _31848_);
  and (_32429_, _31886_, _31847_);
  and (_32430_, _32429_, _32428_);
  and (_32431_, _32430_, _32427_);
  nor (_32432_, _32000_, _31848_);
  and (_32433_, _32432_, _32431_);
  not (_32434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_32435_, _32431_, _32434_);
  or (_35887_, _32435_, _32433_);
  nor (_32436_, _32426_, _32425_);
  nor (_32437_, _32429_, _32428_);
  and (_32438_, _32437_, _31847_);
  and (_32439_, _32438_, _32436_);
  and (_32440_, _31916_, _31847_);
  and (_32441_, _32440_, _32439_);
  not (_32442_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_32443_, _32439_, _32442_);
  or (_35832_, _32443_, _32441_);
  nor (_32444_, _32213_, _31848_);
  and (_32445_, _32444_, _32439_);
  not (_32446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_32447_, _32439_, _32446_);
  or (_35833_, _32447_, _32445_);
  and (_32448_, _32102_, _31847_);
  and (_32449_, _32448_, _32439_);
  not (_32450_, _32439_);
  and (_32451_, _32450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  or (_35834_, _32451_, _32449_);
  and (_32452_, _32048_, _31847_);
  and (_32453_, _32452_, _32439_);
  and (_32454_, _32450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_35835_, _32454_, _32453_);
  nor (_32455_, _32258_, _31848_);
  and (_32456_, _32455_, _32439_);
  and (_32457_, _32450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or (_35836_, _32457_, _32456_);
  nor (_32458_, _32151_, _31848_);
  and (_32459_, _32458_, _32439_);
  and (_32460_, _32450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or (_35837_, _32460_, _32459_);
  nor (_32461_, _32331_, _31848_);
  and (_32462_, _32461_, _32439_);
  and (_32463_, _32450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_35838_, _32463_, _32462_);
  and (_32464_, _32439_, _32432_);
  and (_32465_, _32450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  or (_35839_, _32465_, _32464_);
  and (_32466_, _32425_, _31900_);
  and (_32467_, _32466_, _32437_);
  and (_32468_, _32467_, _32440_);
  not (_32469_, _32467_);
  and (_32470_, _32469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  or (_35888_, _32470_, _32468_);
  and (_32471_, _32467_, _32444_);
  and (_32472_, _32469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  or (_35889_, _32472_, _32471_);
  and (_32473_, _32467_, _32448_);
  and (_32474_, _32469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_35890_, _32474_, _32473_);
  and (_32475_, _32467_, _32452_);
  not (_32476_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_32477_, _32467_, _32476_);
  or (_35891_, _32477_, _32475_);
  and (_32478_, _32467_, _32455_);
  not (_32479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_32480_, _32467_, _32479_);
  or (_35892_, _32480_, _32478_);
  and (_32481_, _32467_, _32458_);
  not (_32482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_32483_, _32467_, _32482_);
  or (_35893_, _32483_, _32481_);
  and (_32484_, _32467_, _32461_);
  not (_32485_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_32486_, _32467_, _32485_);
  or (_35894_, _32486_, _32484_);
  and (_32487_, _32467_, _32432_);
  and (_32488_, _32469_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or (_35895_, _32488_, _32487_);
  and (_32489_, _32426_, _31852_);
  and (_32490_, _32489_, _32437_);
  and (_32491_, _32490_, _32440_);
  not (_32492_, _32490_);
  and (_32493_, _32492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_35896_, _32493_, _32491_);
  and (_32494_, _32490_, _32444_);
  and (_32495_, _32492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_35897_, _32495_, _32494_);
  and (_32496_, _32490_, _32448_);
  not (_32497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_32498_, _32490_, _32497_);
  or (_35898_, _32498_, _32496_);
  and (_32499_, _32490_, _32452_);
  and (_32500_, _32492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_35899_, _32500_, _32499_);
  and (_32501_, _32490_, _32455_);
  not (_32502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_32503_, _32490_, _32502_);
  or (_35900_, _32503_, _32501_);
  and (_32504_, _32490_, _32458_);
  not (_32505_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_32506_, _32490_, _32505_);
  or (_35901_, _32506_, _32504_);
  and (_32507_, _32490_, _32461_);
  and (_32508_, _32492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_35902_, _32508_, _32507_);
  and (_32509_, _32490_, _32432_);
  not (_32510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_32511_, _32490_, _32510_);
  or (_35903_, _32511_, _32509_);
  and (_32512_, _32437_, _32427_);
  and (_32513_, _32512_, _32440_);
  not (_32514_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_32515_, _32512_, _32514_);
  or (_35904_, _32515_, _32513_);
  and (_32516_, _32512_, _32444_);
  not (_32517_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_32518_, _32512_, _32517_);
  or (_35905_, _32518_, _32516_);
  and (_32519_, _32512_, _32448_);
  not (_32520_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_32521_, _32512_, _32520_);
  or (_35906_, _32521_, _32519_);
  and (_32522_, _32512_, _32452_);
  not (_32523_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_32524_, _32512_, _32523_);
  or (_35907_, _32524_, _32522_);
  and (_32525_, _32512_, _32455_);
  not (_32526_, _32512_);
  and (_32527_, _32526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  or (_35908_, _32527_, _32525_);
  and (_32528_, _32512_, _32458_);
  and (_32529_, _32526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  or (_35909_, _32529_, _32528_);
  and (_32530_, _32512_, _32461_);
  not (_32531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor (_32532_, _32512_, _32531_);
  or (_35910_, _32532_, _32530_);
  and (_32533_, _32512_, _32432_);
  nor (_32534_, _32512_, _32375_);
  or (_35911_, _32534_, _32533_);
  and (_32535_, _32428_, _32310_);
  and (_32536_, _32535_, _32436_);
  and (_32537_, _32536_, _32440_);
  not (_32538_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_32539_, _32536_, _32538_);
  or (_35912_, _32539_, _32537_);
  and (_32540_, _32536_, _32444_);
  not (_32541_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_32542_, _32536_, _32541_);
  or (_35913_, _32542_, _32540_);
  and (_32543_, _32536_, _32448_);
  not (_32544_, _32536_);
  and (_32545_, _32544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  or (_35914_, _32545_, _32543_);
  and (_32546_, _32536_, _32452_);
  not (_32547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_32548_, _32536_, _32547_);
  or (_35915_, _32548_, _32546_);
  and (_32549_, _32536_, _32455_);
  and (_32550_, _32544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or (_35916_, _32550_, _32549_);
  and (_32551_, _32536_, _32458_);
  and (_32552_, _32544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or (_35917_, _32552_, _32551_);
  and (_32553_, _32536_, _32461_);
  and (_32554_, _32544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_35918_, _32554_, _32553_);
  and (_32555_, _32536_, _32432_);
  and (_32556_, _32544_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  or (_35919_, _32556_, _32555_);
  and (_32557_, _32535_, _32466_);
  and (_32558_, _32557_, _32440_);
  not (_32559_, _32557_);
  and (_32560_, _32559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  or (_35920_, _32560_, _32558_);
  and (_32561_, _32557_, _32444_);
  and (_32562_, _32559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  or (_35921_, _32562_, _32561_);
  and (_32563_, _32557_, _32448_);
  and (_32564_, _32559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_35922_, _32564_, _32563_);
  and (_32565_, _32557_, _32452_);
  and (_32566_, _32559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_35923_, _32566_, _32565_);
  and (_32567_, _32557_, _32455_);
  not (_32568_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor (_32569_, _32557_, _32568_);
  or (_35924_, _32569_, _32567_);
  and (_32570_, _32557_, _32458_);
  not (_32571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_32572_, _32557_, _32571_);
  or (_35925_, _32572_, _32570_);
  and (_32573_, _32557_, _32461_);
  not (_32574_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_32575_, _32557_, _32574_);
  or (_35926_, _32575_, _32573_);
  and (_32576_, _32557_, _32432_);
  and (_32577_, _32559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or (_35927_, _32577_, _32576_);
  and (_32578_, _32535_, _32489_);
  and (_32579_, _32578_, _32440_);
  not (_32580_, _32578_);
  and (_32581_, _32580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_35928_, _32581_, _32579_);
  and (_32582_, _32578_, _32444_);
  and (_32583_, _32580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_35929_, _32583_, _32582_);
  and (_32584_, _32578_, _32448_);
  not (_32585_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_32586_, _32578_, _32585_);
  or (_35930_, _32586_, _32584_);
  and (_32587_, _32578_, _32452_);
  and (_32588_, _32580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_35931_, _32588_, _32587_);
  and (_32589_, _32578_, _32455_);
  not (_32590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_32591_, _32578_, _32590_);
  or (_35932_, _32591_, _32589_);
  and (_32592_, _32578_, _32458_);
  not (_32593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_32594_, _32578_, _32593_);
  or (_35933_, _32594_, _32592_);
  and (_32595_, _32578_, _32461_);
  and (_32596_, _32580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_35934_, _32596_, _32595_);
  and (_32597_, _32578_, _32432_);
  not (_32598_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_32599_, _32578_, _32598_);
  or (_35935_, _32599_, _32597_);
  and (_32600_, _32535_, _32427_);
  and (_32601_, _32600_, _32440_);
  not (_32602_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_32603_, _32600_, _32602_);
  or (_35936_, _32603_, _32601_);
  and (_32604_, _32600_, _32444_);
  not (_32605_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_32606_, _32600_, _32605_);
  or (_35937_, _32606_, _32604_);
  and (_32607_, _32600_, _32448_);
  not (_32608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_32609_, _32600_, _32608_);
  or (_35938_, _32609_, _32607_);
  and (_32610_, _32600_, _32452_);
  not (_32611_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_32612_, _32600_, _32611_);
  or (_35939_, _32612_, _32610_);
  and (_32613_, _32600_, _32455_);
  not (_32614_, _32600_);
  and (_32615_, _32614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  or (_35940_, _32615_, _32613_);
  and (_32616_, _32600_, _32458_);
  and (_32617_, _32614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  or (_35941_, _32617_, _32616_);
  and (_32618_, _32600_, _32461_);
  not (_32619_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_32620_, _32600_, _32619_);
  or (_35942_, _32620_, _32618_);
  and (_32621_, _32600_, _32432_);
  nor (_32622_, _32600_, _32387_);
  or (_35943_, _32622_, _32621_);
  and (_32623_, _32429_, _31896_);
  and (_32624_, _32623_, _32436_);
  and (_32625_, _32624_, _32440_);
  not (_32626_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_32627_, _32624_, _32626_);
  or (_35944_, _32627_, _32625_);
  and (_32628_, _32624_, _32444_);
  not (_32629_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor (_32630_, _32624_, _32629_);
  or (_35945_, _32630_, _32628_);
  and (_32631_, _32624_, _32448_);
  not (_32632_, _32624_);
  and (_32633_, _32632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_35946_, _32633_, _32631_);
  and (_32634_, _32624_, _32452_);
  and (_32635_, _32632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_35947_, _32635_, _32634_);
  and (_32636_, _32624_, _32455_);
  and (_32637_, _32632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or (_35948_, _32637_, _32636_);
  and (_32638_, _32624_, _32458_);
  and (_32639_, _32632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  or (_35949_, _32639_, _32638_);
  and (_32640_, _32624_, _32461_);
  and (_32641_, _32632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_35950_, _32641_, _32640_);
  and (_32642_, _32624_, _32432_);
  and (_32643_, _32632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  or (_35951_, _32643_, _32642_);
  and (_32644_, _32623_, _32466_);
  and (_32645_, _32644_, _32440_);
  not (_32646_, _32644_);
  and (_32647_, _32646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  or (_35952_, _32647_, _32645_);
  and (_32648_, _32644_, _32444_);
  and (_32649_, _32646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  or (_35953_, _32649_, _32648_);
  and (_32650_, _32644_, _32448_);
  and (_32651_, _32646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  or (_35954_, _32651_, _32650_);
  and (_32652_, _32644_, _32452_);
  and (_32653_, _32646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_35955_, _32653_, _32652_);
  and (_32654_, _32644_, _32455_);
  not (_32655_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_32656_, _32644_, _32655_);
  or (_35956_, _32656_, _32654_);
  and (_32657_, _32644_, _32458_);
  not (_32658_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_32659_, _32644_, _32658_);
  or (_35957_, _32659_, _32657_);
  and (_32660_, _32644_, _32461_);
  and (_32661_, _32646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_35958_, _32661_, _32660_);
  and (_32662_, _32644_, _32432_);
  and (_32663_, _32646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  or (_35959_, _32663_, _32662_);
  and (_32664_, _32623_, _32489_);
  and (_32665_, _32664_, _32440_);
  not (_32666_, _32664_);
  and (_32667_, _32666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  or (_35840_, _32667_, _32665_);
  and (_32668_, _32664_, _32444_);
  and (_32669_, _32666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  or (_35841_, _32669_, _32668_);
  and (_32670_, _32664_, _32448_);
  not (_32671_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_32672_, _32664_, _32671_);
  or (_35842_, _32672_, _32670_);
  and (_32673_, _32664_, _32452_);
  and (_32674_, _32666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_35843_, _32674_, _32673_);
  and (_32675_, _32664_, _32455_);
  not (_32676_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_32677_, _32664_, _32676_);
  or (_35844_, _32677_, _32675_);
  and (_32678_, _32664_, _32458_);
  not (_32679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_32680_, _32664_, _32679_);
  or (_35845_, _32680_, _32678_);
  and (_32681_, _32664_, _32461_);
  not (_32682_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_32683_, _32664_, _32682_);
  or (_35846_, _32683_, _32681_);
  and (_32684_, _32664_, _32432_);
  nor (_32685_, _32664_, _32401_);
  or (_35847_, _32685_, _32684_);
  and (_32686_, _32623_, _32427_);
  and (_32687_, _32686_, _32440_);
  not (_32688_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_32689_, _32686_, _32688_);
  or (_35848_, _32689_, _32687_);
  and (_32690_, _32686_, _32444_);
  not (_32691_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_32692_, _32686_, _32691_);
  or (_35849_, _32692_, _32690_);
  and (_32693_, _32686_, _32448_);
  not (_32694_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_32695_, _32686_, _32694_);
  or (_35850_, _32695_, _32693_);
  and (_32696_, _32686_, _32452_);
  not (_32697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_32698_, _32686_, _32697_);
  or (_35851_, _32698_, _32696_);
  and (_32699_, _32686_, _32455_);
  not (_32700_, _32686_);
  and (_32701_, _32700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  or (_35852_, _32701_, _32699_);
  and (_32702_, _32686_, _32458_);
  and (_32703_, _32700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  or (_35853_, _32703_, _32702_);
  and (_32704_, _32686_, _32461_);
  and (_32705_, _32700_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  or (_35854_, _32705_, _32704_);
  and (_32706_, _32686_, _32432_);
  not (_32707_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_32708_, _32686_, _32707_);
  or (_35855_, _32708_, _32706_);
  and (_32709_, _32436_, _32430_);
  and (_32710_, _32709_, _32440_);
  not (_32711_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_32712_, _32709_, _32711_);
  or (_35856_, _32712_, _32710_);
  and (_32713_, _32709_, _32444_);
  not (_32714_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_32715_, _32709_, _32714_);
  or (_35857_, _32715_, _32713_);
  and (_32716_, _32709_, _32448_);
  not (_32717_, _32709_);
  and (_32718_, _32717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_35858_, _32718_, _32716_);
  and (_32719_, _32709_, _32452_);
  and (_32720_, _32717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  or (_35859_, _32720_, _32719_);
  and (_32721_, _32709_, _32455_);
  and (_32722_, _32717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or (_35860_, _32722_, _32721_);
  and (_32723_, _32709_, _32458_);
  and (_32724_, _32717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  or (_35861_, _32724_, _32723_);
  and (_32725_, _32709_, _32461_);
  and (_32726_, _32717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  or (_35862_, _32726_, _32725_);
  and (_32727_, _32709_, _32432_);
  and (_32728_, _32717_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  or (_35863_, _32728_, _32727_);
  and (_32729_, _32466_, _32430_);
  and (_32730_, _32729_, _32440_);
  not (_32731_, _32729_);
  and (_32732_, _32731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  or (_35864_, _32732_, _32730_);
  and (_32733_, _32729_, _32444_);
  and (_32734_, _32731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  or (_35865_, _32734_, _32733_);
  and (_32735_, _32729_, _32448_);
  and (_32736_, _32731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  or (_35866_, _32736_, _32735_);
  and (_32737_, _32729_, _32452_);
  not (_32738_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_32739_, _32729_, _32738_);
  or (_35867_, _32739_, _32737_);
  and (_32740_, _32729_, _32455_);
  not (_32741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_32742_, _32729_, _32741_);
  or (_35868_, _32742_, _32740_);
  and (_32743_, _32729_, _32458_);
  not (_32744_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_32745_, _32729_, _32744_);
  or (_35869_, _32745_, _32743_);
  and (_32746_, _32729_, _32461_);
  not (_32747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_32748_, _32729_, _32747_);
  or (_35870_, _32748_, _32746_);
  and (_32749_, _32729_, _32432_);
  and (_32750_, _32731_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  or (_35871_, _32750_, _32749_);
  and (_32751_, _32489_, _32430_);
  and (_32752_, _32751_, _32440_);
  not (_32753_, _32751_);
  and (_32754_, _32753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  or (_35872_, _32754_, _32752_);
  and (_32755_, _32751_, _32444_);
  and (_32756_, _32753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  or (_35873_, _32756_, _32755_);
  and (_32757_, _32751_, _32448_);
  not (_32758_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_32759_, _32751_, _32758_);
  or (_35874_, _32759_, _32757_);
  and (_32760_, _32751_, _32452_);
  and (_32761_, _32753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_35875_, _32761_, _32760_);
  and (_32762_, _32751_, _32455_);
  not (_32763_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_32764_, _32751_, _32763_);
  or (_35876_, _32764_, _32762_);
  and (_32765_, _32751_, _32458_);
  not (_32766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_32767_, _32751_, _32766_);
  or (_35877_, _32767_, _32765_);
  and (_32768_, _32751_, _32461_);
  not (_32769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_32770_, _32751_, _32769_);
  or (_35878_, _32770_, _32768_);
  and (_32771_, _32751_, _32432_);
  nor (_32772_, _32751_, _32412_);
  or (_35879_, _32772_, _32771_);
  and (_32773_, _32440_, _32431_);
  not (_32774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_32775_, _32431_, _32774_);
  or (_35880_, _32775_, _32773_);
  and (_32776_, _32444_, _32431_);
  not (_32777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_32778_, _32431_, _32777_);
  or (_35881_, _32778_, _32776_);
  and (_32779_, _32448_, _32431_);
  not (_32780_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_32781_, _32431_, _32780_);
  or (_35882_, _32781_, _32779_);
  and (_32782_, _32452_, _32431_);
  not (_32783_, _32431_);
  and (_32784_, _32783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_35883_, _32784_, _32782_);
  and (_32785_, _32455_, _32431_);
  and (_32786_, _32783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  or (_35884_, _32786_, _32785_);
  and (_32787_, _32458_, _32431_);
  and (_32788_, _32783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  or (_35885_, _32788_, _32787_);
  and (_32789_, _32461_, _32431_);
  and (_32790_, _32783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  or (_35886_, _32790_, _32789_);
  or (_32791_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_32792_, _32089_, _32442_);
  and (_32793_, _32792_, _32303_);
  and (_32794_, _32793_, _32791_);
  nor (_32795_, _32089_, _32514_);
  and (_32796_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or (_32797_, _32796_, _32795_);
  and (_32798_, _32797_, _32374_);
  or (_32799_, _32798_, _32794_);
  or (_32800_, _32799_, _32368_);
  or (_32801_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_32802_, _32089_, _32538_);
  and (_32803_, _32802_, _32303_);
  and (_32804_, _32803_, _32801_);
  nor (_32805_, _32089_, _32602_);
  and (_32806_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or (_32807_, _32806_, _32805_);
  and (_32808_, _32807_, _32374_);
  or (_32809_, _32808_, _32804_);
  or (_32810_, _32809_, _32194_);
  and (_32811_, _32810_, _32382_);
  and (_32812_, _32811_, _32800_);
  nand (_32813_, _32089_, _32626_);
  or (_32814_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_32815_, _32814_, _32813_);
  and (_32816_, _32815_, _32303_);
  and (_32817_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_32818_, _32089_, _32688_);
  or (_32819_, _32818_, _32817_);
  and (_32820_, _32819_, _32374_);
  or (_32821_, _32820_, _32816_);
  or (_32822_, _32821_, _32368_);
  nand (_32823_, _32089_, _32711_);
  or (_32824_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_32825_, _32824_, _32823_);
  and (_32826_, _32825_, _32303_);
  and (_32827_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_32828_, _32089_, _32774_);
  or (_32829_, _32828_, _32827_);
  and (_32830_, _32829_, _32374_);
  or (_32831_, _32830_, _32826_);
  or (_32832_, _32831_, _32194_);
  and (_32833_, _32832_, _32361_);
  and (_32834_, _32833_, _32822_);
  or (_32835_, _32834_, _32812_);
  or (_32836_, _32835_, _32367_);
  or (_32837_, _32422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and (_32838_, _32837_, _35583_);
  and (_35960_[0], _32838_, _32836_);
  or (_32839_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_32840_, _32089_, _32446_);
  and (_32841_, _32840_, _32303_);
  and (_32842_, _32841_, _32839_);
  nor (_32843_, _32089_, _32517_);
  and (_32844_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or (_32845_, _32844_, _32843_);
  and (_32846_, _32845_, _32374_);
  or (_32847_, _32846_, _32842_);
  or (_32848_, _32847_, _32368_);
  or (_32849_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_32850_, _32089_, _32541_);
  and (_32851_, _32850_, _32303_);
  and (_32852_, _32851_, _32849_);
  nor (_32853_, _32089_, _32605_);
  and (_32854_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or (_32855_, _32854_, _32853_);
  and (_32856_, _32855_, _32374_);
  or (_32857_, _32856_, _32852_);
  or (_32858_, _32857_, _32194_);
  and (_32859_, _32858_, _32382_);
  and (_32860_, _32859_, _32848_);
  nand (_32861_, _32089_, _32629_);
  or (_32862_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_32863_, _32862_, _32861_);
  and (_32864_, _32863_, _32303_);
  and (_32865_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_32866_, _32089_, _32691_);
  or (_32867_, _32866_, _32865_);
  and (_32868_, _32867_, _32374_);
  or (_32869_, _32868_, _32864_);
  or (_32870_, _32869_, _32368_);
  nand (_32871_, _32089_, _32714_);
  or (_32872_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_32873_, _32872_, _32871_);
  and (_32874_, _32873_, _32303_);
  and (_32875_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_32876_, _32089_, _32777_);
  or (_32877_, _32876_, _32875_);
  and (_32878_, _32877_, _32374_);
  or (_32879_, _32878_, _32874_);
  or (_32880_, _32879_, _32194_);
  and (_32881_, _32880_, _32361_);
  and (_32882_, _32881_, _32870_);
  or (_32883_, _32882_, _32860_);
  or (_32884_, _32883_, _32367_);
  or (_32885_, _32422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  and (_32886_, _32885_, _35583_);
  and (_35960_[1], _32886_, _32884_);
  and (_32887_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_32888_, _32370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  or (_32889_, _32888_, _32887_);
  and (_32890_, _32889_, _32303_);
  nor (_32891_, _32089_, _32520_);
  and (_32892_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or (_32893_, _32892_, _32891_);
  and (_32894_, _32893_, _32374_);
  or (_32895_, _32894_, _32890_);
  or (_32896_, _32895_, _32368_);
  and (_32897_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_32898_, _32370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  or (_32899_, _32898_, _32897_);
  and (_32900_, _32899_, _32303_);
  nor (_32901_, _32089_, _32608_);
  and (_32902_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_32903_, _32902_, _32901_);
  and (_32904_, _32903_, _32374_);
  or (_32905_, _32904_, _32900_);
  or (_32906_, _32905_, _32194_);
  and (_32907_, _32906_, _32382_);
  and (_32908_, _32907_, _32896_);
  or (_32909_, _32370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  or (_32910_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_32911_, _32910_, _32909_);
  and (_32912_, _32911_, _32303_);
  or (_32913_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand (_32914_, _32089_, _32671_);
  and (_32915_, _32914_, _32913_);
  and (_32916_, _32915_, _32374_);
  or (_32917_, _32916_, _32912_);
  or (_32918_, _32917_, _32368_);
  or (_32919_, _32370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  or (_32920_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_32921_, _32920_, _32919_);
  and (_32922_, _32921_, _32303_);
  or (_32923_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand (_32924_, _32089_, _32758_);
  and (_32925_, _32924_, _32923_);
  and (_32926_, _32925_, _32374_);
  or (_32927_, _32926_, _32922_);
  or (_32928_, _32927_, _32194_);
  and (_32929_, _32928_, _32361_);
  and (_32930_, _32929_, _32918_);
  or (_32931_, _32930_, _32908_);
  or (_32932_, _32931_, _32367_);
  or (_32933_, _32422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and (_32934_, _32933_, _35583_);
  and (_35960_[2], _32934_, _32932_);
  and (_32935_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_32936_, _32089_, _32476_);
  or (_32937_, _32936_, _32935_);
  and (_32938_, _32937_, _32303_);
  nor (_32939_, _32089_, _32523_);
  and (_32940_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_32941_, _32940_, _32939_);
  and (_32942_, _32941_, _32374_);
  or (_32943_, _32942_, _32938_);
  or (_32944_, _32943_, _32368_);
  or (_32945_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nand (_32946_, _32089_, _32547_);
  and (_32947_, _32946_, _32303_);
  and (_32948_, _32947_, _32945_);
  nor (_32949_, _32089_, _32611_);
  and (_32950_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_32951_, _32950_, _32949_);
  and (_32952_, _32951_, _32374_);
  or (_32953_, _32952_, _32948_);
  or (_32954_, _32953_, _32194_);
  and (_32955_, _32954_, _32382_);
  and (_32956_, _32955_, _32944_);
  or (_32957_, _32370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  or (_32958_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_32959_, _32958_, _32957_);
  and (_32960_, _32959_, _32303_);
  and (_32961_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_32962_, _32089_, _32697_);
  or (_32963_, _32962_, _32961_);
  and (_32964_, _32963_, _32374_);
  or (_32965_, _32964_, _32960_);
  or (_32966_, _32965_, _32368_);
  and (_32967_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_32968_, _32089_, _32738_);
  or (_32969_, _32968_, _32967_);
  and (_32970_, _32969_, _32303_);
  or (_32971_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  or (_32972_, _32370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_32973_, _32972_, _32971_);
  and (_32974_, _32973_, _32374_);
  or (_32975_, _32974_, _32970_);
  or (_32976_, _32975_, _32194_);
  and (_32977_, _32976_, _32361_);
  and (_32978_, _32977_, _32966_);
  or (_32979_, _32978_, _32956_);
  or (_32980_, _32979_, _32367_);
  or (_32981_, _32422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  and (_32982_, _32981_, _35583_);
  and (_35960_[3], _32982_, _32980_);
  and (_32983_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_32984_, _32089_, _32479_);
  or (_32985_, _32984_, _32983_);
  and (_32986_, _32985_, _32303_);
  or (_32987_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_32988_, _32089_, _32502_);
  and (_32989_, _32988_, _32987_);
  and (_32990_, _32989_, _32374_);
  or (_32991_, _32990_, _32986_);
  or (_32992_, _32991_, _32368_);
  and (_32993_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_32994_, _32089_, _32568_);
  or (_32995_, _32994_, _32993_);
  and (_32996_, _32995_, _32303_);
  or (_32997_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_32998_, _32089_, _32590_);
  and (_32999_, _32998_, _32997_);
  and (_33000_, _32999_, _32374_);
  or (_33001_, _33000_, _32996_);
  or (_33002_, _33001_, _32194_);
  and (_33003_, _33002_, _32382_);
  and (_33004_, _33003_, _32992_);
  and (_33005_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_33006_, _32089_, _32655_);
  or (_33007_, _33006_, _33005_);
  and (_33008_, _33007_, _32303_);
  or (_33009_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_33010_, _32089_, _32676_);
  and (_33011_, _33010_, _33009_);
  and (_33012_, _33011_, _32374_);
  or (_33013_, _33012_, _33008_);
  or (_33014_, _33013_, _32368_);
  and (_33015_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_33016_, _32089_, _32741_);
  or (_33017_, _33016_, _33015_);
  and (_33018_, _33017_, _32303_);
  or (_33019_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_33020_, _32089_, _32763_);
  and (_33021_, _33020_, _33019_);
  and (_33022_, _33021_, _32374_);
  or (_33023_, _33022_, _33018_);
  or (_33024_, _33023_, _32194_);
  and (_33025_, _33024_, _32361_);
  and (_33026_, _33025_, _33014_);
  or (_33027_, _33026_, _33004_);
  or (_33028_, _33027_, _32367_);
  or (_33029_, _32422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  and (_33030_, _33029_, _35583_);
  and (_35960_[4], _33030_, _33028_);
  and (_33031_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_33032_, _32089_, _32482_);
  or (_33033_, _33032_, _33031_);
  and (_33034_, _33033_, _32303_);
  or (_33035_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_33036_, _32089_, _32505_);
  and (_33037_, _33036_, _33035_);
  and (_33038_, _33037_, _32374_);
  or (_33039_, _33038_, _33034_);
  or (_33040_, _33039_, _32368_);
  and (_33041_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_33042_, _32089_, _32571_);
  or (_33043_, _33042_, _33041_);
  and (_33044_, _33043_, _32303_);
  or (_33045_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_33046_, _32089_, _32593_);
  and (_33047_, _33046_, _33045_);
  and (_33048_, _33047_, _32374_);
  or (_33049_, _33048_, _33044_);
  or (_33050_, _33049_, _32194_);
  and (_33051_, _33050_, _32382_);
  and (_33052_, _33051_, _33040_);
  and (_33053_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_33054_, _32089_, _32658_);
  or (_33055_, _33054_, _33053_);
  and (_33056_, _33055_, _32303_);
  or (_33057_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_33058_, _32089_, _32679_);
  and (_33059_, _33058_, _33057_);
  and (_33060_, _33059_, _32374_);
  or (_33061_, _33060_, _33056_);
  or (_33062_, _33061_, _32368_);
  and (_33063_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_33064_, _32089_, _32744_);
  or (_33065_, _33064_, _33063_);
  and (_33066_, _33065_, _32303_);
  or (_33067_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_33068_, _32089_, _32766_);
  and (_33069_, _33068_, _33067_);
  and (_33070_, _33069_, _32374_);
  or (_33071_, _33070_, _33066_);
  or (_33072_, _33071_, _32194_);
  and (_33073_, _33072_, _32361_);
  and (_33074_, _33073_, _33062_);
  or (_33075_, _33074_, _33052_);
  or (_33076_, _33075_, _32367_);
  or (_33077_, _32422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and (_33078_, _33077_, _35583_);
  and (_35960_[5], _33078_, _33076_);
  and (_33079_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_33080_, _32089_, _32485_);
  or (_33081_, _33080_, _33079_);
  and (_33082_, _33081_, _32303_);
  nor (_33083_, _32089_, _32531_);
  and (_33084_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_33085_, _33084_, _33083_);
  and (_33086_, _33085_, _32374_);
  or (_33087_, _33086_, _33082_);
  or (_33088_, _33087_, _32368_);
  and (_33089_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_33090_, _32089_, _32574_);
  or (_33091_, _33090_, _33089_);
  and (_33092_, _33091_, _32303_);
  nor (_33093_, _32089_, _32619_);
  and (_33094_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_33095_, _33094_, _33093_);
  and (_33096_, _33095_, _32374_);
  or (_33097_, _33096_, _33092_);
  or (_33098_, _33097_, _32194_);
  and (_33099_, _33098_, _32382_);
  and (_33100_, _33099_, _33088_);
  or (_33101_, _32370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  or (_33102_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_33103_, _33102_, _33101_);
  and (_33104_, _33103_, _32303_);
  or (_33105_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_33106_, _32089_, _32682_);
  and (_33107_, _33106_, _33105_);
  and (_33108_, _33107_, _32374_);
  or (_33109_, _33108_, _33104_);
  or (_33110_, _33109_, _32368_);
  and (_33111_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_33112_, _32089_, _32747_);
  or (_33113_, _33112_, _33111_);
  and (_33114_, _33113_, _32303_);
  or (_33115_, _32089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_33116_, _32089_, _32769_);
  and (_33117_, _33116_, _33115_);
  and (_33118_, _33117_, _32374_);
  or (_33119_, _33118_, _33114_);
  or (_33120_, _33119_, _32194_);
  and (_33121_, _33120_, _32361_);
  and (_33122_, _33121_, _33110_);
  or (_33123_, _33122_, _33100_);
  or (_33124_, _33123_, _32367_);
  or (_33125_, _32422_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and (_33126_, _33125_, _35583_);
  and (_35960_[6], _33126_, _33124_);
  or (_33127_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not (_33128_, \oc8051_gm_cxrom_1.cell0.valid );
  or (_33129_, _33128_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand (_33130_, _33129_, _33127_);
  nand (_33131_, _33130_, _35583_);
  or (_33132_, \oc8051_gm_cxrom_1.cell0.data [7], _35583_);
  and (_35582_[7], _33132_, _33131_);
  or (_33133_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33134_, \oc8051_gm_cxrom_1.cell0.data [0], _33128_);
  nand (_33135_, _33134_, _33133_);
  nand (_33136_, _33135_, _35583_);
  or (_33137_, \oc8051_gm_cxrom_1.cell0.data [0], _35583_);
  and (_35582_[0], _33137_, _33136_);
  or (_33138_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33139_, \oc8051_gm_cxrom_1.cell0.data [1], _33128_);
  nand (_33140_, _33139_, _33138_);
  nand (_33141_, _33140_, _35583_);
  or (_33142_, \oc8051_gm_cxrom_1.cell0.data [1], _35583_);
  and (_35582_[1], _33142_, _33141_);
  or (_33143_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33144_, \oc8051_gm_cxrom_1.cell0.data [2], _33128_);
  nand (_33145_, _33144_, _33143_);
  nand (_33146_, _33145_, _35583_);
  or (_33147_, \oc8051_gm_cxrom_1.cell0.data [2], _35583_);
  and (_35582_[2], _33147_, _33146_);
  or (_33148_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33149_, \oc8051_gm_cxrom_1.cell0.data [3], _33128_);
  nand (_33150_, _33149_, _33148_);
  nand (_33151_, _33150_, _35583_);
  or (_33152_, \oc8051_gm_cxrom_1.cell0.data [3], _35583_);
  and (_35582_[3], _33152_, _33151_);
  or (_33153_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33154_, \oc8051_gm_cxrom_1.cell0.data [4], _33128_);
  nand (_33155_, _33154_, _33153_);
  nand (_33156_, _33155_, _35583_);
  or (_33157_, \oc8051_gm_cxrom_1.cell0.data [4], _35583_);
  and (_35582_[4], _33157_, _33156_);
  or (_33158_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33159_, \oc8051_gm_cxrom_1.cell0.data [5], _33128_);
  nand (_33160_, _33159_, _33158_);
  nand (_33161_, _33160_, _35583_);
  or (_33162_, \oc8051_gm_cxrom_1.cell0.data [5], _35583_);
  and (_35582_[5], _33162_, _33161_);
  or (_33163_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or (_33164_, \oc8051_gm_cxrom_1.cell0.data [6], _33128_);
  nand (_33165_, _33164_, _33163_);
  nand (_33166_, _33165_, _35583_);
  or (_33167_, \oc8051_gm_cxrom_1.cell0.data [6], _35583_);
  and (_35582_[6], _33167_, _33166_);
  or (_33168_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not (_33169_, \oc8051_gm_cxrom_1.cell1.valid );
  or (_33170_, _33169_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand (_33171_, _33170_, _33168_);
  nand (_33172_, _33171_, _35583_);
  or (_33173_, \oc8051_gm_cxrom_1.cell1.data [7], _35583_);
  and (_35584_[7], _33173_, _33172_);
  or (_33174_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33175_, \oc8051_gm_cxrom_1.cell1.data [0], _33169_);
  nand (_33176_, _33175_, _33174_);
  nand (_33177_, _33176_, _35583_);
  or (_33178_, \oc8051_gm_cxrom_1.cell1.data [0], _35583_);
  and (_35584_[0], _33178_, _33177_);
  or (_33179_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33180_, \oc8051_gm_cxrom_1.cell1.data [1], _33169_);
  nand (_33181_, _33180_, _33179_);
  nand (_33182_, _33181_, _35583_);
  or (_33183_, \oc8051_gm_cxrom_1.cell1.data [1], _35583_);
  and (_35584_[1], _33183_, _33182_);
  or (_33184_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33185_, \oc8051_gm_cxrom_1.cell1.data [2], _33169_);
  nand (_33186_, _33185_, _33184_);
  nand (_33187_, _33186_, _35583_);
  or (_33188_, \oc8051_gm_cxrom_1.cell1.data [2], _35583_);
  and (_35584_[2], _33188_, _33187_);
  or (_33189_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33190_, \oc8051_gm_cxrom_1.cell1.data [3], _33169_);
  nand (_33191_, _33190_, _33189_);
  nand (_33192_, _33191_, _35583_);
  or (_33193_, \oc8051_gm_cxrom_1.cell1.data [3], _35583_);
  and (_35584_[3], _33193_, _33192_);
  or (_33194_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33195_, \oc8051_gm_cxrom_1.cell1.data [4], _33169_);
  nand (_33196_, _33195_, _33194_);
  nand (_33197_, _33196_, _35583_);
  or (_33198_, \oc8051_gm_cxrom_1.cell1.data [4], _35583_);
  and (_35584_[4], _33198_, _33197_);
  or (_33199_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33200_, \oc8051_gm_cxrom_1.cell1.data [5], _33169_);
  nand (_33201_, _33200_, _33199_);
  nand (_33202_, _33201_, _35583_);
  or (_33203_, \oc8051_gm_cxrom_1.cell1.data [5], _35583_);
  and (_35584_[5], _33203_, _33202_);
  or (_33204_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or (_33205_, \oc8051_gm_cxrom_1.cell1.data [6], _33169_);
  nand (_33206_, _33205_, _33204_);
  nand (_33207_, _33206_, _35583_);
  or (_33208_, \oc8051_gm_cxrom_1.cell1.data [6], _35583_);
  and (_35584_[6], _33208_, _33207_);
  or (_33209_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not (_33210_, \oc8051_gm_cxrom_1.cell2.valid );
  or (_33211_, _33210_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand (_33212_, _33211_, _33209_);
  nand (_33213_, _33212_, _35583_);
  or (_33214_, \oc8051_gm_cxrom_1.cell2.data [7], _35583_);
  and (_35598_[7], _33214_, _33213_);
  or (_33215_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33216_, \oc8051_gm_cxrom_1.cell2.data [0], _33210_);
  nand (_33217_, _33216_, _33215_);
  nand (_33218_, _33217_, _35583_);
  or (_33219_, \oc8051_gm_cxrom_1.cell2.data [0], _35583_);
  and (_35598_[0], _33219_, _33218_);
  or (_33220_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33221_, \oc8051_gm_cxrom_1.cell2.data [1], _33210_);
  nand (_33222_, _33221_, _33220_);
  nand (_33223_, _33222_, _35583_);
  or (_33224_, \oc8051_gm_cxrom_1.cell2.data [1], _35583_);
  and (_35598_[1], _33224_, _33223_);
  or (_33225_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33226_, \oc8051_gm_cxrom_1.cell2.data [2], _33210_);
  nand (_33227_, _33226_, _33225_);
  nand (_33228_, _33227_, _35583_);
  or (_33229_, \oc8051_gm_cxrom_1.cell2.data [2], _35583_);
  and (_35598_[2], _33229_, _33228_);
  or (_33230_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33231_, \oc8051_gm_cxrom_1.cell2.data [3], _33210_);
  nand (_33232_, _33231_, _33230_);
  nand (_33233_, _33232_, _35583_);
  or (_33234_, \oc8051_gm_cxrom_1.cell2.data [3], _35583_);
  and (_35598_[3], _33234_, _33233_);
  or (_33235_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33236_, \oc8051_gm_cxrom_1.cell2.data [4], _33210_);
  nand (_33237_, _33236_, _33235_);
  nand (_33238_, _33237_, _35583_);
  or (_33239_, \oc8051_gm_cxrom_1.cell2.data [4], _35583_);
  and (_35598_[4], _33239_, _33238_);
  or (_33240_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33241_, \oc8051_gm_cxrom_1.cell2.data [5], _33210_);
  nand (_33242_, _33241_, _33240_);
  nand (_33243_, _33242_, _35583_);
  or (_33244_, \oc8051_gm_cxrom_1.cell2.data [5], _35583_);
  and (_35598_[5], _33244_, _33243_);
  or (_33245_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or (_33246_, \oc8051_gm_cxrom_1.cell2.data [6], _33210_);
  nand (_33247_, _33246_, _33245_);
  nand (_33248_, _33247_, _35583_);
  or (_33249_, \oc8051_gm_cxrom_1.cell2.data [6], _35583_);
  and (_35598_[6], _33249_, _33248_);
  or (_33250_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not (_33251_, \oc8051_gm_cxrom_1.cell3.valid );
  or (_33252_, _33251_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand (_33253_, _33252_, _33250_);
  nand (_33254_, _33253_, _35583_);
  or (_33255_, \oc8051_gm_cxrom_1.cell3.data [7], _35583_);
  and (_35600_[7], _33255_, _33254_);
  or (_33256_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33257_, \oc8051_gm_cxrom_1.cell3.data [0], _33251_);
  nand (_33258_, _33257_, _33256_);
  nand (_33259_, _33258_, _35583_);
  or (_33260_, \oc8051_gm_cxrom_1.cell3.data [0], _35583_);
  and (_35600_[0], _33260_, _33259_);
  or (_33261_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33262_, \oc8051_gm_cxrom_1.cell3.data [1], _33251_);
  nand (_33263_, _33262_, _33261_);
  nand (_33264_, _33263_, _35583_);
  or (_33265_, \oc8051_gm_cxrom_1.cell3.data [1], _35583_);
  and (_35600_[1], _33265_, _33264_);
  or (_33266_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33267_, \oc8051_gm_cxrom_1.cell3.data [2], _33251_);
  nand (_33268_, _33267_, _33266_);
  nand (_33269_, _33268_, _35583_);
  or (_33270_, \oc8051_gm_cxrom_1.cell3.data [2], _35583_);
  and (_35600_[2], _33270_, _33269_);
  or (_33271_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33272_, \oc8051_gm_cxrom_1.cell3.data [3], _33251_);
  nand (_33273_, _33272_, _33271_);
  nand (_33274_, _33273_, _35583_);
  or (_33275_, \oc8051_gm_cxrom_1.cell3.data [3], _35583_);
  and (_35600_[3], _33275_, _33274_);
  or (_33276_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33277_, \oc8051_gm_cxrom_1.cell3.data [4], _33251_);
  nand (_33278_, _33277_, _33276_);
  nand (_33279_, _33278_, _35583_);
  or (_33280_, \oc8051_gm_cxrom_1.cell3.data [4], _35583_);
  and (_35600_[4], _33280_, _33279_);
  or (_33281_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33282_, \oc8051_gm_cxrom_1.cell3.data [5], _33251_);
  nand (_33283_, _33282_, _33281_);
  nand (_33284_, _33283_, _35583_);
  or (_33285_, \oc8051_gm_cxrom_1.cell3.data [5], _35583_);
  and (_35600_[5], _33285_, _33284_);
  or (_33286_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or (_33287_, \oc8051_gm_cxrom_1.cell3.data [6], _33251_);
  nand (_33288_, _33287_, _33286_);
  nand (_33289_, _33288_, _35583_);
  or (_33290_, \oc8051_gm_cxrom_1.cell3.data [6], _35583_);
  and (_35600_[6], _33290_, _33289_);
  or (_33291_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not (_33292_, \oc8051_gm_cxrom_1.cell4.valid );
  or (_33293_, _33292_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand (_33294_, _33293_, _33291_);
  nand (_33295_, _33294_, _35583_);
  or (_33296_, \oc8051_gm_cxrom_1.cell4.data [7], _35583_);
  and (_35602_[7], _33296_, _33295_);
  or (_33297_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33298_, \oc8051_gm_cxrom_1.cell4.data [0], _33292_);
  nand (_33299_, _33298_, _33297_);
  nand (_33300_, _33299_, _35583_);
  or (_33301_, \oc8051_gm_cxrom_1.cell4.data [0], _35583_);
  and (_35602_[0], _33301_, _33300_);
  or (_33302_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33303_, \oc8051_gm_cxrom_1.cell4.data [1], _33292_);
  nand (_33304_, _33303_, _33302_);
  nand (_33305_, _33304_, _35583_);
  or (_33306_, \oc8051_gm_cxrom_1.cell4.data [1], _35583_);
  and (_35602_[1], _33306_, _33305_);
  or (_33307_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33308_, \oc8051_gm_cxrom_1.cell4.data [2], _33292_);
  nand (_33309_, _33308_, _33307_);
  nand (_33310_, _33309_, _35583_);
  or (_33311_, \oc8051_gm_cxrom_1.cell4.data [2], _35583_);
  and (_35602_[2], _33311_, _33310_);
  or (_33312_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33313_, \oc8051_gm_cxrom_1.cell4.data [3], _33292_);
  nand (_33314_, _33313_, _33312_);
  nand (_33315_, _33314_, _35583_);
  or (_33316_, \oc8051_gm_cxrom_1.cell4.data [3], _35583_);
  and (_35602_[3], _33316_, _33315_);
  or (_33317_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33318_, \oc8051_gm_cxrom_1.cell4.data [4], _33292_);
  nand (_33319_, _33318_, _33317_);
  nand (_33320_, _33319_, _35583_);
  or (_33321_, \oc8051_gm_cxrom_1.cell4.data [4], _35583_);
  and (_35602_[4], _33321_, _33320_);
  or (_33322_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33323_, \oc8051_gm_cxrom_1.cell4.data [5], _33292_);
  nand (_33324_, _33323_, _33322_);
  nand (_33325_, _33324_, _35583_);
  or (_33326_, \oc8051_gm_cxrom_1.cell4.data [5], _35583_);
  and (_35602_[5], _33326_, _33325_);
  or (_33327_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or (_33328_, \oc8051_gm_cxrom_1.cell4.data [6], _33292_);
  nand (_33329_, _33328_, _33327_);
  nand (_33330_, _33329_, _35583_);
  or (_33331_, \oc8051_gm_cxrom_1.cell4.data [6], _35583_);
  and (_35602_[6], _33331_, _33330_);
  or (_33332_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not (_33333_, \oc8051_gm_cxrom_1.cell5.valid );
  or (_33334_, _33333_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand (_33335_, _33334_, _33332_);
  nand (_33336_, _33335_, _35583_);
  or (_33337_, \oc8051_gm_cxrom_1.cell5.data [7], _35583_);
  and (_35604_[7], _33337_, _33336_);
  or (_33338_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33339_, \oc8051_gm_cxrom_1.cell5.data [0], _33333_);
  nand (_33340_, _33339_, _33338_);
  nand (_33341_, _33340_, _35583_);
  or (_33342_, \oc8051_gm_cxrom_1.cell5.data [0], _35583_);
  and (_35604_[0], _33342_, _33341_);
  or (_33343_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33344_, \oc8051_gm_cxrom_1.cell5.data [1], _33333_);
  nand (_33345_, _33344_, _33343_);
  nand (_33346_, _33345_, _35583_);
  or (_33347_, \oc8051_gm_cxrom_1.cell5.data [1], _35583_);
  and (_35604_[1], _33347_, _33346_);
  or (_33348_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33349_, \oc8051_gm_cxrom_1.cell5.data [2], _33333_);
  nand (_33350_, _33349_, _33348_);
  nand (_33351_, _33350_, _35583_);
  or (_33352_, \oc8051_gm_cxrom_1.cell5.data [2], _35583_);
  and (_35604_[2], _33352_, _33351_);
  or (_33353_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33354_, \oc8051_gm_cxrom_1.cell5.data [3], _33333_);
  nand (_33355_, _33354_, _33353_);
  nand (_33356_, _33355_, _35583_);
  or (_33357_, \oc8051_gm_cxrom_1.cell5.data [3], _35583_);
  and (_35604_[3], _33357_, _33356_);
  or (_33358_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33359_, \oc8051_gm_cxrom_1.cell5.data [4], _33333_);
  nand (_33360_, _33359_, _33358_);
  nand (_33361_, _33360_, _35583_);
  or (_33362_, \oc8051_gm_cxrom_1.cell5.data [4], _35583_);
  and (_35604_[4], _33362_, _33361_);
  or (_33363_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33364_, \oc8051_gm_cxrom_1.cell5.data [5], _33333_);
  nand (_33365_, _33364_, _33363_);
  nand (_33366_, _33365_, _35583_);
  or (_33367_, \oc8051_gm_cxrom_1.cell5.data [5], _35583_);
  and (_35604_[5], _33367_, _33366_);
  or (_33368_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or (_33369_, \oc8051_gm_cxrom_1.cell5.data [6], _33333_);
  nand (_33370_, _33369_, _33368_);
  nand (_33371_, _33370_, _35583_);
  or (_33372_, \oc8051_gm_cxrom_1.cell5.data [6], _35583_);
  and (_35604_[6], _33372_, _33371_);
  or (_33373_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not (_33374_, \oc8051_gm_cxrom_1.cell6.valid );
  or (_33375_, _33374_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand (_33376_, _33375_, _33373_);
  nand (_33377_, _33376_, _35583_);
  or (_33378_, \oc8051_gm_cxrom_1.cell6.data [7], _35583_);
  and (_35606_[7], _33378_, _33377_);
  or (_33379_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33380_, \oc8051_gm_cxrom_1.cell6.data [0], _33374_);
  nand (_33381_, _33380_, _33379_);
  nand (_33382_, _33381_, _35583_);
  or (_33383_, \oc8051_gm_cxrom_1.cell6.data [0], _35583_);
  and (_35606_[0], _33383_, _33382_);
  or (_33384_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33385_, \oc8051_gm_cxrom_1.cell6.data [1], _33374_);
  nand (_33386_, _33385_, _33384_);
  nand (_33387_, _33386_, _35583_);
  or (_33388_, \oc8051_gm_cxrom_1.cell6.data [1], _35583_);
  and (_35606_[1], _33388_, _33387_);
  or (_33389_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33390_, \oc8051_gm_cxrom_1.cell6.data [2], _33374_);
  nand (_33391_, _33390_, _33389_);
  nand (_33392_, _33391_, _35583_);
  or (_33393_, \oc8051_gm_cxrom_1.cell6.data [2], _35583_);
  and (_35606_[2], _33393_, _33392_);
  or (_33394_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33395_, \oc8051_gm_cxrom_1.cell6.data [3], _33374_);
  nand (_33396_, _33395_, _33394_);
  nand (_33397_, _33396_, _35583_);
  or (_33398_, \oc8051_gm_cxrom_1.cell6.data [3], _35583_);
  and (_35606_[3], _33398_, _33397_);
  or (_33399_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33400_, \oc8051_gm_cxrom_1.cell6.data [4], _33374_);
  nand (_33401_, _33400_, _33399_);
  nand (_33402_, _33401_, _35583_);
  or (_33403_, \oc8051_gm_cxrom_1.cell6.data [4], _35583_);
  and (_35606_[4], _33403_, _33402_);
  or (_33404_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33405_, \oc8051_gm_cxrom_1.cell6.data [5], _33374_);
  nand (_33406_, _33405_, _33404_);
  nand (_33407_, _33406_, _35583_);
  or (_33408_, \oc8051_gm_cxrom_1.cell6.data [5], _35583_);
  and (_35606_[5], _33408_, _33407_);
  or (_33409_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or (_33410_, \oc8051_gm_cxrom_1.cell6.data [6], _33374_);
  nand (_33411_, _33410_, _33409_);
  nand (_33412_, _33411_, _35583_);
  or (_33413_, \oc8051_gm_cxrom_1.cell6.data [6], _35583_);
  and (_35606_[6], _33413_, _33412_);
  or (_33414_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not (_33415_, \oc8051_gm_cxrom_1.cell7.valid );
  or (_33416_, _33415_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand (_33417_, _33416_, _33414_);
  nand (_33418_, _33417_, _35583_);
  or (_33419_, \oc8051_gm_cxrom_1.cell7.data [7], _35583_);
  and (_35608_[7], _33419_, _33418_);
  or (_33420_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33421_, \oc8051_gm_cxrom_1.cell7.data [0], _33415_);
  nand (_33422_, _33421_, _33420_);
  nand (_33423_, _33422_, _35583_);
  or (_33424_, \oc8051_gm_cxrom_1.cell7.data [0], _35583_);
  and (_35608_[0], _33424_, _33423_);
  or (_33425_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33426_, \oc8051_gm_cxrom_1.cell7.data [1], _33415_);
  nand (_33427_, _33426_, _33425_);
  nand (_33428_, _33427_, _35583_);
  or (_33429_, \oc8051_gm_cxrom_1.cell7.data [1], _35583_);
  and (_35608_[1], _33429_, _33428_);
  or (_33430_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33431_, \oc8051_gm_cxrom_1.cell7.data [2], _33415_);
  nand (_33432_, _33431_, _33430_);
  nand (_33433_, _33432_, _35583_);
  or (_33434_, \oc8051_gm_cxrom_1.cell7.data [2], _35583_);
  and (_35608_[2], _33434_, _33433_);
  or (_33435_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33436_, \oc8051_gm_cxrom_1.cell7.data [3], _33415_);
  nand (_33437_, _33436_, _33435_);
  nand (_33438_, _33437_, _35583_);
  or (_33439_, \oc8051_gm_cxrom_1.cell7.data [3], _35583_);
  and (_35608_[3], _33439_, _33438_);
  or (_33440_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33441_, \oc8051_gm_cxrom_1.cell7.data [4], _33415_);
  nand (_33442_, _33441_, _33440_);
  nand (_33443_, _33442_, _35583_);
  or (_33444_, \oc8051_gm_cxrom_1.cell7.data [4], _35583_);
  and (_35608_[4], _33444_, _33443_);
  or (_33445_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33446_, \oc8051_gm_cxrom_1.cell7.data [5], _33415_);
  nand (_33447_, _33446_, _33445_);
  nand (_33448_, _33447_, _35583_);
  or (_33449_, \oc8051_gm_cxrom_1.cell7.data [5], _35583_);
  and (_35608_[5], _33449_, _33448_);
  or (_33450_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or (_33451_, \oc8051_gm_cxrom_1.cell7.data [6], _33415_);
  nand (_33452_, _33451_, _33450_);
  nand (_33453_, _33452_, _35583_);
  or (_33454_, \oc8051_gm_cxrom_1.cell7.data [6], _35583_);
  and (_35608_[6], _33454_, _33453_);
  or (_33455_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not (_33456_, \oc8051_gm_cxrom_1.cell8.valid );
  or (_33457_, _33456_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand (_33458_, _33457_, _33455_);
  nand (_33459_, _33458_, _35583_);
  or (_33460_, \oc8051_gm_cxrom_1.cell8.data [7], _35583_);
  and (_35610_[7], _33460_, _33459_);
  or (_33461_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33462_, \oc8051_gm_cxrom_1.cell8.data [0], _33456_);
  nand (_33463_, _33462_, _33461_);
  nand (_33464_, _33463_, _35583_);
  or (_33465_, \oc8051_gm_cxrom_1.cell8.data [0], _35583_);
  and (_35610_[0], _33465_, _33464_);
  or (_33466_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33467_, \oc8051_gm_cxrom_1.cell8.data [1], _33456_);
  nand (_33468_, _33467_, _33466_);
  nand (_33469_, _33468_, _35583_);
  or (_33470_, \oc8051_gm_cxrom_1.cell8.data [1], _35583_);
  and (_35610_[1], _33470_, _33469_);
  or (_33471_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33472_, \oc8051_gm_cxrom_1.cell8.data [2], _33456_);
  nand (_33473_, _33472_, _33471_);
  nand (_33474_, _33473_, _35583_);
  or (_33475_, \oc8051_gm_cxrom_1.cell8.data [2], _35583_);
  and (_35610_[2], _33475_, _33474_);
  or (_33476_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33477_, \oc8051_gm_cxrom_1.cell8.data [3], _33456_);
  nand (_33478_, _33477_, _33476_);
  nand (_33479_, _33478_, _35583_);
  or (_33480_, \oc8051_gm_cxrom_1.cell8.data [3], _35583_);
  and (_35610_[3], _33480_, _33479_);
  or (_33481_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33482_, \oc8051_gm_cxrom_1.cell8.data [4], _33456_);
  nand (_33483_, _33482_, _33481_);
  nand (_33484_, _33483_, _35583_);
  or (_33485_, \oc8051_gm_cxrom_1.cell8.data [4], _35583_);
  and (_35610_[4], _33485_, _33484_);
  or (_33486_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33487_, \oc8051_gm_cxrom_1.cell8.data [5], _33456_);
  nand (_33488_, _33487_, _33486_);
  nand (_33489_, _33488_, _35583_);
  or (_33490_, \oc8051_gm_cxrom_1.cell8.data [5], _35583_);
  and (_35610_[5], _33490_, _33489_);
  or (_33491_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or (_33492_, \oc8051_gm_cxrom_1.cell8.data [6], _33456_);
  nand (_33493_, _33492_, _33491_);
  nand (_33494_, _33493_, _35583_);
  or (_33495_, \oc8051_gm_cxrom_1.cell8.data [6], _35583_);
  and (_35610_[6], _33495_, _33494_);
  or (_33496_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not (_33497_, \oc8051_gm_cxrom_1.cell9.valid );
  or (_33498_, _33497_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand (_33499_, _33498_, _33496_);
  nand (_33500_, _33499_, _35583_);
  or (_33501_, \oc8051_gm_cxrom_1.cell9.data [7], _35583_);
  and (_35612_[7], _33501_, _33500_);
  or (_33502_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33503_, \oc8051_gm_cxrom_1.cell9.data [0], _33497_);
  nand (_33504_, _33503_, _33502_);
  nand (_33505_, _33504_, _35583_);
  or (_33506_, \oc8051_gm_cxrom_1.cell9.data [0], _35583_);
  and (_35612_[0], _33506_, _33505_);
  or (_33507_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33508_, \oc8051_gm_cxrom_1.cell9.data [1], _33497_);
  nand (_33509_, _33508_, _33507_);
  nand (_33510_, _33509_, _35583_);
  or (_33511_, \oc8051_gm_cxrom_1.cell9.data [1], _35583_);
  and (_35612_[1], _33511_, _33510_);
  or (_33512_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33513_, \oc8051_gm_cxrom_1.cell9.data [2], _33497_);
  nand (_33514_, _33513_, _33512_);
  nand (_33515_, _33514_, _35583_);
  or (_33516_, \oc8051_gm_cxrom_1.cell9.data [2], _35583_);
  and (_35612_[2], _33516_, _33515_);
  or (_33517_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33518_, \oc8051_gm_cxrom_1.cell9.data [3], _33497_);
  nand (_33519_, _33518_, _33517_);
  nand (_33520_, _33519_, _35583_);
  or (_33521_, \oc8051_gm_cxrom_1.cell9.data [3], _35583_);
  and (_35612_[3], _33521_, _33520_);
  or (_33522_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33523_, \oc8051_gm_cxrom_1.cell9.data [4], _33497_);
  nand (_33524_, _33523_, _33522_);
  nand (_33525_, _33524_, _35583_);
  or (_33526_, \oc8051_gm_cxrom_1.cell9.data [4], _35583_);
  and (_35612_[4], _33526_, _33525_);
  or (_33527_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33528_, \oc8051_gm_cxrom_1.cell9.data [5], _33497_);
  nand (_33529_, _33528_, _33527_);
  nand (_33530_, _33529_, _35583_);
  or (_33531_, \oc8051_gm_cxrom_1.cell9.data [5], _35583_);
  and (_35612_[5], _33531_, _33530_);
  or (_33532_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or (_33533_, \oc8051_gm_cxrom_1.cell9.data [6], _33497_);
  nand (_33534_, _33533_, _33532_);
  nand (_33535_, _33534_, _35583_);
  or (_33536_, \oc8051_gm_cxrom_1.cell9.data [6], _35583_);
  and (_35612_[6], _33536_, _33535_);
  or (_33537_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not (_33538_, \oc8051_gm_cxrom_1.cell10.valid );
  or (_33539_, _33538_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand (_33540_, _33539_, _33537_);
  nand (_33541_, _33540_, _35583_);
  or (_33542_, \oc8051_gm_cxrom_1.cell10.data [7], _35583_);
  and (_35586_[7], _33542_, _33541_);
  or (_33543_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33544_, \oc8051_gm_cxrom_1.cell10.data [0], _33538_);
  nand (_33545_, _33544_, _33543_);
  nand (_33546_, _33545_, _35583_);
  or (_33547_, \oc8051_gm_cxrom_1.cell10.data [0], _35583_);
  and (_35586_[0], _33547_, _33546_);
  or (_33548_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33549_, \oc8051_gm_cxrom_1.cell10.data [1], _33538_);
  nand (_33550_, _33549_, _33548_);
  nand (_33551_, _33550_, _35583_);
  or (_33552_, \oc8051_gm_cxrom_1.cell10.data [1], _35583_);
  and (_35586_[1], _33552_, _33551_);
  or (_33553_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33554_, \oc8051_gm_cxrom_1.cell10.data [2], _33538_);
  nand (_33555_, _33554_, _33553_);
  nand (_33556_, _33555_, _35583_);
  or (_33557_, \oc8051_gm_cxrom_1.cell10.data [2], _35583_);
  and (_35586_[2], _33557_, _33556_);
  or (_33558_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33559_, \oc8051_gm_cxrom_1.cell10.data [3], _33538_);
  nand (_33560_, _33559_, _33558_);
  nand (_33561_, _33560_, _35583_);
  or (_33562_, \oc8051_gm_cxrom_1.cell10.data [3], _35583_);
  and (_35586_[3], _33562_, _33561_);
  or (_33563_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33564_, \oc8051_gm_cxrom_1.cell10.data [4], _33538_);
  nand (_33565_, _33564_, _33563_);
  nand (_33566_, _33565_, _35583_);
  or (_33567_, \oc8051_gm_cxrom_1.cell10.data [4], _35583_);
  and (_35586_[4], _33567_, _33566_);
  or (_33568_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33569_, \oc8051_gm_cxrom_1.cell10.data [5], _33538_);
  nand (_33570_, _33569_, _33568_);
  nand (_33571_, _33570_, _35583_);
  or (_33572_, \oc8051_gm_cxrom_1.cell10.data [5], _35583_);
  and (_35586_[5], _33572_, _33571_);
  or (_33573_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or (_33574_, \oc8051_gm_cxrom_1.cell10.data [6], _33538_);
  nand (_33575_, _33574_, _33573_);
  nand (_33576_, _33575_, _35583_);
  or (_33577_, \oc8051_gm_cxrom_1.cell10.data [6], _35583_);
  and (_35586_[6], _33577_, _33576_);
  or (_33578_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not (_33579_, \oc8051_gm_cxrom_1.cell11.valid );
  or (_33580_, _33579_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand (_33581_, _33580_, _33578_);
  nand (_33582_, _33581_, _35583_);
  or (_33583_, \oc8051_gm_cxrom_1.cell11.data [7], _35583_);
  and (_35588_[7], _33583_, _33582_);
  or (_33584_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33585_, \oc8051_gm_cxrom_1.cell11.data [0], _33579_);
  nand (_33586_, _33585_, _33584_);
  nand (_33587_, _33586_, _35583_);
  or (_33588_, \oc8051_gm_cxrom_1.cell11.data [0], _35583_);
  and (_35588_[0], _33588_, _33587_);
  or (_33589_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33590_, \oc8051_gm_cxrom_1.cell11.data [1], _33579_);
  nand (_33591_, _33590_, _33589_);
  nand (_33592_, _33591_, _35583_);
  or (_33593_, \oc8051_gm_cxrom_1.cell11.data [1], _35583_);
  and (_35588_[1], _33593_, _33592_);
  or (_33594_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33595_, \oc8051_gm_cxrom_1.cell11.data [2], _33579_);
  nand (_33596_, _33595_, _33594_);
  nand (_33597_, _33596_, _35583_);
  or (_33598_, \oc8051_gm_cxrom_1.cell11.data [2], _35583_);
  and (_35588_[2], _33598_, _33597_);
  or (_33599_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33600_, \oc8051_gm_cxrom_1.cell11.data [3], _33579_);
  nand (_33601_, _33600_, _33599_);
  nand (_33602_, _33601_, _35583_);
  or (_33603_, \oc8051_gm_cxrom_1.cell11.data [3], _35583_);
  and (_35588_[3], _33603_, _33602_);
  or (_33604_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33605_, \oc8051_gm_cxrom_1.cell11.data [4], _33579_);
  nand (_33606_, _33605_, _33604_);
  nand (_33607_, _33606_, _35583_);
  or (_33608_, \oc8051_gm_cxrom_1.cell11.data [4], _35583_);
  and (_35588_[4], _33608_, _33607_);
  or (_33609_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33610_, \oc8051_gm_cxrom_1.cell11.data [5], _33579_);
  nand (_33611_, _33610_, _33609_);
  nand (_33612_, _33611_, _35583_);
  or (_33613_, \oc8051_gm_cxrom_1.cell11.data [5], _35583_);
  and (_35588_[5], _33613_, _33612_);
  or (_33614_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or (_33615_, \oc8051_gm_cxrom_1.cell11.data [6], _33579_);
  nand (_33616_, _33615_, _33614_);
  nand (_33617_, _33616_, _35583_);
  or (_33618_, \oc8051_gm_cxrom_1.cell11.data [6], _35583_);
  and (_35588_[6], _33618_, _33617_);
  or (_33619_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not (_33620_, \oc8051_gm_cxrom_1.cell12.valid );
  or (_33621_, _33620_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand (_33622_, _33621_, _33619_);
  nand (_33623_, _33622_, _35583_);
  or (_33624_, \oc8051_gm_cxrom_1.cell12.data [7], _35583_);
  and (_35590_[7], _33624_, _33623_);
  or (_33625_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33626_, \oc8051_gm_cxrom_1.cell12.data [0], _33620_);
  nand (_33627_, _33626_, _33625_);
  nand (_33628_, _33627_, _35583_);
  or (_33629_, \oc8051_gm_cxrom_1.cell12.data [0], _35583_);
  and (_35590_[0], _33629_, _33628_);
  or (_33630_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33631_, \oc8051_gm_cxrom_1.cell12.data [1], _33620_);
  nand (_33632_, _33631_, _33630_);
  nand (_33633_, _33632_, _35583_);
  or (_33634_, \oc8051_gm_cxrom_1.cell12.data [1], _35583_);
  and (_35590_[1], _33634_, _33633_);
  or (_33635_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33636_, \oc8051_gm_cxrom_1.cell12.data [2], _33620_);
  nand (_33637_, _33636_, _33635_);
  nand (_33638_, _33637_, _35583_);
  or (_33639_, \oc8051_gm_cxrom_1.cell12.data [2], _35583_);
  and (_35590_[2], _33639_, _33638_);
  or (_33640_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33641_, \oc8051_gm_cxrom_1.cell12.data [3], _33620_);
  nand (_33642_, _33641_, _33640_);
  nand (_33643_, _33642_, _35583_);
  or (_33644_, \oc8051_gm_cxrom_1.cell12.data [3], _35583_);
  and (_35590_[3], _33644_, _33643_);
  or (_33645_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33646_, \oc8051_gm_cxrom_1.cell12.data [4], _33620_);
  nand (_33647_, _33646_, _33645_);
  nand (_33648_, _33647_, _35583_);
  or (_33649_, \oc8051_gm_cxrom_1.cell12.data [4], _35583_);
  and (_35590_[4], _33649_, _33648_);
  or (_33650_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33651_, \oc8051_gm_cxrom_1.cell12.data [5], _33620_);
  nand (_33652_, _33651_, _33650_);
  nand (_33653_, _33652_, _35583_);
  or (_33654_, \oc8051_gm_cxrom_1.cell12.data [5], _35583_);
  and (_35590_[5], _33654_, _33653_);
  or (_33655_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or (_33656_, \oc8051_gm_cxrom_1.cell12.data [6], _33620_);
  nand (_33657_, _33656_, _33655_);
  nand (_33658_, _33657_, _35583_);
  or (_33659_, \oc8051_gm_cxrom_1.cell12.data [6], _35583_);
  and (_35590_[6], _33659_, _33658_);
  or (_33660_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not (_33661_, \oc8051_gm_cxrom_1.cell13.valid );
  or (_33662_, _33661_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand (_33663_, _33662_, _33660_);
  nand (_33664_, _33663_, _35583_);
  or (_33665_, \oc8051_gm_cxrom_1.cell13.data [7], _35583_);
  and (_35592_[7], _33665_, _33664_);
  or (_33666_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33667_, \oc8051_gm_cxrom_1.cell13.data [0], _33661_);
  nand (_33668_, _33667_, _33666_);
  nand (_33669_, _33668_, _35583_);
  or (_33670_, \oc8051_gm_cxrom_1.cell13.data [0], _35583_);
  and (_35592_[0], _33670_, _33669_);
  or (_33671_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33672_, \oc8051_gm_cxrom_1.cell13.data [1], _33661_);
  nand (_33673_, _33672_, _33671_);
  nand (_33674_, _33673_, _35583_);
  or (_33675_, \oc8051_gm_cxrom_1.cell13.data [1], _35583_);
  and (_35592_[1], _33675_, _33674_);
  or (_33676_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33677_, \oc8051_gm_cxrom_1.cell13.data [2], _33661_);
  nand (_33678_, _33677_, _33676_);
  nand (_33679_, _33678_, _35583_);
  or (_33680_, \oc8051_gm_cxrom_1.cell13.data [2], _35583_);
  and (_35592_[2], _33680_, _33679_);
  or (_33681_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33682_, \oc8051_gm_cxrom_1.cell13.data [3], _33661_);
  nand (_33683_, _33682_, _33681_);
  nand (_33684_, _33683_, _35583_);
  or (_33685_, \oc8051_gm_cxrom_1.cell13.data [3], _35583_);
  and (_35592_[3], _33685_, _33684_);
  or (_33686_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33687_, \oc8051_gm_cxrom_1.cell13.data [4], _33661_);
  nand (_33688_, _33687_, _33686_);
  nand (_33689_, _33688_, _35583_);
  or (_33690_, \oc8051_gm_cxrom_1.cell13.data [4], _35583_);
  and (_35592_[4], _33690_, _33689_);
  or (_33691_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33692_, \oc8051_gm_cxrom_1.cell13.data [5], _33661_);
  nand (_33693_, _33692_, _33691_);
  nand (_33694_, _33693_, _35583_);
  or (_33695_, \oc8051_gm_cxrom_1.cell13.data [5], _35583_);
  and (_35592_[5], _33695_, _33694_);
  or (_33696_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or (_33697_, \oc8051_gm_cxrom_1.cell13.data [6], _33661_);
  nand (_33698_, _33697_, _33696_);
  nand (_33699_, _33698_, _35583_);
  or (_33700_, \oc8051_gm_cxrom_1.cell13.data [6], _35583_);
  and (_35592_[6], _33700_, _33699_);
  or (_33701_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not (_33702_, \oc8051_gm_cxrom_1.cell14.valid );
  or (_33703_, _33702_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand (_33704_, _33703_, _33701_);
  nand (_33705_, _33704_, _35583_);
  or (_33706_, \oc8051_gm_cxrom_1.cell14.data [7], _35583_);
  and (_35594_[7], _33706_, _33705_);
  or (_33707_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33708_, \oc8051_gm_cxrom_1.cell14.data [0], _33702_);
  nand (_33709_, _33708_, _33707_);
  nand (_33710_, _33709_, _35583_);
  or (_33711_, \oc8051_gm_cxrom_1.cell14.data [0], _35583_);
  and (_35594_[0], _33711_, _33710_);
  or (_33712_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33713_, \oc8051_gm_cxrom_1.cell14.data [1], _33702_);
  nand (_33714_, _33713_, _33712_);
  nand (_33715_, _33714_, _35583_);
  or (_33716_, \oc8051_gm_cxrom_1.cell14.data [1], _35583_);
  and (_35594_[1], _33716_, _33715_);
  or (_33717_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33718_, \oc8051_gm_cxrom_1.cell14.data [2], _33702_);
  nand (_33719_, _33718_, _33717_);
  nand (_33720_, _33719_, _35583_);
  or (_33721_, \oc8051_gm_cxrom_1.cell14.data [2], _35583_);
  and (_35594_[2], _33721_, _33720_);
  or (_33722_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33723_, \oc8051_gm_cxrom_1.cell14.data [3], _33702_);
  nand (_33724_, _33723_, _33722_);
  nand (_33725_, _33724_, _35583_);
  or (_33726_, \oc8051_gm_cxrom_1.cell14.data [3], _35583_);
  and (_35594_[3], _33726_, _33725_);
  or (_33727_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33728_, \oc8051_gm_cxrom_1.cell14.data [4], _33702_);
  nand (_33729_, _33728_, _33727_);
  nand (_33730_, _33729_, _35583_);
  or (_33731_, \oc8051_gm_cxrom_1.cell14.data [4], _35583_);
  and (_35594_[4], _33731_, _33730_);
  or (_33732_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33733_, \oc8051_gm_cxrom_1.cell14.data [5], _33702_);
  nand (_33734_, _33733_, _33732_);
  nand (_33735_, _33734_, _35583_);
  or (_33736_, \oc8051_gm_cxrom_1.cell14.data [5], _35583_);
  and (_35594_[5], _33736_, _33735_);
  or (_33737_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or (_33738_, \oc8051_gm_cxrom_1.cell14.data [6], _33702_);
  nand (_33739_, _33738_, _33737_);
  nand (_33740_, _33739_, _35583_);
  or (_33741_, \oc8051_gm_cxrom_1.cell14.data [6], _35583_);
  and (_35594_[6], _33741_, _33740_);
  or (_33742_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not (_33743_, \oc8051_gm_cxrom_1.cell15.valid );
  or (_33744_, _33743_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand (_33745_, _33744_, _33742_);
  nand (_33746_, _33745_, _35583_);
  or (_33747_, \oc8051_gm_cxrom_1.cell15.data [7], _35583_);
  and (_35596_[7], _33747_, _33746_);
  or (_33748_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33749_, \oc8051_gm_cxrom_1.cell15.data [0], _33743_);
  nand (_33750_, _33749_, _33748_);
  nand (_33751_, _33750_, _35583_);
  or (_33752_, \oc8051_gm_cxrom_1.cell15.data [0], _35583_);
  and (_35596_[0], _33752_, _33751_);
  or (_33753_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33754_, \oc8051_gm_cxrom_1.cell15.data [1], _33743_);
  nand (_33755_, _33754_, _33753_);
  nand (_33756_, _33755_, _35583_);
  or (_33757_, \oc8051_gm_cxrom_1.cell15.data [1], _35583_);
  and (_35596_[1], _33757_, _33756_);
  or (_33758_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33759_, \oc8051_gm_cxrom_1.cell15.data [2], _33743_);
  nand (_33760_, _33759_, _33758_);
  nand (_33761_, _33760_, _35583_);
  or (_33762_, \oc8051_gm_cxrom_1.cell15.data [2], _35583_);
  and (_35596_[2], _33762_, _33761_);
  or (_33763_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33764_, \oc8051_gm_cxrom_1.cell15.data [3], _33743_);
  nand (_33765_, _33764_, _33763_);
  nand (_33766_, _33765_, _35583_);
  or (_33767_, \oc8051_gm_cxrom_1.cell15.data [3], _35583_);
  and (_35596_[3], _33767_, _33766_);
  or (_33768_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33769_, \oc8051_gm_cxrom_1.cell15.data [4], _33743_);
  nand (_33770_, _33769_, _33768_);
  nand (_33771_, _33770_, _35583_);
  or (_33772_, \oc8051_gm_cxrom_1.cell15.data [4], _35583_);
  and (_35596_[4], _33772_, _33771_);
  or (_33773_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33774_, \oc8051_gm_cxrom_1.cell15.data [5], _33743_);
  nand (_33775_, _33774_, _33773_);
  nand (_33776_, _33775_, _35583_);
  or (_33777_, \oc8051_gm_cxrom_1.cell15.data [5], _35583_);
  and (_35596_[5], _33777_, _33776_);
  or (_33778_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or (_33779_, \oc8051_gm_cxrom_1.cell15.data [6], _33743_);
  nand (_33780_, _33779_, _33778_);
  nand (_33781_, _33780_, _35583_);
  or (_33782_, \oc8051_gm_cxrom_1.cell15.data [6], _35583_);
  and (_35596_[6], _33782_, _33781_);
  nor (_35779_[2], _30720_, rst);
  and (_33783_, _30335_, _35583_);
  nand (_33784_, _33783_, _30556_);
  nor (_33785_, _30588_, _30547_);
  or (_35780_[2], _33785_, _33784_);
  not (_33786_, _30416_);
  and (_33787_, _33786_, _30394_);
  not (_33788_, _30509_);
  not (_33789_, _30487_);
  nor (_33790_, _33789_, _30464_);
  and (_33791_, _33790_, _30442_);
  and (_33792_, _33791_, _30540_);
  and (_33793_, _33792_, _33788_);
  and (_33794_, _33793_, _33787_);
  not (_33795_, _30394_);
  and (_33796_, _30416_, _33795_);
  and (_33797_, _30487_, _30464_);
  and (_33798_, _33797_, _30442_);
  and (_33799_, _33798_, _30540_);
  and (_33800_, _33799_, _30509_);
  and (_33801_, _33800_, _33796_);
  or (_33802_, _33801_, _33794_);
  not (_33803_, _30442_);
  and (_33804_, _33797_, _33803_);
  nor (_33805_, _30370_, _30509_);
  nor (_33806_, _30416_, _30394_);
  and (_33807_, _33806_, _33805_);
  and (_33808_, _33807_, _33804_);
  nor (_33809_, _30370_, _33788_);
  and (_33810_, _33809_, _33787_);
  and (_33811_, _33810_, _33791_);
  or (_33812_, _33811_, _33808_);
  and (_33813_, _33806_, _33809_);
  and (_33814_, _33813_, _33804_);
  nor (_33815_, _33788_, _30487_);
  and (_33816_, _33806_, _30370_);
  and (_33817_, _33816_, _33815_);
  or (_33818_, _33817_, _33814_);
  or (_33819_, _33818_, _33812_);
  and (_33820_, _33787_, _30370_);
  not (_33821_, _30540_);
  and (_33822_, _33804_, _33821_);
  and (_33823_, _33822_, _33820_);
  not (_33824_, _30370_);
  and (_33825_, _33806_, _33824_);
  and (_33826_, _33825_, _33799_);
  or (_33827_, _33826_, _33823_);
  or (_33828_, _33827_, _33819_);
  or (_33829_, _33828_, _33802_);
  and (_33830_, _30370_, _33788_);
  and (_33831_, _33796_, _33830_);
  and (_33832_, _33831_, _33799_);
  and (_33833_, _30416_, _30394_);
  and (_33834_, _33833_, _33809_);
  and (_33835_, _33834_, _33799_);
  not (_33836_, _33798_);
  and (_33837_, _33796_, _33805_);
  nor (_33838_, _33837_, _33821_);
  nor (_33839_, _33838_, _33836_);
  or (_33840_, _33839_, _33835_);
  nor (_33841_, _33840_, _33832_);
  and (_33842_, _33804_, _30540_);
  and (_33843_, _33833_, _30370_);
  and (_33844_, _33843_, _33842_);
  and (_33845_, _33833_, _33824_);
  and (_33846_, _33842_, _33845_);
  and (_33847_, _33787_, _33824_);
  nor (_33848_, _33788_, _30442_);
  and (_33849_, _33848_, _33790_);
  or (_33850_, _33849_, _33815_);
  and (_33851_, _33850_, _33847_);
  or (_33852_, _33851_, _33846_);
  or (_33853_, _33852_, _33844_);
  and (_33854_, _33809_, _33796_);
  and (_33855_, _33822_, _33854_);
  and (_33856_, _30370_, _30509_);
  and (_33857_, _33806_, _33856_);
  and (_33858_, _33791_, _33821_);
  and (_33859_, _33858_, _33857_);
  or (_33860_, _33859_, _33855_);
  nor (_33861_, _33856_, _33805_);
  not (_33862_, _33861_);
  and (_33863_, _33862_, _33833_);
  and (_33864_, _33863_, _33799_);
  and (_33865_, _33830_, _33787_);
  and (_33866_, _33799_, _33865_);
  or (_33867_, _33866_, _33864_);
  or (_33868_, _33867_, _33860_);
  nor (_33869_, _33868_, _33853_);
  nand (_33870_, _33869_, _33841_);
  or (_33871_, _33870_, _33829_);
  and (_33872_, _33871_, _30336_);
  not (_33873_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_33874_, _30334_, _15093_);
  and (_33875_, _33874_, _30601_);
  nor (_33876_, _33875_, _33873_);
  or (_33877_, _33876_, rst);
  or (_35781_[1], _33877_, _33872_);
  nand (_33878_, _30416_, _30330_);
  or (_33879_, _30330_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_33880_, _33879_, _35583_);
  and (_35782_[7], _33880_, _33878_);
  and (_33881_, \oc8051_top_1.oc8051_sfr1.wait_data , _35583_);
  and (_33882_, _33881_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  or (_33883_, _30692_, _30627_);
  and (_33884_, _30626_, _30575_);
  and (_33885_, _30594_, _30588_);
  and (_33886_, _30586_, _30547_);
  or (_33887_, _33886_, _33885_);
  or (_33888_, _33887_, _33884_);
  or (_33889_, _33888_, _33883_);
  not (_33890_, _30675_);
  and (_33891_, _30709_, _30656_);
  and (_33892_, _30575_, _30563_);
  and (_33893_, _33892_, _30513_);
  or (_33894_, _33893_, _33891_);
  or (_33895_, _33894_, _33890_);
  or (_33896_, _33895_, _33889_);
  and (_33897_, _33896_, _33783_);
  or (_35783_, _33897_, _33882_);
  and (_33898_, _30552_, _30374_);
  nor (_33899_, _30514_, _30491_);
  and (_33900_, _33899_, _33898_);
  and (_33901_, _33900_, _30421_);
  or (_33902_, _33901_, _30562_);
  and (_33903_, _30614_, _30446_);
  and (_33904_, _33903_, _30626_);
  or (_33905_, _33904_, _33902_);
  and (_33906_, _30588_, _30582_);
  or (_33907_, _33906_, _30576_);
  or (_33908_, _33907_, _33905_);
  and (_33909_, _33908_, _30335_);
  and (_33910_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_33911_, \oc8051_top_1.oc8051_decoder1.state [0], _15093_);
  and (_33912_, _33911_, _33873_);
  not (_33913_, _30712_);
  and (_33914_, _33913_, _33912_);
  or (_33915_, _33914_, _33910_);
  or (_33916_, _33915_, _33909_);
  and (_35784_[1], _33916_, _35583_);
  and (_33917_, _33881_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_33918_, _30709_, _30676_);
  nor (_33919_, _30676_, _30586_);
  nor (_33920_, _33919_, _30654_);
  or (_33921_, _33920_, _33918_);
  and (_33922_, _33903_, _30632_);
  or (_33923_, _33922_, _33921_);
  not (_33924_, _30522_);
  nor (_33925_, _33919_, _30491_);
  nor (_33926_, _30513_, _30491_);
  and (_33927_, _33926_, _30520_);
  or (_33928_, _33927_, _33925_);
  or (_33929_, _33928_, _33924_);
  and (_33930_, _30709_, _30650_);
  and (_33931_, _30624_, _30680_);
  or (_33932_, _33931_, _33930_);
  or (_33933_, _33932_, _33907_);
  or (_33934_, _33933_, _33929_);
  or (_33935_, _33934_, _33923_);
  and (_33936_, _33935_, _33783_);
  or (_35785_[1], _33936_, _33917_);
  and (_33937_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_33938_, _30643_, _30335_);
  or (_33939_, _33938_, _33937_);
  or (_33940_, _33939_, _33914_);
  and (_35786_[2], _33940_, _35583_);
  not (_33941_, _33785_);
  and (_33942_, _33941_, _30656_);
  nor (_33943_, _33942_, _33892_);
  not (_33944_, _33943_);
  and (_33945_, _33944_, _33912_);
  or (_33946_, _33945_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_33947_, _30615_, _30546_);
  and (_33948_, _30548_, _30520_);
  nor (_33949_, _33948_, _33947_);
  nor (_33950_, _33949_, _30513_);
  not (_33951_, _30331_);
  and (_33952_, _33893_, _33951_);
  or (_33953_, _33952_, _33950_);
  and (_33954_, _33953_, _30601_);
  or (_33955_, _33954_, _33946_);
  or (_33956_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _15093_);
  and (_33957_, _33956_, _35583_);
  and (_35787_[2], _33957_, _33955_);
  and (_33958_, _33881_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  and (_33959_, _33926_, _30561_);
  or (_33960_, _33927_, _33959_);
  or (_33961_, _30617_, _30576_);
  or (_33962_, _33961_, _33960_);
  and (_33963_, _30548_, _30423_);
  or (_33964_, _33922_, _33886_);
  or (_33965_, _33964_, _33963_);
  or (_33966_, _30632_, _30626_);
  and (_33967_, _33966_, _30518_);
  or (_33968_, _33901_, _30665_);
  or (_33969_, _33968_, _33967_);
  or (_33970_, _33969_, _33965_);
  or (_33971_, _33970_, _33962_);
  and (_33972_, _33971_, _33783_);
  or (_35788_[1], _33972_, _33958_);
  and (_33973_, _33881_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  or (_33974_, _33904_, _30634_);
  and (_33975_, _30575_, _30519_);
  and (_33976_, _33903_, _30591_);
  or (_33977_, _33976_, _33975_);
  or (_33978_, _33977_, _33974_);
  or (_33979_, _33978_, _33928_);
  and (_33980_, _30561_, _30516_);
  and (_33981_, _33898_, _30551_);
  or (_33982_, _33981_, _30592_);
  or (_33983_, _33982_, _33980_);
  not (_33984_, _30622_);
  and (_33985_, _30709_, _30620_);
  or (_33986_, _33985_, _33984_);
  or (_33987_, _33986_, _33983_);
  or (_33988_, _33987_, _33979_);
  nor (_33989_, _30640_, _30521_);
  not (_33990_, _30631_);
  and (_33991_, _33899_, _30579_);
  or (_33992_, _33991_, _33900_);
  nor (_33993_, _33992_, _33990_);
  nand (_33994_, _33993_, _33989_);
  or (_33995_, _33994_, _33923_);
  or (_33996_, _33995_, _33988_);
  and (_33997_, _33996_, _33783_);
  or (_35789_[3], _33997_, _33973_);
  and (_33998_, _30582_, _30518_);
  and (_33999_, _33926_, _30563_);
  and (_34000_, _30549_, _30680_);
  and (_34001_, _30549_, _30518_);
  and (_34002_, _33903_, _30549_);
  or (_34003_, _34002_, _34001_);
  or (_34004_, _34003_, _34000_);
  or (_34005_, _34004_, _33999_);
  or (_34006_, _34005_, _33998_);
  and (_34007_, _30616_, _30582_);
  and (_34008_, _30709_, _30582_);
  or (_34009_, _34008_, _34007_);
  or (_34010_, _34009_, _34006_);
  and (_34011_, _34010_, _30335_);
  and (_34012_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_34013_, _34012_, _30717_);
  or (_34014_, _34013_, _34011_);
  and (_35790_[1], _34014_, _35583_);
  or (_34015_, _30665_, _30661_);
  not (_34016_, _30628_);
  or (_34017_, _33920_, _34016_);
  or (_34018_, _34017_, _34015_);
  and (_34019_, _30578_, _30514_);
  and (_34020_, _34019_, _30616_);
  or (_34021_, _34020_, _30633_);
  and (_34022_, _30632_, _30548_);
  or (_34023_, _34022_, _30621_);
  nor (_34024_, _34023_, _34021_);
  nand (_34025_, _34024_, _30645_);
  or (_34026_, _34025_, _34018_);
  and (_34027_, _34019_, _30518_);
  or (_34028_, _34027_, _30521_);
  or (_34029_, _34028_, _30679_);
  and (_34030_, _33926_, _30578_);
  or (_34031_, _34030_, _30647_);
  and (_34032_, _33947_, _30514_);
  or (_34033_, _34032_, _30595_);
  or (_34034_, _34033_, _34031_);
  or (_34035_, _34034_, _34029_);
  and (_34036_, _33899_, _30563_);
  or (_34037_, _33902_, _30681_);
  or (_34038_, _34037_, _34036_);
  or (_34039_, _34038_, _33928_);
  or (_34040_, _34039_, _34035_);
  or (_34041_, _34040_, _34026_);
  and (_34042_, _34041_, _30335_);
  and (_34043_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_34044_, _30698_, _30603_);
  or (_34045_, _34022_, _34032_);
  and (_34046_, _34045_, _30603_);
  or (_34047_, _34046_, _33914_);
  or (_34048_, _34047_, _34044_);
  or (_34049_, _34048_, _34043_);
  or (_34050_, _34049_, _34042_);
  and (_35791_, _34050_, _35583_);
  nor (_35779_[0], _30609_, rst);
  nor (_35779_[1], _30704_, rst);
  nand (_35780_[0], _33944_, _33783_);
  nand (_34051_, _33892_, _33783_);
  or (_34052_, _33784_, _30671_);
  and (_35780_[1], _34052_, _34051_);
  or (_34053_, _33823_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_34054_, _34053_, _33846_);
  or (_34055_, _34054_, _33794_);
  and (_34056_, _34055_, _33875_);
  nor (_34057_, _33874_, _30601_);
  or (_34058_, _34057_, rst);
  or (_35781_[0], _34058_, _34056_);
  nand (_34059_, _30540_, _30330_);
  or (_34060_, _30330_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_34061_, _34060_, _35583_);
  and (_35782_[0], _34061_, _34059_);
  nand (_34062_, _30442_, _30330_);
  or (_34063_, _30330_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_34064_, _34063_, _35583_);
  and (_35782_[1], _34064_, _34062_);
  nand (_34065_, _30464_, _30330_);
  or (_34066_, _30330_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_34067_, _34066_, _35583_);
  and (_35782_[2], _34067_, _34065_);
  nand (_34068_, _30487_, _30330_);
  or (_34069_, _30330_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_34070_, _34069_, _35583_);
  and (_35782_[3], _34070_, _34068_);
  or (_34071_, _30509_, _30716_);
  or (_34072_, _30330_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_34073_, _34072_, _35583_);
  and (_35782_[4], _34073_, _34071_);
  nand (_34074_, _30370_, _30330_);
  or (_34075_, _30330_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_34076_, _34075_, _35583_);
  and (_35782_[5], _34076_, _34074_);
  nand (_34077_, _30394_, _30330_);
  or (_34078_, _30330_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_34079_, _34078_, _35583_);
  and (_35782_[6], _34079_, _34077_);
  or (_34080_, _33906_, _30629_);
  or (_34081_, _34080_, _33985_);
  and (_34082_, _30556_, _30514_);
  and (_34083_, _34082_, _30709_);
  and (_34084_, _30709_, _30580_);
  and (_34085_, _33926_, _30554_);
  or (_34086_, _34085_, _34084_);
  or (_34087_, _34086_, _34083_);
  or (_34088_, _34087_, _34005_);
  or (_34089_, _34088_, _34081_);
  or (_34090_, _30592_, _33998_);
  or (_34091_, _30657_, _30576_);
  or (_34092_, _34091_, _34090_);
  or (_34093_, _30586_, _30520_);
  and (_34094_, _34093_, _30709_);
  and (_34095_, _33899_, _30554_);
  or (_34096_, _34095_, _30558_);
  or (_34097_, _34096_, _34094_);
  or (_34098_, _34097_, _34092_);
  and (_34099_, _33903_, _30582_);
  and (_34100_, _33903_, _30568_);
  or (_34101_, _34100_, _34099_);
  and (_34102_, _30656_, _30680_);
  and (_34103_, _30568_, _30518_);
  or (_34104_, _34103_, _34102_);
  or (_34105_, _34104_, _34101_);
  or (_34106_, _33991_, _33891_);
  or (_34107_, _34106_, _33977_);
  or (_34108_, _34107_, _34105_);
  or (_34109_, _34108_, _34098_);
  or (_34110_, _34109_, _34089_);
  and (_34111_, _34110_, _30335_);
  and (_34112_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34113_, _34112_, _33945_);
  or (_34114_, _34113_, _34111_);
  and (_35784_[0], _34114_, _35583_);
  and (_34115_, _33881_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_34116_, _30620_, _30591_);
  and (_34117_, _34116_, _30548_);
  or (_34118_, _34117_, _33992_);
  and (_34119_, _30398_, _30375_);
  and (_34120_, _33926_, _34119_);
  and (_34121_, _34120_, _30421_);
  nor (_34122_, _34121_, _30517_);
  not (_34123_, _30709_);
  or (_34124_, _34123_, _30569_);
  nand (_34125_, _34124_, _34122_);
  or (_34126_, _34125_, _34118_);
  or (_34127_, _34081_, _33983_);
  and (_34128_, _30709_, _30591_);
  nor (_34129_, _34128_, _33930_);
  nand (_34130_, _34129_, _30666_);
  or (_34131_, _34130_, _33894_);
  or (_34132_, _34131_, _34127_);
  or (_34133_, _34132_, _34126_);
  and (_34134_, _34133_, _33783_);
  or (_35785_[0], _34134_, _34115_);
  or (_34135_, _34036_, _30647_);
  or (_34136_, _34135_, _34033_);
  or (_34137_, _34136_, _34026_);
  and (_34138_, _34137_, _30335_);
  and (_34139_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34140_, _34139_, _34048_);
  or (_34141_, _34140_, _34138_);
  and (_35786_[0], _34141_, _35583_);
  and (_34142_, _30639_, _30513_);
  or (_34143_, _34142_, _30562_);
  or (_34144_, _34143_, _34029_);
  or (_34145_, _34144_, _33950_);
  and (_34146_, _34145_, _30335_);
  and (_34147_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34148_, _34147_, _34047_);
  or (_34149_, _34148_, _34146_);
  and (_35786_[1], _34149_, _35583_);
  and (_34150_, _30568_, _30548_);
  and (_34151_, _34020_, _30421_);
  or (_34152_, _34151_, _34128_);
  or (_34153_, _34152_, _34150_);
  or (_34154_, _34153_, _33950_);
  and (_34155_, _30554_, _30516_);
  or (_34156_, _34001_, _34155_);
  or (_34157_, _33999_, _34156_);
  or (_34158_, _33892_, _30711_);
  and (_34159_, _34002_, _30514_);
  or (_34160_, _34159_, _34100_);
  or (_34161_, _34160_, _34158_);
  or (_34162_, _34161_, _34157_);
  or (_34163_, _34162_, _34154_);
  and (_34164_, _33903_, _30624_);
  or (_34165_, _34164_, _33891_);
  or (_34166_, _34083_, _30710_);
  or (_34167_, _34166_, _34094_);
  or (_34168_, _34167_, _34165_);
  or (_34169_, _34085_, _34000_);
  and (_34170_, _30709_, _30626_);
  or (_34171_, _34099_, _33975_);
  or (_34172_, _34171_, _34170_);
  or (_34173_, _34172_, _34169_);
  and (_34174_, _34002_, _30513_);
  or (_34175_, _34174_, _30581_);
  or (_34176_, _34030_, _34027_);
  or (_34177_, _34176_, _33998_);
  or (_34178_, _34084_, _33985_);
  or (_34179_, _34178_, _34177_);
  or (_34180_, _34179_, _34175_);
  or (_34181_, _34180_, _34173_);
  or (_34182_, _34181_, _34168_);
  or (_34183_, _34182_, _34163_);
  and (_34184_, _34183_, _30335_);
  and (_34185_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34186_, _33945_, _30718_);
  or (_34187_, _34186_, _34185_);
  or (_34188_, _34187_, _34184_);
  and (_35787_[0], _34188_, _35583_);
  or (_34189_, _30640_, _30621_);
  and (_34190_, _34189_, _30574_);
  or (_34191_, _30711_, _30647_);
  and (_34192_, _30556_, _30516_);
  or (_34193_, _34192_, _33906_);
  or (_34194_, _34193_, _34191_);
  or (_34195_, _34194_, _34157_);
  or (_34196_, _34195_, _34190_);
  and (_34197_, _33926_, _30556_);
  or (_34198_, _34197_, _34020_);
  nor (_34199_, _34198_, _33998_);
  nand (_34200_, _34199_, _30584_);
  or (_34201_, _34200_, _30655_);
  or (_34202_, _34201_, _34173_);
  or (_34203_, _34202_, _34168_);
  or (_34204_, _34203_, _34196_);
  and (_34205_, _34204_, _30335_);
  and (_34206_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34207_, _34206_, _34186_);
  or (_34208_, _34207_, _34205_);
  and (_35787_[1], _34208_, _35583_);
  and (_34209_, _33881_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_34210_, _34001_, _30514_);
  and (_34211_, _30575_, _30624_);
  and (_34212_, _30575_, _30672_);
  or (_34213_, _34212_, _34211_);
  or (_34214_, _34213_, _34210_);
  or (_34215_, _34214_, _33962_);
  and (_34216_, _30575_, _30520_);
  and (_34217_, _34216_, _30514_);
  and (_34218_, _33886_, _30574_);
  or (_34219_, _34218_, _34217_);
  not (_34220_, _31856_);
  or (_34221_, _34099_, _34220_);
  or (_34222_, _34221_, _34219_);
  or (_34223_, _34222_, _34215_);
  or (_34224_, _33999_, _33901_);
  and (_34225_, _30709_, _30586_);
  or (_34226_, _34225_, _33922_);
  or (_34227_, _34226_, _34015_);
  or (_34228_, _34227_, _34224_);
  and (_34229_, _33926_, _30549_);
  or (_34230_, _34229_, _33998_);
  or (_34231_, _34159_, _30642_);
  or (_34232_, _34231_, _34230_);
  not (_34233_, _31855_);
  or (_34234_, _33967_, _34233_);
  or (_34235_, _34234_, _34232_);
  or (_34236_, _34235_, _34228_);
  or (_34237_, _34236_, _34223_);
  and (_34238_, _34237_, _33783_);
  or (_35788_[0], _34238_, _34209_);
  or (_34239_, _33904_, _30629_);
  or (_34240_, _33981_, _33980_);
  or (_34241_, _34240_, _34239_);
  or (_34242_, _34241_, _33986_);
  or (_34243_, _34242_, _34161_);
  or (_34244_, _34212_, _34225_);
  or (_34245_, _34217_, _34169_);
  or (_34246_, _34245_, _34244_);
  or (_34247_, _33900_, _31945_);
  or (_34248_, _34247_, _30576_);
  or (_34249_, _34248_, _30570_);
  or (_34250_, _34175_, _30649_);
  or (_34251_, _34250_, _34249_);
  or (_34252_, _34251_, _34246_);
  or (_34253_, _34252_, _34243_);
  or (_34254_, _30711_, _33951_);
  or (_34255_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _15093_);
  and (_34256_, _34255_, _35583_);
  and (_34257_, _34256_, _34254_);
  and (_35789_[0], _34257_, _34253_);
  and (_34258_, _30575_, _30549_);
  or (_34259_, _34099_, _33931_);
  or (_34260_, _34259_, _34258_);
  or (_34261_, _30630_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_34262_, _33904_, _30711_);
  or (_34263_, _34262_, _34261_);
  or (_34264_, _34263_, _34260_);
  or (_34265_, _34083_, _30625_);
  or (_34266_, _34265_, _34211_);
  not (_34267_, _30646_);
  nor (_34268_, _34100_, _30647_);
  and (_34269_, _34268_, _34267_);
  not (_34270_, _34269_);
  or (_34271_, _34270_, _34266_);
  or (_34272_, _34271_, _34264_);
  or (_34273_, _34165_, _30566_);
  or (_34274_, _34085_, _34155_);
  or (_34275_, _34274_, _34224_);
  or (_34276_, _34275_, _34273_);
  or (_34277_, _34276_, _33929_);
  or (_34278_, _34277_, _33923_);
  or (_34279_, _34278_, _34272_);
  or (_34280_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _15093_);
  and (_34281_, _34280_, _35583_);
  and (_34282_, _34281_, _34254_);
  and (_35789_[1], _34282_, _34279_);
  or (_34283_, _34226_, _33968_);
  not (_34284_, _34268_);
  or (_34285_, _34274_, _34284_);
  or (_34286_, _34285_, _34283_);
  or (_34287_, _30562_, _30521_);
  nor (_34288_, _34287_, _34216_);
  nand (_34289_, _34288_, _31856_);
  or (_34290_, _34289_, _33928_);
  or (_34291_, _34266_, _33921_);
  or (_34292_, _34291_, _34290_);
  or (_34293_, _34292_, _34286_);
  and (_34294_, _34293_, _30335_);
  and (_34295_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_34296_, _30710_, _15093_);
  or (_34297_, _34296_, _34295_);
  or (_34298_, _34297_, _34294_);
  and (_35789_[2], _34298_, _35583_);
  and (_34299_, _33881_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_34300_, _33884_, _30662_);
  nand (_34301_, _34300_, _31855_);
  not (_34302_, _30546_);
  or (_34303_, _30575_, _34302_);
  and (_34304_, _34303_, _30624_);
  or (_34305_, _34304_, _34244_);
  or (_34306_, _34305_, _34301_);
  or (_34307_, _34306_, _34222_);
  or (_34308_, _34307_, _34006_);
  and (_34309_, _34308_, _33783_);
  or (_35790_[0], _34309_, _34299_);
  nor (_35776_[7], _30416_, rst);
  nor (_35777_[7], _32030_, rst);
  nor (_34310_, _30426_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and (_34311_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_34312_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_34313_, _34312_, _34311_);
  and (_34314_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_34315_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_34316_, _34315_, _34314_);
  and (_34317_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_34318_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_34319_, _34318_, _34317_);
  and (_34320_, _34319_, _34316_);
  and (_34321_, _34320_, _34313_);
  and (_34322_, _34321_, _30426_);
  nor (_34323_, _34322_, _34310_);
  nor (_34324_, _34323_, _31945_);
  nor (_34325_, _30335_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  nor (_34326_, _34325_, _34324_);
  and (_35778_[7], _34326_, _35583_);
  nor (_35776_[0], _30540_, rst);
  nor (_35776_[1], _30442_, rst);
  nor (_35776_[2], _30464_, rst);
  nor (_35776_[3], _30487_, rst);
  and (_35776_[4], _30509_, _35583_);
  nor (_35776_[5], _30370_, rst);
  nor (_35776_[6], _30394_, rst);
  nor (_35777_[0], _31961_, rst);
  nor (_35777_[1], _32241_, rst);
  nor (_35777_[2], _32134_, rst);
  nor (_35777_[3], _32081_, rst);
  nor (_35777_[4], _32290_, rst);
  nor (_35777_[5], _32186_, rst);
  nor (_35777_[6], _32352_, rst);
  nor (_34327_, _30426_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and (_34328_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_34329_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_34330_, _34329_, _34328_);
  and (_34331_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_34332_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_34333_, _34332_, _34331_);
  and (_34334_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_34335_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_34336_, _34335_, _34334_);
  and (_34337_, _34336_, _34333_);
  and (_34338_, _34337_, _34330_);
  and (_34339_, _34338_, _30426_);
  nor (_34340_, _34339_, _34327_);
  nor (_34341_, _34340_, _31945_);
  nor (_34342_, _30335_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  nor (_34343_, _34342_, _34341_);
  and (_35778_[0], _34343_, _35583_);
  nor (_34344_, _30426_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and (_34345_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_34346_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_34347_, _34346_, _34345_);
  and (_34348_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_34349_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_34350_, _34349_, _34348_);
  and (_34351_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_34352_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_34353_, _34352_, _34351_);
  and (_34354_, _34353_, _34350_);
  and (_34355_, _34354_, _34347_);
  and (_34356_, _34355_, _30426_);
  nor (_34357_, _34356_, _34344_);
  nor (_34358_, _34357_, _31945_);
  nor (_34359_, _30335_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  nor (_34360_, _34359_, _34358_);
  and (_35778_[1], _34360_, _35583_);
  nor (_34361_, _30426_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and (_34362_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_34363_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_34364_, _34363_, _34362_);
  and (_34365_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_34366_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_34367_, _34366_, _34365_);
  and (_34368_, _34367_, _34364_);
  and (_34369_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_34370_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_34371_, _34370_, _34369_);
  and (_34372_, _34371_, _34368_);
  and (_34373_, _34372_, _30426_);
  nor (_34374_, _34373_, _34361_);
  nor (_34375_, _34374_, _31945_);
  nor (_34376_, _30335_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  nor (_34377_, _34376_, _34375_);
  and (_35778_[2], _34377_, _35583_);
  nor (_34378_, _30426_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and (_34379_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_34380_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_34381_, _34380_, _34379_);
  and (_34382_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_34383_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_34384_, _34383_, _34382_);
  and (_34385_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_34386_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_34387_, _34386_, _34385_);
  and (_34388_, _34387_, _34384_);
  and (_34389_, _34388_, _34381_);
  and (_34390_, _34389_, _30426_);
  nor (_34391_, _34390_, _34378_);
  nor (_34392_, _34391_, _31945_);
  nor (_34393_, _30335_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  nor (_34394_, _34393_, _34392_);
  and (_35778_[3], _34394_, _35583_);
  nor (_34395_, _30426_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and (_34396_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_34397_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_34398_, _34397_, _34396_);
  and (_34399_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_34400_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_34401_, _34400_, _34399_);
  and (_34402_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_34403_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_34404_, _34403_, _34402_);
  and (_34405_, _34404_, _34401_);
  and (_34406_, _34405_, _34398_);
  and (_34407_, _34406_, _30426_);
  nor (_34408_, _34407_, _34395_);
  nor (_34409_, _34408_, _31945_);
  nor (_34410_, _30335_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  nor (_34411_, _34410_, _34409_);
  and (_35778_[4], _34411_, _35583_);
  nor (_34412_, _30426_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and (_34413_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_34414_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_34415_, _34414_, _34413_);
  and (_34416_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_34417_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_34418_, _34417_, _34416_);
  and (_34419_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_34420_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_34421_, _34420_, _34419_);
  and (_34422_, _34421_, _34418_);
  and (_34423_, _34422_, _34415_);
  and (_34424_, _34423_, _30426_);
  nor (_34425_, _34424_, _34412_);
  nor (_34426_, _34425_, _31945_);
  nor (_34427_, _30335_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  nor (_34428_, _34427_, _34426_);
  and (_35778_[5], _34428_, _35583_);
  nor (_34429_, _30426_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and (_34430_, _30344_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_34431_, _30348_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_34432_, _34431_, _34430_);
  and (_34433_, _30352_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_34434_, _30356_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_34435_, _34434_, _34433_);
  and (_34436_, _34435_, _34432_);
  and (_34437_, _30360_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_34438_, _30362_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_34439_, _34438_, _34437_);
  and (_34440_, _34439_, _34436_);
  and (_34441_, _34440_, _30426_);
  nor (_34442_, _34441_, _34429_);
  nor (_34443_, _34442_, _31945_);
  nor (_34444_, _30335_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  nor (_34445_, _34444_, _34443_);
  and (_35778_[6], _34445_, _35583_);
  and (_34446_, _30336_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or (_34447_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_34448_, _34446_, _30901_);
  and (_34449_, _34448_, _35583_);
  and (_35793_[15], _34449_, _34447_);
  not (_34450_, _34446_);
  or (_34451_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_00000_, _34446_, _35583_);
  and (_34452_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _35583_);
  or (_34453_, _34452_, _00000_);
  and (_35794_[15], _34453_, _34451_);
  nor (_35795_, _32036_, rst);
  nor (_35796_[4], _32293_, rst);
  and (_35797_[7], _32013_, _35583_);
  nor (_34454_, _32359_, _30725_);
  and (_34455_, _32359_, _30725_);
  nor (_34456_, _34455_, _34454_);
  and (_34457_, _32036_, _28082_);
  nor (_34458_, _32036_, _28082_);
  nor (_34459_, _34458_, _34457_);
  and (_34460_, _34459_, _34456_);
  nor (_34461_, _32191_, _24295_);
  and (_34462_, _32191_, _24295_);
  nor (_34463_, _34462_, _34461_);
  nor (_34464_, _32300_, _31897_);
  and (_34465_, _32300_, _31897_);
  nor (_34466_, _34465_, _34464_);
  and (_34467_, _34466_, _34463_);
  and (_34468_, _34467_, _34460_);
  and (_34469_, _32086_, _24020_);
  nor (_34470_, _32086_, _24020_);
  or (_34471_, _34470_, _34469_);
  not (_34472_, _34471_);
  and (_34473_, _34472_, _34468_);
  or (_34474_, _32246_, _30016_);
  nand (_34475_, _32246_, _30016_);
  and (_34476_, _34475_, _34474_);
  and (_34477_, _34476_, _27507_);
  nor (_34478_, _31966_, _24416_);
  and (_34479_, _31966_, _24416_);
  or (_34480_, _34479_, _34478_);
  nor (_34481_, _32139_, _24668_);
  and (_34482_, _32139_, _24668_);
  or (_34483_, _34482_, _34481_);
  and (_34484_, _34483_, _34480_);
  and (_34485_, _34484_, _34477_);
  and (_34486_, _34485_, _34473_);
  nor (_34487_, _23812_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_34488_, _34487_, _34486_);
  not (_34489_, _34488_);
  nor (_34490_, _30675_, _33911_);
  and (_34491_, _30317_, _27518_);
  and (_34492_, _34491_, _34490_);
  and (_34493_, _34492_, _34473_);
  nor (_34494_, _30613_, _30446_);
  and (_34495_, _30574_, _30491_);
  and (_34496_, _34495_, _34494_);
  and (_34497_, _34496_, _30580_);
  nor (_34498_, _34497_, _33885_);
  and (_34499_, _29570_, _25437_);
  and (_34500_, _34499_, _30051_);
  nor (_34501_, _30117_, _28278_);
  and (_34502_, _34501_, _30192_);
  and (_34503_, _34502_, _34500_);
  and (_34504_, _34503_, _30268_);
  nor (_34505_, _34490_, _30693_);
  and (_34506_, _34505_, _34504_);
  and (_34507_, _34506_, _26053_);
  and (_34508_, _34490_, _25800_);
  or (_34509_, _34490_, _30374_);
  and (_34510_, _34509_, _30693_);
  and (_34511_, _34510_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_34512_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_34513_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_34514_, _34513_, _34512_);
  nor (_34515_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_34516_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_34517_, _34516_, _34515_);
  and (_34518_, _34517_, _34514_);
  and (_34519_, _34518_, _30605_);
  or (_34520_, _34519_, _34511_);
  or (_34521_, _34520_, _34508_);
  nor (_34522_, _34521_, _34507_);
  not (_34523_, _33959_);
  nor (_34524_, _34164_, _30617_);
  and (_34525_, _34524_, _34523_);
  and (_34526_, _34525_, _34122_);
  or (_34527_, _30580_, _30672_);
  nor (_34528_, _34527_, _30568_);
  or (_34529_, _34528_, _30671_);
  nand (_34530_, _34529_, _34526_);
  nand (_34531_, _34530_, _34522_);
  nand (_34532_, _30692_, _30513_);
  and (_34533_, _34532_, _30699_);
  or (_34534_, _34533_, _34522_);
  and (_34535_, _34534_, _34531_);
  and (_34536_, _34535_, _34498_);
  or (_34537_, _34536_, _30694_);
  nor (_34538_, _33949_, _30331_);
  nor (_34539_, _34538_, _30606_);
  and (_34540_, _34539_, _34537_);
  nor (_34541_, _31329_, _31313_);
  nand (_34542_, _34541_, _31323_);
  and (_34543_, _34542_, _30605_);
  or (_34544_, _31217_, _31211_);
  or (_34545_, _34544_, _31204_);
  and (_34546_, _34545_, _34510_);
  or (_34547_, _34546_, _34543_);
  nor (_34548_, _34547_, _34540_);
  not (_34549_, _34548_);
  nor (_34550_, _34549_, _34493_);
  and (_34551_, _34550_, _34489_);
  nor (_34552_, _30607_, rst);
  and (_35800_, _34552_, _34551_);
  and (_35801_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _35583_);
  and (_35802_[7], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _35583_);
  and (_34553_, _31969_, _31980_);
  and (_34554_, _34122_, _34553_);
  nand (_34555_, _34554_, _34524_);
  and (_34556_, _34555_, _30603_);
  not (_34557_, _34556_);
  not (_34558_, _30607_);
  and (_34559_, _33948_, _33951_);
  and (_34560_, _30669_, _33951_);
  nor (_34561_, _34560_, _34559_);
  and (_34562_, _34561_, _34558_);
  and (_34563_, _34562_, _34557_);
  and (_34564_, _34563_, _32030_);
  nor (_34565_, _34563_, _34326_);
  nor (_34566_, _34565_, _34564_);
  and (_34567_, _34566_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_34568_, _34566_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_34569_, _34563_, _32352_);
  nor (_34570_, _34563_, _34445_);
  nor (_34571_, _34570_, _34569_);
  and (_34572_, _34571_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_34573_, _34571_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_34574_, _34573_, _34572_);
  and (_34575_, _34563_, _32186_);
  nor (_34576_, _34563_, _34428_);
  nor (_34577_, _34576_, _34575_);
  and (_34578_, _34577_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_34579_, _34577_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_34580_, _34563_, _32290_);
  nor (_34581_, _34563_, _34411_);
  nor (_34582_, _34581_, _34580_);
  nand (_34583_, _34582_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_34584_, _34563_, _32081_);
  nor (_34585_, _34563_, _34394_);
  nor (_34586_, _34585_, _34584_);
  and (_34587_, _34586_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_34588_, _34586_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_34589_, _34563_, _32134_);
  nor (_34590_, _34563_, _34377_);
  nor (_34591_, _34590_, _34589_);
  and (_34592_, _34591_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_34593_, _34563_, _32241_);
  nor (_34594_, _34563_, _34360_);
  nor (_34595_, _34594_, _34593_);
  and (_34596_, _34595_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_34597_, _34563_, _31961_);
  nor (_34598_, _34563_, _34343_);
  nor (_34599_, _34598_, _34597_);
  and (_34600_, _34599_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_34601_, _34595_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_34602_, _34601_, _34596_);
  and (_34603_, _34602_, _34600_);
  nor (_34604_, _34603_, _34596_);
  not (_34605_, _34604_);
  nor (_34606_, _34591_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_34607_, _34606_, _34592_);
  and (_34608_, _34607_, _34605_);
  nor (_34609_, _34608_, _34592_);
  nor (_34610_, _34609_, _34588_);
  or (_34611_, _34610_, _34587_);
  or (_34612_, _34582_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_34613_, _34612_, _34583_);
  nand (_34614_, _34613_, _34611_);
  and (_34615_, _34614_, _34583_);
  nor (_34616_, _34615_, _34579_);
  or (_34617_, _34616_, _34578_);
  and (_34618_, _34617_, _34574_);
  nor (_34619_, _34618_, _34572_);
  nor (_34620_, _34619_, _34568_);
  or (_34621_, _34620_, _34567_);
  and (_34622_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_34623_, \oc8051_top_1.oc8051_memory_interface1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_34624_, _34623_, _34622_);
  and (_34625_, _34624_, _34621_);
  and (_34626_, _34625_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_34627_, _34626_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_34628_, _34627_, _34566_);
  not (_34629_, _34566_);
  nor (_34630_, _34621_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_34631_, _34630_, _30879_);
  and (_34632_, _34631_, _30884_);
  and (_34633_, _34632_, _30869_);
  nor (_34634_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_34635_, _34634_, _34633_);
  nor (_34636_, _34635_, _34629_);
  nor (_34637_, _34636_, _34628_);
  or (_34638_, _34566_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_34639_, _34566_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_34640_, _34639_, _34638_);
  nand (_34641_, _34640_, _34637_);
  nand (_34642_, _34641_, _30901_);
  not (_34643_, _34563_);
  and (_34644_, _30603_, _30581_);
  nor (_34645_, _34644_, _34538_);
  nor (_34646_, _34645_, _34643_);
  or (_34647_, _33885_, _30581_);
  nor (_34648_, _34647_, _30692_);
  and (_34649_, _34648_, _30675_);
  nand (_34650_, _34649_, _34526_);
  and (_34651_, _34650_, _30603_);
  nor (_34652_, _34651_, _34560_);
  nor (_34653_, _34652_, _34646_);
  or (_34654_, _34641_, _30901_);
  and (_34655_, _34654_, _34653_);
  and (_34656_, _34655_, _34642_);
  nor (_34657_, _34558_, _27441_);
  not (_34658_, _34644_);
  or (_34659_, _34658_, _30950_);
  not (_34660_, _33947_);
  and (_34661_, _30676_, _30548_);
  nor (_34662_, _34661_, _34022_);
  and (_34663_, _34662_, _34660_);
  nor (_34664_, _34663_, _30331_);
  nor (_34665_, _30544_, _30446_);
  and (_34666_, _34665_, _30546_);
  and (_34667_, _34666_, _30580_);
  and (_34668_, _30603_, _34667_);
  nor (_34669_, _34668_, _34664_);
  not (_34670_, _31968_);
  and (_34671_, _34662_, _34670_);
  and (_34672_, _34671_, _31980_);
  nor (_34673_, _34672_, _30331_);
  not (_34674_, _34673_);
  nor (_34675_, _34556_, _30690_);
  and (_34676_, _34675_, _34674_);
  nor (_34677_, _31968_, _30697_);
  nor (_34678_, _34677_, _30331_);
  nor (_34679_, _34678_, _34651_);
  and (_34680_, _34679_, _34676_);
  and (_34681_, _34680_, _34669_);
  and (_34682_, _34681_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_34683_, _34622_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_34684_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_34685_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_34686_, _34685_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_34687_, _34686_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_34688_, _34687_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_34689_, _34688_, _34684_);
  and (_34690_, _34689_, _34683_);
  and (_34691_, _34690_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_34692_, _34691_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_34693_, _34692_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_34694_, _34693_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_34695_, _34694_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_34696_, _34694_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_34697_, _34696_, _34695_);
  and (_34698_, _34498_, _34525_);
  and (_34699_, _34698_, _34554_);
  nor (_34700_, _34699_, _30694_);
  nor (_34701_, _34700_, _30693_);
  and (_34702_, _30549_, _33951_);
  and (_34703_, _34702_, _30588_);
  or (_34704_, _34559_, _30690_);
  or (_34705_, _34704_, _34556_);
  nor (_34706_, _34705_, _34703_);
  and (_34707_, _34497_, _30603_);
  nor (_34708_, _34707_, _34538_);
  not (_34709_, _34708_);
  and (_34710_, _34709_, _34706_);
  and (_34711_, _34710_, _34701_);
  and (_34712_, _34711_, _34697_);
  or (_34713_, _34712_, _34682_);
  and (_34714_, _34559_, _32031_);
  nor (_34715_, _34714_, _34713_);
  and (_34716_, _34715_, _34659_);
  nand (_34717_, _34716_, _34551_);
  or (_34718_, _34717_, _34657_);
  or (_34719_, _34718_, _34656_);
  nor (_34720_, _30343_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_34721_, _34720_, _31945_);
  nor (_34722_, _34721_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_34723_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_34724_, _34723_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_34725_, _34724_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not (_34726_, _34725_);
  nor (_34727_, _34726_, _34722_);
  and (_34728_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_34729_, _34728_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_34730_, _34729_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_34731_, _34730_, _34727_);
  and (_34732_, _34731_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_34733_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_34734_, _34733_, _34732_);
  and (_34735_, _34734_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_34736_, _34735_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_34737_, _34736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_34738_, _34736_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_34739_, _34738_, _34737_);
  or (_34740_, _34739_, _34551_);
  and (_34741_, _34740_, _35583_);
  and (_35803_[15], _34741_, _34719_);
  not (_34742_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_34743_, _30335_, _34742_);
  not (_34744_, _34743_);
  not (_34745_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_34746_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_34747_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_34748_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_34749_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_34750_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_34751_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_34752_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_34753_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_34754_, _34753_, _34751_);
  and (_34755_, _34754_, _34752_);
  nor (_34756_, _34755_, _34751_);
  nor (_34757_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_34758_, _34757_, _34750_);
  not (_34759_, _34758_);
  nor (_34760_, _34759_, _34756_);
  nor (_34761_, _34760_, _34750_);
  not (_34762_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_34763_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_34764_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_34765_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_34766_, _34765_, _34764_);
  and (_34767_, _34766_, _34763_);
  and (_34768_, _34767_, _34762_);
  nor (_34769_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_34770_, _34769_, _34768_);
  and (_34771_, _34770_, _34761_);
  and (_34772_, _34771_, _34749_);
  and (_34773_, _34772_, _34748_);
  and (_34774_, _34773_, _34747_);
  and (_34775_, _34774_, _34746_);
  and (_34776_, _34775_, _34745_);
  nor (_34777_, _34775_, _34745_);
  nor (_34778_, _34777_, _34776_);
  not (_34779_, _34778_);
  nor (_34780_, _34774_, _34746_);
  nor (_34781_, _34780_, _34775_);
  not (_34782_, _34781_);
  nor (_34783_, _34773_, _34747_);
  nor (_34784_, _34783_, _34774_);
  not (_34785_, _34784_);
  nor (_34786_, _34772_, _34748_);
  nor (_34787_, _34786_, _34773_);
  not (_34788_, _34787_);
  nor (_34789_, _34771_, _34749_);
  or (_34790_, _34789_, _34772_);
  not (_34791_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_34792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_34793_, _34768_, _34761_);
  and (_34794_, _34793_, _34792_);
  nor (_34795_, _34794_, _34791_);
  nor (_34796_, _34795_, _34771_);
  not (_34797_, _34796_);
  and (_34798_, _34766_, _34761_);
  and (_34799_, _34798_, _34763_);
  nor (_34800_, _34799_, _34762_);
  nor (_34801_, _34800_, _34793_);
  not (_34802_, _34801_);
  nor (_34803_, _34798_, _34763_);
  or (_34804_, _34803_, _34799_);
  and (_34805_, _34765_, _34761_);
  nor (_34806_, _34805_, _34764_);
  nor (_34807_, _34806_, _34798_);
  not (_34808_, _34807_);
  not (_34809_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_34810_, _34761_, _34809_);
  nor (_34811_, _34761_, _34809_);
  nor (_34812_, _34811_, _34810_);
  not (_34813_, _34812_);
  not (_34814_, _33858_);
  and (_34815_, _33856_, _33787_);
  and (_34816_, _33806_, _33830_);
  nor (_34817_, _34816_, _34815_);
  nor (_34818_, _34817_, _34814_);
  not (_34819_, _34818_);
  not (_34820_, _33842_);
  nor (_34821_, _34816_, _33810_);
  nor (_34822_, _34821_, _34820_);
  nor (_34823_, _33831_, _33813_);
  nor (_34824_, _34823_, _34814_);
  nor (_34825_, _34824_, _34822_);
  and (_34826_, _34825_, _34819_);
  nor (_34827_, _33854_, _33865_);
  nor (_34828_, _34827_, _34814_);
  not (_34829_, _33799_);
  and (_34830_, _33805_, _33787_);
  nor (_34831_, _33816_, _34830_);
  nor (_34832_, _34831_, _34829_);
  nor (_34833_, _34832_, _34828_);
  and (_34834_, _33834_, _33792_);
  nor (_34835_, _33857_, _33854_);
  nor (_34836_, _34835_, _34820_);
  nor (_34837_, _34836_, _34834_);
  and (_34838_, _34837_, _34833_);
  and (_34839_, _34838_, _34826_);
  and (_34840_, _34839_, _33841_);
  and (_34841_, _33800_, _33787_);
  nor (_34842_, _34841_, _33801_);
  not (_34843_, _34830_);
  and (_34844_, _34827_, _34843_);
  nor (_34845_, _34844_, _30487_);
  and (_34846_, _33842_, _33787_);
  and (_34847_, _34846_, _33830_);
  nor (_34848_, _34847_, _34845_);
  and (_34849_, _34848_, _34842_);
  nor (_34850_, _33833_, _33807_);
  nor (_34851_, _34850_, _34814_);
  nor (_34852_, _34851_, _33844_);
  and (_34853_, _33831_, _33822_);
  nor (_34854_, _34815_, _33854_);
  not (_34855_, _34854_);
  and (_34856_, _34855_, _33792_);
  nor (_34857_, _34856_, _34853_);
  and (_34858_, _34857_, _34852_);
  and (_34859_, _33796_, _33824_);
  and (_34860_, _33849_, _34859_);
  not (_34861_, _34860_);
  nor (_34862_, _30509_, _30442_);
  and (_34863_, _34862_, _33790_);
  and (_34864_, _34863_, _33787_);
  nor (_34865_, _34864_, _33817_);
  and (_34866_, _34865_, _34861_);
  nor (_34867_, _33866_, _33851_);
  and (_34868_, _34867_, _34866_);
  and (_34869_, _34868_, _34858_);
  and (_34870_, _34869_, _34849_);
  and (_34871_, _33858_, _33810_);
  and (_34872_, _33856_, _33796_);
  and (_34873_, _33822_, _34872_);
  nor (_34874_, _34873_, _34871_);
  nor (_34875_, _33864_, _33859_);
  nand (_34876_, _33811_, _30540_);
  and (_34877_, _34876_, _34875_);
  and (_34878_, _34877_, _34874_);
  not (_34879_, _34872_);
  nor (_34880_, _33842_, _33791_);
  nor (_34881_, _34880_, _34879_);
  nor (_34882_, _33804_, _33791_);
  and (_34883_, _33831_, _30540_);
  nor (_34884_, _34883_, _33837_);
  nor (_34885_, _34884_, _34882_);
  nor (_34886_, _34885_, _34881_);
  and (_34887_, _33845_, _33793_);
  and (_34888_, _34846_, _33862_);
  nor (_34889_, _34888_, _34887_);
  and (_34890_, _34889_, _34886_);
  and (_34891_, _34890_, _34878_);
  and (_34892_, _34891_, _34870_);
  and (_34893_, _34892_, _34840_);
  not (_34894_, _34893_);
  nor (_34895_, _34754_, _34752_);
  nor (_34896_, _34895_, _34755_);
  nand (_34897_, _34896_, _34894_);
  nand (_34898_, _34841_, _30370_);
  nor (_34899_, _33851_, _33844_);
  nor (_34900_, _34853_, _33835_);
  and (_34901_, _33837_, _33822_);
  nor (_34902_, _34901_, _34828_);
  and (_34903_, _34902_, _34900_);
  and (_34904_, _34903_, _34899_);
  and (_34905_, _34904_, _34898_);
  nand (_34906_, _34905_, _34878_);
  nor (_34907_, _34906_, _34893_);
  not (_34908_, _34907_);
  nor (_34909_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_34910_, _34909_, _34752_);
  and (_34911_, _34910_, _34908_);
  or (_34912_, _34896_, _34894_);
  and (_34913_, _34912_, _34897_);
  nand (_34914_, _34913_, _34911_);
  and (_34915_, _34914_, _34897_);
  not (_34916_, _34915_);
  and (_34917_, _34759_, _34756_);
  nor (_34918_, _34917_, _34760_);
  and (_34919_, _34918_, _34916_);
  and (_34920_, _34919_, _34813_);
  not (_34921_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_34922_, _34810_, _34921_);
  or (_34923_, _34922_, _34805_);
  and (_34924_, _34923_, _34920_);
  and (_34925_, _34924_, _34808_);
  and (_34926_, _34925_, _34804_);
  and (_34927_, _34926_, _34802_);
  nor (_34928_, _34793_, _34792_);
  or (_34929_, _34928_, _34794_);
  and (_34930_, _34929_, _34927_);
  and (_34931_, _34930_, _34797_);
  and (_34932_, _34931_, _34790_);
  and (_34933_, _34932_, _34788_);
  and (_34934_, _34933_, _34785_);
  and (_34935_, _34934_, _34782_);
  and (_34936_, _34935_, _34779_);
  nor (_34937_, _34936_, _34744_);
  nor (_34938_, _34743_, _30901_);
  not (_34939_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_34940_, _34776_, _34939_);
  nor (_34941_, _34776_, _34939_);
  nor (_34942_, _34941_, _34940_);
  and (_34943_, _34942_, _34743_);
  or (_34944_, _34943_, _34938_);
  or (_34945_, _34944_, _34937_);
  nand (_34946_, _34942_, _34937_);
  nor (_34947_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and (_34948_, _34947_, _34946_);
  and (_34949_, _34948_, _34945_);
  and (_34950_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _35583_);
  and (_34951_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_35804_[15], _34951_, _34949_);
  nor (_34952_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_35805_, _34952_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_35806_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _35583_);
  and (_34953_, \oc8051_top_1.oc8051_rom1.ea_int , _30332_);
  nand (_34954_, _34953_, _30335_);
  and (_35807_, _34954_, _35806_);
  and (_35808_[7], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _35583_);
  nor (_34955_, _34722_, _31945_);
  or (_34956_, _34893_, _30354_);
  nor (_34957_, _34907_, _30346_);
  nand (_34958_, _34893_, _30354_);
  and (_34959_, _34958_, _34956_);
  nand (_34960_, _34959_, _34957_);
  and (_34961_, _34960_, _34956_);
  nor (_34962_, _34961_, _31945_);
  and (_34963_, _34962_, _30342_);
  nor (_34964_, _34962_, _30342_);
  nor (_34965_, _34964_, _34963_);
  nor (_34966_, _34965_, _34955_);
  and (_34967_, _30355_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_34968_, _34967_, _34955_);
  and (_34969_, _34968_, _34906_);
  or (_34970_, _34969_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_34971_, _34970_, _34966_);
  and (_35809_[2], _34971_, _35583_);
  not (_34972_, _30483_);
  and (_34973_, _30366_, _34972_);
  nor (_34974_, _30412_, _30390_);
  and (_34975_, _34974_, _34973_);
  and (_34976_, _30336_, _35583_);
  and (_34977_, _34976_, _30459_);
  and (_34978_, _34977_, _30503_);
  nor (_34979_, _30536_, _30438_);
  and (_34980_, _34979_, _34978_);
  and (_35812_, _34980_, _34975_);
  nor (_34981_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and (_34982_, _34981_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and (_34983_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and (_35814_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _35583_);
  and (_34984_, _35814_, _34983_);
  or (_35813_[7], _34984_, _34982_);
  not (_34985_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_34986_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_34987_, _34986_, _34985_);
  and (_34988_, _34986_, _34985_);
  nor (_34989_, _34988_, _34987_);
  not (_34990_, _34989_);
  and (_34991_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_34992_, _34991_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_34993_, _34991_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_34994_, _34993_, _34992_);
  or (_34995_, _34994_, _34986_);
  and (_34996_, _34995_, _34990_);
  nor (_34997_, _34987_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_34998_, _34987_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_34999_, _34998_, _34997_);
  or (_35000_, _34992_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_35816_[3], _35000_, _35583_);
  and (_35001_, _35816_[3], _34999_);
  and (_35815_, _35001_, _34996_);
  not (_35002_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor (_35003_, _34722_, _35002_);
  and (_35004_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not (_35005_, _35003_);
  and (_35006_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_35007_, _35006_, _35004_);
  and (_35817_[31], _35007_, _35583_);
  and (_35008_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_35009_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_35010_, _35009_, _35008_);
  and (_35818_[31], _35010_, _35583_);
  and (_35011_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not (_35012_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_35013_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _35012_);
  and (_35014_, _35013_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_35015_, _35014_, _35011_);
  and (_35819_[7], _35015_, _35583_);
  and (_35016_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_35017_, _35016_, _35013_);
  and (_35820_, _35017_, _35583_);
  or (_35018_, _35012_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and (_35821_, _35018_, _35583_);
  not (_35019_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_35020_, _35019_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_35021_, _35020_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_35022_, _35012_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and (_35023_, _35022_, _35583_);
  and (_35822_[15], _35023_, _35021_);
  or (_35024_, _35012_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and (_35823_, _35024_, _35583_);
  nor (_35025_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and (_35026_, _35025_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_35027_, _35026_, _35583_);
  and (_35028_, _35814_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_35824_, _35028_, _35027_);
  and (_35029_, _35002_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_35030_, _35029_, _35026_);
  and (_35825_, _35030_, _35583_);
  nand (_35031_, _35026_, _30950_);
  or (_35032_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and (_35033_, _35032_, _35583_);
  and (_35826_[15], _35033_, _35031_);
  and (_35827_, _30723_, _31866_);
  or (_35034_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_35035_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_35036_, _34446_, _35035_);
  and (_35037_, _35036_, _35583_);
  and (_35793_[0], _35037_, _35034_);
  or (_35038_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_35039_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_35040_, _34446_, _35039_);
  and (_35041_, _35040_, _35583_);
  and (_35793_[1], _35041_, _35038_);
  or (_35042_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_35043_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_35044_, _34446_, _35043_);
  and (_35045_, _35044_, _35583_);
  and (_35793_[2], _35045_, _35042_);
  or (_35046_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_35047_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_35048_, _34446_, _35047_);
  and (_35049_, _35048_, _35583_);
  and (_35793_[3], _35049_, _35046_);
  or (_35050_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not (_35051_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_35052_, _34446_, _35051_);
  and (_35053_, _35052_, _35583_);
  and (_35793_[4], _35053_, _35050_);
  or (_35054_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_35055_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_35056_, _34446_, _35055_);
  and (_35057_, _35056_, _35583_);
  and (_35793_[5], _35057_, _35054_);
  or (_35058_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_35059_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_35060_, _34446_, _35059_);
  and (_35061_, _35060_, _35583_);
  and (_35793_[6], _35061_, _35058_);
  or (_35062_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not (_35063_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_35064_, _34446_, _35063_);
  and (_35065_, _35064_, _35583_);
  and (_35793_[7], _35065_, _35062_);
  or (_35066_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_35067_, _34446_, _30873_);
  and (_35068_, _35067_, _35583_);
  and (_35793_[8], _35068_, _35066_);
  or (_35069_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_35070_, _34446_, _30879_);
  and (_35071_, _35070_, _35583_);
  and (_35793_[9], _35071_, _35069_);
  or (_35072_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_35073_, _34446_, _30884_);
  and (_35074_, _35073_, _35583_);
  and (_35793_[10], _35074_, _35072_);
  or (_35075_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_35076_, _34446_, _30869_);
  and (_35077_, _35076_, _35583_);
  and (_35793_[11], _35077_, _35075_);
  or (_35078_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_35079_, _34446_, _30890_);
  and (_35080_, _35079_, _35583_);
  and (_35793_[12], _35080_, _35078_);
  or (_35081_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_35082_, _34446_, _30865_);
  and (_35083_, _35082_, _35583_);
  and (_35793_[13], _35083_, _35081_);
  or (_35084_, _34446_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_35085_, _34446_, _30896_);
  and (_35086_, _35085_, _35583_);
  and (_35793_[14], _35086_, _35084_);
  or (_35087_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_35088_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _35583_);
  or (_35089_, _35088_, _00000_);
  and (_35794_[0], _35089_, _35087_);
  or (_35090_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_35091_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _35583_);
  or (_35092_, _35091_, _00000_);
  and (_35794_[1], _35092_, _35090_);
  or (_35093_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_35094_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _35583_);
  or (_35095_, _35094_, _00000_);
  and (_35794_[2], _35095_, _35093_);
  or (_35096_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_35097_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _35583_);
  or (_35098_, _35097_, _00000_);
  and (_35794_[3], _35098_, _35096_);
  or (_35099_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_35100_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _35583_);
  or (_35101_, _35100_, _00000_);
  and (_35794_[4], _35101_, _35099_);
  or (_35102_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_35103_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _35583_);
  or (_35104_, _35103_, _00000_);
  and (_35794_[5], _35104_, _35102_);
  or (_35105_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and (_35106_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _35583_);
  or (_35107_, _35106_, _00000_);
  and (_35794_[6], _35107_, _35105_);
  or (_35108_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_35109_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _35583_);
  or (_35110_, _35109_, _00000_);
  and (_35794_[7], _35110_, _35108_);
  or (_35111_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_35112_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _35583_);
  or (_35113_, _35112_, _00000_);
  and (_35794_[8], _35113_, _35111_);
  or (_35114_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_35115_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _35583_);
  or (_35116_, _35115_, _00000_);
  and (_35794_[9], _35116_, _35114_);
  or (_35117_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_35118_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _35583_);
  or (_35119_, _35118_, _00000_);
  and (_35794_[10], _35119_, _35117_);
  or (_35120_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_35121_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _35583_);
  or (_35122_, _35121_, _00000_);
  and (_35794_[11], _35122_, _35120_);
  or (_35123_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_35124_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _35583_);
  or (_35125_, _35124_, _00000_);
  and (_35794_[12], _35125_, _35123_);
  or (_35126_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_35127_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _35583_);
  or (_35128_, _35127_, _00000_);
  and (_35794_[13], _35128_, _35126_);
  or (_35129_, _34450_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_35130_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _35583_);
  or (_35131_, _35130_, _00000_);
  and (_35794_[14], _35131_, _35129_);
  and (_35132_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_35133_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or (_35134_, _35133_, _35132_);
  and (_35817_[0], _35134_, _35583_);
  and (_35135_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_35136_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_35137_, _35136_, _35135_);
  and (_35817_[1], _35137_, _35583_);
  and (_35138_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_35139_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_35140_, _35139_, _35138_);
  and (_35817_[2], _35140_, _35583_);
  and (_35141_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_35142_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or (_35143_, _35142_, _35141_);
  and (_35817_[3], _35143_, _35583_);
  and (_35144_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_35145_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or (_35146_, _35145_, _35144_);
  and (_35817_[4], _35146_, _35583_);
  and (_35147_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_35148_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_35149_, _35148_, _35147_);
  and (_35817_[5], _35149_, _35583_);
  and (_35150_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_35151_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_35152_, _35151_, _35150_);
  and (_35817_[6], _35152_, _35583_);
  and (_35153_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_35154_, _35003_, _34983_);
  or (_35155_, _35154_, _35153_);
  and (_35817_[7], _35155_, _35583_);
  and (_35156_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and (_35157_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or (_35158_, _35157_, _35156_);
  and (_35817_[8], _35158_, _35583_);
  and (_35159_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and (_35160_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_35161_, _35160_, _35159_);
  and (_35817_[9], _35161_, _35583_);
  and (_35162_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and (_35163_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_35164_, _35163_, _35162_);
  and (_35817_[10], _35164_, _35583_);
  and (_35165_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and (_35166_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_35167_, _35166_, _35165_);
  and (_35817_[11], _35167_, _35583_);
  and (_35168_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and (_35169_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_35170_, _35169_, _35168_);
  and (_35817_[12], _35170_, _35583_);
  and (_35171_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and (_35172_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_35173_, _35172_, _35171_);
  and (_35817_[13], _35173_, _35583_);
  and (_35174_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and (_35175_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_35176_, _35175_, _35174_);
  and (_35817_[14], _35176_, _35583_);
  and (_35177_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and (_35178_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_35179_, _35178_, _35177_);
  and (_35817_[15], _35179_, _35583_);
  and (_35180_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and (_35181_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_35182_, _35181_, _35180_);
  and (_35817_[16], _35182_, _35583_);
  and (_35183_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and (_35184_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_35185_, _35184_, _35183_);
  and (_35817_[17], _35185_, _35583_);
  and (_35186_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and (_35187_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or (_35188_, _35187_, _35186_);
  and (_35817_[18], _35188_, _35583_);
  and (_35189_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and (_35190_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or (_35191_, _35190_, _35189_);
  and (_35817_[19], _35191_, _35583_);
  and (_35192_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and (_35193_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_35194_, _35193_, _35192_);
  and (_35817_[20], _35194_, _35583_);
  and (_35195_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and (_35196_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_35197_, _35196_, _35195_);
  and (_35817_[21], _35197_, _35583_);
  and (_35198_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and (_35199_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_35200_, _35199_, _35198_);
  and (_35817_[22], _35200_, _35583_);
  and (_35201_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and (_35202_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or (_35203_, _35202_, _35201_);
  and (_35817_[23], _35203_, _35583_);
  and (_35204_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and (_35205_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_35206_, _35205_, _35204_);
  and (_35817_[24], _35206_, _35583_);
  and (_35207_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and (_35208_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_35209_, _35208_, _35207_);
  and (_35817_[25], _35209_, _35583_);
  and (_35210_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and (_35211_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_35212_, _35211_, _35210_);
  and (_35817_[26], _35212_, _35583_);
  and (_35213_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and (_35214_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_35215_, _35214_, _35213_);
  and (_35817_[27], _35215_, _35583_);
  and (_35216_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and (_35217_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_35218_, _35217_, _35216_);
  and (_35817_[28], _35218_, _35583_);
  and (_35219_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and (_35220_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or (_35221_, _35220_, _35219_);
  and (_35817_[29], _35221_, _35583_);
  and (_35222_, _35003_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and (_35223_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_35224_, _35223_, _35222_);
  and (_35817_[30], _35224_, _35583_);
  nor (_35796_[0], _30544_, rst);
  nor (_35796_[1], _30446_, rst);
  nor (_35796_[2], _30468_, rst);
  nor (_35796_[3], _31878_, rst);
  and (_35797_[0], _31933_, _35583_);
  and (_35797_[1], _32226_, _35583_);
  and (_35797_[2], _32114_, _35583_);
  and (_35797_[3], _32060_, _35583_);
  nor (_35797_[4], _32271_, rst);
  nor (_35797_[5], _32164_, rst);
  nor (_35797_[6], _32335_, rst);
  and (_35802_[0], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _35583_);
  and (_35802_[1], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _35583_);
  and (_35802_[2], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _35583_);
  and (_35802_[3], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _35583_);
  and (_35802_[4], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _35583_);
  and (_35802_[5], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _35583_);
  and (_35802_[6], \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _35583_);
  or (_35225_, _34551_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_35226_, _35225_, _35583_);
  not (_35227_, _34651_);
  and (_35228_, _34645_, _34563_);
  and (_35229_, _35228_, _35227_);
  or (_35230_, _35229_, _34644_);
  and (_35231_, _35230_, _28567_);
  or (_35232_, _34599_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_35233_, _34600_);
  and (_35234_, _34653_, _35233_);
  and (_35235_, _35234_, _35232_);
  and (_35236_, _34559_, _34343_);
  and (_35237_, _30607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_35238_, _35227_, _34646_);
  and (_35239_, _35238_, _31962_);
  or (_35240_, _35239_, _35237_);
  or (_35241_, _35240_, _35236_);
  nor (_35242_, _35241_, _35235_);
  nand (_35243_, _35242_, _34551_);
  or (_35244_, _35243_, _35231_);
  and (_35803_[0], _35244_, _35226_);
  or (_35245_, _34551_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_35246_, _35245_, _35583_);
  and (_35247_, _35230_, _29253_);
  or (_35248_, _34602_, _34600_);
  not (_35249_, _34603_);
  and (_35250_, _34653_, _35249_);
  and (_35251_, _35250_, _35248_);
  and (_35252_, _34559_, _34360_);
  and (_35253_, _35238_, _32242_);
  and (_35254_, _30607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_35255_, _35254_, _35253_);
  or (_35256_, _35255_, _35252_);
  nor (_35257_, _35256_, _35251_);
  nand (_35258_, _35257_, _34551_);
  or (_35259_, _35258_, _35247_);
  and (_35803_[1], _35259_, _35246_);
  not (_35260_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_35261_, _34722_, _35260_);
  and (_35262_, _34722_, _35260_);
  nor (_35263_, _35262_, _35261_);
  or (_35264_, _35263_, _34551_);
  and (_35265_, _35264_, _35583_);
  and (_35266_, _35230_, _29898_);
  or (_35267_, _34607_, _34605_);
  not (_35268_, _34608_);
  and (_35269_, _34653_, _35268_);
  and (_35270_, _35269_, _35267_);
  and (_35271_, _34559_, _34377_);
  and (_35272_, _35238_, _32135_);
  and (_35273_, _30607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_35274_, _35273_, _35272_);
  or (_35275_, _35274_, _35271_);
  nor (_35276_, _35275_, _35270_);
  nand (_35277_, _35276_, _34551_);
  or (_35278_, _35277_, _35266_);
  and (_35803_[2], _35278_, _35265_);
  and (_35279_, _35261_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_35280_, _35261_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_35281_, _35280_, _35279_);
  or (_35282_, _35281_, _34551_);
  and (_35283_, _35282_, _35583_);
  and (_35284_, _35230_, _30093_);
  or (_35285_, _34588_, _34587_);
  or (_35286_, _35285_, _34609_);
  nand (_35287_, _35285_, _34609_);
  and (_35288_, _35287_, _34653_);
  and (_35289_, _35288_, _35286_);
  and (_35290_, _34559_, _34394_);
  and (_35291_, _35238_, _32082_);
  and (_35292_, _30607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_35293_, _35292_, _35291_);
  or (_35294_, _35293_, _35290_);
  nor (_35295_, _35294_, _35289_);
  nand (_35296_, _35295_, _34551_);
  or (_35297_, _35296_, _35284_);
  and (_35803_[3], _35297_, _35283_);
  not (_35298_, _34722_);
  and (_35299_, _34724_, _35298_);
  nor (_35300_, _35279_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_35301_, _35300_, _35299_);
  or (_35302_, _35301_, _34551_);
  and (_35303_, _35302_, _35583_);
  and (_35304_, _35230_, _30162_);
  or (_35305_, _34613_, _34611_);
  and (_35306_, _34653_, _34614_);
  and (_35307_, _35306_, _35305_);
  and (_35308_, _34559_, _34411_);
  and (_35309_, _35238_, _32291_);
  and (_35310_, _30607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_35311_, _35310_, _35309_);
  or (_35312_, _35311_, _35308_);
  nor (_35313_, _35312_, _35307_);
  nand (_35314_, _35313_, _34551_);
  or (_35315_, _35314_, _35304_);
  and (_35803_[4], _35315_, _35303_);
  nor (_35316_, _35299_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_35317_, _35316_, _34727_);
  or (_35318_, _35317_, _34551_);
  and (_35319_, _35318_, _35583_);
  and (_35320_, _35230_, _30237_);
  or (_35321_, _34579_, _34578_);
  or (_35322_, _35321_, _34615_);
  nand (_35323_, _35321_, _34615_);
  and (_35324_, _35323_, _34653_);
  and (_35325_, _35324_, _35322_);
  and (_35326_, _35238_, _32187_);
  and (_35327_, _34559_, _34428_);
  and (_35328_, _30607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_35329_, _35328_, _35327_);
  or (_35330_, _35329_, _35326_);
  nor (_35331_, _35330_, _35325_);
  nand (_35332_, _35331_, _34551_);
  or (_35333_, _35332_, _35320_);
  and (_35803_[5], _35333_, _35319_);
  nor (_35334_, _34727_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_35335_, _34727_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_35336_, _35335_, _35334_);
  or (_35337_, _35336_, _34551_);
  and (_35338_, _35337_, _35583_);
  and (_35339_, _35230_, _30310_);
  or (_35340_, _34617_, _34574_);
  not (_35341_, _34618_);
  and (_35342_, _34653_, _35341_);
  nand (_35343_, _35342_, _35340_);
  nand (_35344_, _34559_, _34445_);
  nand (_35345_, _35238_, _32353_);
  nand (_35346_, _30607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_35347_, _35346_, _35345_);
  and (_35348_, _35347_, _35344_);
  and (_35349_, _35348_, _35343_);
  nand (_35350_, _35349_, _34551_);
  or (_35351_, _35350_, _35339_);
  and (_35803_[6], _35351_, _35338_);
  nor (_35352_, _35335_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_35353_, _35335_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_35354_, _35353_, _35352_);
  or (_35355_, _35354_, _34551_);
  and (_35356_, _35355_, _35583_);
  and (_35357_, _35230_, _27452_);
  or (_35358_, _34567_, _34568_);
  or (_35359_, _35358_, _34619_);
  nand (_35360_, _35358_, _34619_);
  and (_35361_, _35360_, _34653_);
  and (_35362_, _35361_, _35359_);
  nand (_35363_, _34559_, _34326_);
  nand (_35364_, _35238_, _32031_);
  nand (_35365_, _30607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_35366_, _35365_, _35364_);
  and (_35367_, _35366_, _35363_);
  nand (_35368_, _35367_, _34551_);
  or (_35369_, _35368_, _35362_);
  or (_35370_, _35369_, _35357_);
  and (_35803_[7], _35370_, _35356_);
  or (_35371_, _35353_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand (_35372_, _34729_, _34727_);
  and (_35373_, _35372_, _35371_);
  or (_35374_, _35373_, _34551_);
  and (_35375_, _35374_, _35583_);
  nor (_35376_, _34558_, _28556_);
  nor (_35377_, _34658_, _30988_);
  and (_35378_, _34621_, _30873_);
  nor (_35379_, _34621_, _30873_);
  nor (_35380_, _35379_, _35378_);
  nand (_35381_, _35380_, _34629_);
  or (_35382_, _35380_, _34629_);
  and (_35383_, _35382_, _34653_);
  and (_35384_, _35383_, _35381_);
  nand (_35385_, _35238_, _33824_);
  and (_35386_, _34681_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_35387_, _34559_, _31962_);
  nor (_35388_, _35387_, _35386_);
  and (_35389_, _35388_, _35385_);
  nand (_35390_, _35389_, _34551_);
  or (_35391_, _35390_, _35384_);
  or (_35392_, _35391_, _35377_);
  or (_35393_, _35392_, _35376_);
  and (_35803_[8], _35393_, _35375_);
  nand (_35394_, _35372_, _34791_);
  or (_35395_, _35372_, _34791_);
  and (_35396_, _35395_, _35394_);
  or (_35397_, _35396_, _34551_);
  and (_35398_, _35397_, _35583_);
  nor (_35399_, _30691_, _29242_);
  and (_35400_, _34486_, _28082_);
  and (_35401_, _35400_, _27474_);
  not (_35402_, _35401_);
  and (_35403_, _30588_, _30579_);
  and (_35404_, _35403_, _30603_);
  and (_35405_, _34542_, _35404_);
  or (_35406_, _35405_, _34540_);
  and (_35407_, _30693_, _30374_);
  and (_35408_, _34545_, _35407_);
  nor (_35409_, _34553_, _33911_);
  and (_35410_, _35409_, _30317_);
  and (_35411_, _35410_, _27518_);
  and (_35412_, _35411_, _34473_);
  or (_35413_, _35412_, _35408_);
  nor (_35414_, _35413_, _35406_);
  and (_35415_, _35414_, _35402_);
  nor (_35416_, _34658_, _31019_);
  and (_35417_, _34681_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_35418_, _35238_, _33795_);
  and (_35419_, _34559_, _32242_);
  or (_35420_, _35419_, _35418_);
  or (_35421_, _35420_, _35417_);
  or (_35422_, _35421_, _35416_);
  not (_35423_, _34701_);
  nor (_35424_, _35423_, _34703_);
  nor (_35425_, _35424_, _34710_);
  and (_35426_, _34621_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_35427_, _35426_, _34629_);
  and (_35428_, _34630_, _34566_);
  nor (_35429_, _35428_, _35427_);
  and (_35430_, _35429_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_35431_, _35429_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_35432_, _35431_, _35430_);
  and (_35433_, _35432_, _35425_);
  nor (_35434_, _35433_, _35422_);
  nand (_35435_, _35434_, _35415_);
  or (_35436_, _35435_, _35399_);
  and (_35803_[9], _35436_, _35398_);
  nor (_35437_, _34731_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_35438_, _35437_, _34732_);
  or (_35439_, _35438_, _34551_);
  and (_35440_, _35439_, _35583_);
  not (_35441_, _35415_);
  and (_35442_, _34631_, _34566_);
  and (_35443_, _35427_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_35444_, _35443_, _35442_);
  nor (_35445_, _35444_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_35446_, _35444_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_35447_, _35446_, _35445_);
  and (_35448_, _35447_, _35425_);
  nor (_35449_, _34658_, _31049_);
  and (_35450_, _34681_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_35451_, _34711_, _33786_);
  or (_35452_, _35451_, _35450_);
  and (_35453_, _34559_, _32135_);
  or (_35454_, _35453_, _35452_);
  or (_35455_, _35454_, _35449_);
  nor (_35456_, _30691_, _29887_);
  or (_35457_, _35456_, _35455_);
  or (_35458_, _35457_, _35448_);
  or (_35459_, _35458_, _35441_);
  and (_35803_[10], _35459_, _35440_);
  nor (_35460_, _34732_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_35461_, _34725_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_35462_, _35461_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_35463_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_35464_, _35463_, _35462_);
  and (_35465_, _35464_, _35298_);
  and (_35466_, _35465_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_35467_, _35466_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_35468_, _35467_, _35460_);
  or (_35469_, _35468_, _34551_);
  and (_35470_, _35469_, _35583_);
  nor (_35471_, _30691_, _30092_);
  nor (_35472_, _34658_, _31078_);
  and (_35473_, _34681_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_35474_, _34559_, _32082_);
  nor (_35475_, _34690_, _30869_);
  and (_35476_, _34690_, _30869_);
  or (_35477_, _35476_, _35475_);
  and (_35478_, _35477_, _35238_);
  or (_35479_, _35478_, _35474_);
  or (_35480_, _35479_, _35473_);
  or (_35481_, _35480_, _35472_);
  and (_35482_, _34683_, _34621_);
  and (_35483_, _35482_, _34629_);
  and (_35484_, _34632_, _34566_);
  nor (_35485_, _35484_, _35483_);
  or (_35486_, _35485_, _30869_);
  nand (_35487_, _35485_, _30869_);
  and (_35488_, _35487_, _35486_);
  and (_35489_, _35488_, _35425_);
  or (_35490_, _35489_, _35481_);
  or (_35491_, _35490_, _35471_);
  or (_35492_, _35491_, _35441_);
  and (_35803_[11], _35492_, _35470_);
  nor (_35493_, _35467_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_35494_, _35493_, _34734_);
  or (_35495_, _35494_, _34551_);
  and (_35496_, _35495_, _35583_);
  nor (_35497_, _34558_, _30161_);
  and (_35498_, _34625_, _34629_);
  and (_35499_, _34566_, _30869_);
  and (_35500_, _35499_, _34632_);
  nor (_35501_, _35500_, _35498_);
  nand (_35502_, _35501_, _30890_);
  or (_35503_, _35501_, _30890_);
  and (_35504_, _35503_, _34653_);
  and (_35505_, _35504_, _35502_);
  or (_35506_, _34658_, _31110_);
  and (_35507_, _34681_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_35508_, _34691_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_35509_, _35508_, _34692_);
  and (_35510_, _35509_, _34711_);
  or (_35511_, _35510_, _35507_);
  and (_35512_, _34559_, _32291_);
  nor (_35513_, _35512_, _35511_);
  and (_35514_, _35513_, _35506_);
  nand (_35515_, _35514_, _34551_);
  or (_35516_, _35515_, _35505_);
  or (_35517_, _35516_, _35497_);
  and (_35803_[12], _35517_, _35496_);
  nor (_35518_, _34734_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_35519_, _35518_, _34735_);
  or (_35520_, _35519_, _34551_);
  and (_35521_, _35520_, _35583_);
  nor (_35522_, _34558_, _30236_);
  and (_35523_, _34626_, _34629_);
  and (_35524_, _35500_, _30890_);
  nor (_35525_, _35524_, _35523_);
  nand (_35526_, _35525_, _30865_);
  or (_35527_, _35525_, _30865_);
  and (_35528_, _35527_, _34653_);
  and (_35529_, _35528_, _35526_);
  or (_35530_, _34658_, _31143_);
  and (_35531_, _34681_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_35532_, _34689_, _34624_);
  and (_35533_, _35532_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_35534_, _35533_, _30865_);
  and (_35535_, _35533_, _30865_);
  or (_35536_, _35535_, _35534_);
  and (_35537_, _35536_, _34711_);
  or (_35538_, _35537_, _35531_);
  and (_35539_, _34559_, _32187_);
  nor (_35540_, _35539_, _35538_);
  and (_35541_, _35540_, _35530_);
  nand (_35542_, _35541_, _34551_);
  or (_35543_, _35542_, _35529_);
  or (_35544_, _35543_, _35522_);
  and (_35803_[13], _35544_, _35521_);
  or (_35545_, _34735_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_35546_, _35545_, _34736_);
  or (_35547_, _35546_, _34551_);
  and (_35548_, _35547_, _35583_);
  nand (_35549_, _34637_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_35550_, _34637_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_35551_, _35550_, _34653_);
  and (_35552_, _35551_, _35549_);
  nor (_35553_, _34558_, _30309_);
  or (_35554_, _34658_, _31175_);
  and (_35555_, _34681_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_35556_, _34693_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_35557_, _35556_, _34694_);
  and (_35558_, _35557_, _34711_);
  or (_35559_, _35558_, _35555_);
  and (_35560_, _34559_, _32353_);
  nor (_35561_, _35560_, _35559_);
  and (_35562_, _35561_, _35554_);
  nand (_35563_, _35562_, _34551_);
  or (_35564_, _35563_, _35553_);
  or (_35565_, _35564_, _35552_);
  and (_35803_[14], _35565_, _35548_);
  and (_35566_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_35567_, _34910_, _34908_);
  nor (_35568_, _35567_, _34911_);
  or (_35569_, _35568_, _34744_);
  or (_35570_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_35571_, _35570_, _34947_);
  and (_35572_, _35571_, _35569_);
  or (_35804_[0], _35572_, _35566_);
  and (_35573_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_35574_, _34913_, _34911_);
  and (_35575_, _35574_, _34914_);
  or (_35576_, _35575_, _34744_);
  or (_35577_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_35578_, _35577_, _34947_);
  and (_35579_, _35578_, _35576_);
  or (_35804_[1], _35579_, _35573_);
  or (_35580_, _34918_, _34916_);
  nor (_35581_, _34919_, _34744_);
  and (_00008_, _35581_, _35580_);
  nor (_00009_, _34743_, _35043_);
  or (_00010_, _00009_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00011_, _00010_, _00008_);
  or (_00012_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _30332_);
  and (_00013_, _00012_, _35583_);
  and (_35804_[2], _00013_, _00011_);
  nor (_00014_, _34919_, _34813_);
  nor (_00015_, _00014_, _34920_);
  or (_00016_, _00015_, _34744_);
  or (_00017_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00018_, _00017_, _34947_);
  and (_00019_, _00018_, _00016_);
  and (_00020_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_35804_[3], _00020_, _00019_);
  nor (_00021_, _34923_, _34920_);
  nor (_00022_, _00021_, _34924_);
  or (_00023_, _00022_, _34744_);
  or (_00024_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00025_, _00024_, _34947_);
  and (_00026_, _00025_, _00023_);
  and (_00027_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_35804_[4], _00027_, _00026_);
  and (_00028_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_00029_, _34924_, _34808_);
  nor (_00030_, _00029_, _34925_);
  or (_00031_, _00030_, _34744_);
  or (_00032_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_00033_, _00032_, _34947_);
  and (_00034_, _00033_, _00031_);
  or (_35804_[5], _00034_, _00028_);
  and (_00035_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00036_, _34925_, _34804_);
  nor (_00037_, _00036_, _34926_);
  or (_00038_, _00037_, _34744_);
  or (_00039_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00040_, _00039_, _34947_);
  and (_00041_, _00040_, _00038_);
  or (_35804_[6], _00041_, _00035_);
  and (_00042_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_00043_, _34926_, _34802_);
  nor (_00044_, _00043_, _34927_);
  or (_00045_, _00044_, _34744_);
  or (_00046_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_00047_, _00046_, _34947_);
  and (_00048_, _00047_, _00045_);
  or (_35804_[7], _00048_, _00042_);
  nor (_00049_, _34929_, _34927_);
  nor (_00050_, _00049_, _34930_);
  or (_00051_, _00050_, _34744_);
  or (_00052_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00053_, _00052_, _34947_);
  and (_00054_, _00053_, _00051_);
  and (_00055_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_35804_[8], _00055_, _00054_);
  nor (_00056_, _34930_, _34797_);
  nor (_00057_, _00056_, _34931_);
  or (_00058_, _00057_, _34744_);
  or (_00059_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00060_, _00059_, _34947_);
  and (_00061_, _00060_, _00058_);
  and (_00062_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_35804_[9], _00062_, _00061_);
  nor (_00063_, _34931_, _34790_);
  nor (_00064_, _00063_, _34932_);
  or (_00065_, _00064_, _34744_);
  or (_00066_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00067_, _00066_, _34947_);
  and (_00068_, _00067_, _00065_);
  and (_00069_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_35804_[10], _00069_, _00068_);
  nor (_00070_, _34932_, _34788_);
  nor (_00071_, _00070_, _34933_);
  or (_00072_, _00071_, _34744_);
  or (_00073_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00074_, _00073_, _34947_);
  and (_00075_, _00074_, _00072_);
  and (_00076_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_35804_[11], _00076_, _00075_);
  nor (_00077_, _34933_, _34785_);
  nor (_00078_, _00077_, _34934_);
  or (_00079_, _00078_, _34744_);
  or (_00080_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00081_, _00080_, _34947_);
  and (_00082_, _00081_, _00079_);
  and (_00083_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_35804_[12], _00083_, _00082_);
  nor (_00084_, _34934_, _34782_);
  nor (_00085_, _00084_, _34935_);
  or (_00086_, _00085_, _34744_);
  or (_00087_, _34743_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00088_, _00087_, _34947_);
  and (_00089_, _00088_, _00086_);
  and (_00090_, _34950_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_35804_[13], _00090_, _00089_);
  or (_00091_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _30332_);
  and (_00092_, _00091_, _35583_);
  or (_00093_, _34935_, _34779_);
  and (_00094_, _00093_, _34937_);
  nor (_00095_, _34743_, _30896_);
  or (_00096_, _00095_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00097_, _00096_, _00094_);
  and (_35804_[14], _00097_, _00092_);
  and (_35808_[0], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _35583_);
  and (_35808_[1], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _35583_);
  and (_35808_[2], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _35583_);
  and (_35808_[3], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _35583_);
  and (_35808_[4], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _35583_);
  and (_35808_[5], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _35583_);
  and (_35808_[6], \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _35583_);
  nor (_00098_, _34907_, _31945_);
  nand (_00099_, _00098_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_00100_, _00098_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_00101_, _00100_, _34947_);
  and (_35809_[0], _00101_, _00099_);
  or (_00102_, _34959_, _34957_);
  and (_00103_, _00102_, _34960_);
  or (_00104_, _00103_, _31945_);
  or (_00105_, _30335_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00106_, _00105_, _34947_);
  and (_35809_[1], _00106_, _00104_);
  and (_00107_, _34981_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and (_00108_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and (_00109_, _00108_, _35814_);
  or (_35813_[0], _00109_, _00107_);
  and (_00110_, _34981_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and (_00111_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and (_00112_, _00111_, _35814_);
  or (_35813_[1], _00112_, _00110_);
  and (_00113_, _34981_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and (_00114_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and (_00115_, _00114_, _35814_);
  or (_35813_[2], _00115_, _00113_);
  and (_00116_, _34981_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and (_00117_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and (_00118_, _00117_, _35814_);
  or (_35813_[3], _00118_, _00116_);
  and (_00119_, _34981_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and (_00120_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and (_00121_, _00120_, _35814_);
  or (_35813_[4], _00121_, _00119_);
  and (_00122_, _34981_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_00123_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and (_00124_, _00123_, _35814_);
  or (_35813_[5], _00124_, _00122_);
  and (_00125_, _34981_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and (_00126_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and (_00127_, _00126_, _35814_);
  or (_35813_[6], _00127_, _00125_);
  and (_35816_[0], _34989_, _35583_);
  nor (_35816_[1], _34999_, rst);
  and (_35816_[2], _34995_, _35583_);
  and (_00128_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_00129_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or (_00130_, _00129_, _00128_);
  and (_35818_[0], _00130_, _35583_);
  and (_00131_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_00132_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or (_00133_, _00132_, _00131_);
  and (_35818_[1], _00133_, _35583_);
  and (_00134_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_00135_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or (_00136_, _00135_, _00134_);
  and (_35818_[2], _00136_, _35583_);
  and (_00137_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_00138_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or (_00139_, _00138_, _00137_);
  and (_35818_[3], _00139_, _35583_);
  and (_00140_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_00141_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or (_00142_, _00141_, _00140_);
  and (_35818_[4], _00142_, _35583_);
  and (_00143_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_00144_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or (_00145_, _00144_, _00143_);
  and (_35818_[5], _00145_, _35583_);
  and (_00146_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_00147_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or (_00148_, _00147_, _00146_);
  and (_35818_[6], _00148_, _35583_);
  and (_00149_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_00150_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or (_00151_, _00150_, _00149_);
  and (_35818_[7], _00151_, _35583_);
  and (_00152_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_00153_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or (_00154_, _00153_, _00152_);
  and (_35818_[8], _00154_, _35583_);
  and (_00155_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_00156_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or (_00157_, _00156_, _00155_);
  and (_35818_[9], _00157_, _35583_);
  and (_00158_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_00159_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or (_00160_, _00159_, _00158_);
  and (_35818_[10], _00160_, _35583_);
  and (_00161_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_00162_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or (_00163_, _00162_, _00161_);
  and (_35818_[11], _00163_, _35583_);
  and (_00164_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_00165_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or (_00166_, _00165_, _00164_);
  and (_35818_[12], _00166_, _35583_);
  and (_00167_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_00168_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or (_00169_, _00168_, _00167_);
  and (_35818_[13], _00169_, _35583_);
  and (_00170_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_00171_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_00172_, _00171_, _00170_);
  and (_35818_[14], _00172_, _35583_);
  and (_00173_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_00174_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or (_00175_, _00174_, _00173_);
  and (_35818_[15], _00175_, _35583_);
  and (_00176_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_00177_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or (_00178_, _00177_, _00176_);
  and (_35818_[16], _00178_, _35583_);
  and (_00179_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00180_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_00181_, _00180_, _00179_);
  and (_35818_[17], _00181_, _35583_);
  and (_00182_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_00183_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_00184_, _00183_, _00182_);
  and (_35818_[18], _00184_, _35583_);
  and (_00185_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_00186_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_00187_, _00186_, _00185_);
  and (_35818_[19], _00187_, _35583_);
  and (_00188_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_00189_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_00190_, _00189_, _00188_);
  and (_35818_[20], _00190_, _35583_);
  and (_00191_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_00192_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_00193_, _00192_, _00191_);
  and (_35818_[21], _00193_, _35583_);
  and (_00194_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_00195_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_00196_, _00195_, _00194_);
  and (_35818_[22], _00196_, _35583_);
  and (_00197_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00198_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_00199_, _00198_, _00197_);
  and (_35818_[23], _00199_, _35583_);
  and (_00200_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00201_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or (_00202_, _00201_, _00200_);
  and (_35818_[24], _00202_, _35583_);
  and (_00203_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00204_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_00205_, _00204_, _00203_);
  and (_35818_[25], _00205_, _35583_);
  and (_00206_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00207_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_00208_, _00207_, _00206_);
  and (_35818_[26], _00208_, _35583_);
  and (_00209_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00210_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_00211_, _00210_, _00209_);
  and (_35818_[27], _00211_, _35583_);
  and (_00212_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_00213_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_00214_, _00213_, _00212_);
  and (_35818_[28], _00214_, _35583_);
  and (_00215_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_00216_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_00217_, _00216_, _00215_);
  and (_35818_[29], _00217_, _35583_);
  and (_00218_, _35003_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_00219_, _35005_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_00220_, _00219_, _00218_);
  and (_35818_[30], _00220_, _35583_);
  and (_00221_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00222_, _35013_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00223_, _00222_, _00221_);
  and (_35819_[0], _00223_, _35583_);
  and (_00224_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00225_, _35013_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00226_, _00225_, _00224_);
  and (_35819_[1], _00226_, _35583_);
  and (_00227_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00228_, _35013_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00229_, _00228_, _00227_);
  and (_35819_[2], _00229_, _35583_);
  and (_00230_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00231_, _35013_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00232_, _00231_, _00230_);
  and (_35819_[3], _00232_, _35583_);
  and (_00233_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00234_, _35013_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_00235_, _00234_, _00233_);
  and (_35819_[4], _00235_, _35583_);
  and (_00236_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00237_, _35013_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_00238_, _00237_, _00236_);
  and (_35819_[5], _00238_, _35583_);
  and (_00239_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_00240_, _35013_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_00241_, _00240_, _00239_);
  and (_35819_[6], _00241_, _35583_);
  and (_00242_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00243_, _31933_, _35019_);
  or (_00244_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00245_, _00244_, _35012_);
  and (_00246_, _00245_, _00243_);
  or (_00247_, _00246_, _00242_);
  and (_35822_[0], _00247_, _35583_);
  and (_00248_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00249_, _32226_, _35019_);
  or (_00250_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00251_, _00250_, _35012_);
  and (_00252_, _00251_, _00249_);
  or (_00253_, _00252_, _00248_);
  and (_35822_[1], _00253_, _35583_);
  and (_00254_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00255_, _32114_, _35019_);
  or (_00256_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00257_, _00256_, _35012_);
  and (_00258_, _00257_, _00255_);
  or (_00259_, _00258_, _00254_);
  and (_35822_[2], _00259_, _35583_);
  and (_00260_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00261_, _32060_, _35019_);
  or (_00262_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00263_, _00262_, _35012_);
  and (_00264_, _00263_, _00261_);
  or (_00265_, _00264_, _00260_);
  and (_35822_[3], _00265_, _35583_);
  and (_00266_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00267_, _32271_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00268_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00269_, _00268_, _35012_);
  and (_00270_, _00269_, _00267_);
  or (_00271_, _00270_, _00266_);
  and (_35822_[4], _00271_, _35583_);
  and (_00272_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00273_, _32164_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00274_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_00275_, _00274_, _35012_);
  and (_00276_, _00275_, _00273_);
  or (_00277_, _00276_, _00272_);
  and (_35822_[5], _00277_, _35583_);
  and (_00278_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand (_00279_, _32335_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or (_00280_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_00281_, _00280_, _35012_);
  and (_00282_, _00281_, _00279_);
  or (_00283_, _00282_, _00278_);
  and (_35822_[6], _00283_, _35583_);
  and (_00284_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00285_, _32013_, _35019_);
  or (_00286_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_00287_, _00286_, _35012_);
  and (_00288_, _00287_, _00285_);
  or (_00289_, _00288_, _00284_);
  and (_35822_[7], _00289_, _35583_);
  and (_00290_, _35019_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_00291_, _00290_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00292_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _35012_);
  and (_00293_, _00292_, _35583_);
  and (_35822_[8], _00293_, _00291_);
  and (_00294_, _35019_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00295_, _00294_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00296_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _35012_);
  and (_00297_, _00296_, _35583_);
  and (_35822_[9], _00297_, _00295_);
  and (_00298_, _35019_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00299_, _00298_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00300_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _35012_);
  and (_00301_, _00300_, _35583_);
  and (_35822_[10], _00301_, _00299_);
  and (_00302_, _35019_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_00303_, _00302_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00304_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _35012_);
  and (_00305_, _00304_, _35583_);
  and (_35822_[11], _00305_, _00303_);
  and (_00306_, _35019_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_00307_, _00306_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00308_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _35012_);
  and (_00309_, _00308_, _35583_);
  and (_35822_[12], _00309_, _00307_);
  and (_00310_, _35019_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_00311_, _00310_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00312_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _35012_);
  and (_00313_, _00312_, _35583_);
  and (_35822_[13], _00313_, _00311_);
  and (_00314_, _35019_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_00315_, _00314_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or (_00316_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _35012_);
  and (_00317_, _00316_, _35583_);
  and (_35822_[14], _00317_, _00315_);
  nand (_00318_, _35026_, _28556_);
  or (_00319_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_00320_, _00319_, _35583_);
  and (_35826_[0], _00320_, _00318_);
  nand (_00321_, _35026_, _29242_);
  or (_00322_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00323_, _00322_, _35583_);
  and (_35826_[1], _00323_, _00321_);
  nand (_00324_, _35026_, _29887_);
  or (_00325_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00326_, _00325_, _35583_);
  and (_35826_[2], _00326_, _00324_);
  nand (_00327_, _35026_, _30092_);
  or (_00328_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_00329_, _00328_, _35583_);
  and (_35826_[3], _00329_, _00327_);
  nand (_00330_, _35026_, _30161_);
  or (_00331_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and (_00332_, _00331_, _35583_);
  and (_35826_[4], _00332_, _00330_);
  nand (_00333_, _35026_, _30236_);
  or (_00334_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and (_00335_, _00334_, _35583_);
  and (_35826_[5], _00335_, _00333_);
  nand (_00336_, _35026_, _30309_);
  or (_00337_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and (_00338_, _00337_, _35583_);
  and (_35826_[6], _00338_, _00336_);
  nand (_00339_, _35026_, _27441_);
  or (_00340_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and (_00341_, _00340_, _35583_);
  and (_35826_[7], _00341_, _00339_);
  nand (_00342_, _35026_, _30988_);
  or (_00343_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and (_00344_, _00343_, _35583_);
  and (_35826_[8], _00344_, _00342_);
  nand (_00345_, _35026_, _31019_);
  or (_00346_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and (_00347_, _00346_, _35583_);
  and (_35826_[9], _00347_, _00345_);
  nand (_00348_, _35026_, _31049_);
  or (_00349_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and (_00350_, _00349_, _35583_);
  and (_35826_[10], _00350_, _00348_);
  nand (_00351_, _35026_, _31078_);
  or (_00352_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and (_00353_, _00352_, _35583_);
  and (_35826_[11], _00353_, _00351_);
  nand (_00354_, _35026_, _31110_);
  or (_00355_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and (_00356_, _00355_, _35583_);
  and (_35826_[12], _00356_, _00354_);
  nand (_00357_, _35026_, _31143_);
  or (_00358_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and (_00359_, _00358_, _35583_);
  and (_35826_[13], _00359_, _00357_);
  nand (_00360_, _35026_, _31175_);
  or (_00361_, _35026_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and (_00362_, _00361_, _35583_);
  and (_35826_[14], _00362_, _00360_);
  nor (_35792_, _31864_, rst);
  nor (_00363_, _32087_, _32036_);
  and (_00364_, _00363_, _32359_);
  not (_00365_, _00364_);
  nor (_00366_, _32359_, _32191_);
  and (_00367_, _00366_, _00363_);
  nor (_00368_, _32359_, _32036_);
  and (_00369_, _32301_, _32191_);
  and (_00370_, _00369_, _32086_);
  and (_00371_, _00370_, _00368_);
  nor (_00372_, _00371_, _00367_);
  and (_00373_, _00372_, _00365_);
  not (_00374_, _00373_);
  and (_00375_, _30554_, _30680_);
  nor (_00376_, _00375_, _30664_);
  nor (_00377_, _30677_, _30661_);
  and (_00378_, _00377_, _00376_);
  not (_00379_, _33925_);
  and (_00380_, _33989_, _00379_);
  and (_00381_, _00380_, _00378_);
  nor (_00382_, _33991_, _33927_);
  and (_00383_, _30553_, _30551_);
  nor (_00384_, _00383_, _34103_);
  and (_00385_, _00384_, _00382_);
  and (_00386_, _00385_, _34269_);
  and (_00387_, _00386_, _00381_);
  and (_00388_, _00387_, _30638_);
  nor (_00389_, _00388_, _30331_);
  not (_00390_, _00389_);
  nand (_00391_, _00390_, _00364_);
  and (_00392_, _00391_, _31216_);
  and (_00393_, _00392_, _34473_);
  and (_00394_, _00393_, _00374_);
  not (_00395_, _32139_);
  nor (_00396_, _31361_, _31350_);
  and (_00397_, _31361_, _31350_);
  nor (_00398_, _00397_, _00396_);
  nor (_00399_, _31390_, _31376_);
  and (_00400_, _31390_, _31376_);
  nor (_00401_, _00400_, _00399_);
  nor (_00402_, _00401_, _00398_);
  and (_00403_, _00401_, _00398_);
  nor (_00404_, _00403_, _00402_);
  nor (_00405_, _31412_, _31401_);
  and (_00406_, _31412_, _31401_);
  nor (_00407_, _00406_, _00405_);
  not (_00408_, _31339_);
  nor (_00409_, _31423_, _00408_);
  and (_00410_, _31423_, _00408_);
  nor (_00411_, _00410_, _00409_);
  nor (_00412_, _00411_, _00407_);
  and (_00413_, _00411_, _00407_);
  or (_00414_, _00413_, _00412_);
  or (_00415_, _00414_, _00404_);
  nand (_00416_, _00414_, _00404_);
  and (_00417_, _00416_, _00415_);
  or (_00418_, _00417_, _00395_);
  and (_00419_, _31966_, _32246_);
  or (_00420_, _32139_, _31285_);
  and (_00421_, _00420_, _00419_);
  and (_00422_, _00421_, _00418_);
  or (_00423_, _00395_, _31230_);
  not (_00424_, _31966_);
  and (_00425_, _00424_, _32246_);
  or (_00426_, _32139_, _31294_);
  and (_00427_, _00426_, _00425_);
  and (_00428_, _00427_, _00423_);
  nor (_00429_, _31966_, _32246_);
  and (_00430_, _00429_, _32139_);
  and (_00431_, _00430_, _31274_);
  and (_00432_, _00429_, _00395_);
  and (_00433_, _00432_, _31221_);
  or (_00434_, _00433_, _00431_);
  or (_00435_, _00434_, _00428_);
  or (_00436_, _00395_, _31266_);
  nor (_00437_, _00424_, _32246_);
  or (_00438_, _32139_, _31311_);
  and (_00439_, _00438_, _00437_);
  and (_00440_, _00439_, _00436_);
  or (_00441_, _00440_, _00435_);
  or (_00442_, _00441_, _00422_);
  and (_00443_, _00442_, _00371_);
  and (_00444_, _34450_, p1in_reg[4]);
  and (_00445_, _34446_, p1_in[4]);
  or (_00446_, _00445_, _00444_);
  or (_00447_, _00446_, _00389_);
  or (_00448_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_00449_, _00448_, _00447_);
  or (_00450_, _00449_, _32139_);
  and (_00451_, _34450_, p1in_reg[0]);
  and (_00452_, _34446_, p1_in[0]);
  or (_00453_, _00452_, _00451_);
  or (_00454_, _00453_, _00389_);
  nand (_00455_, _00389_, _31588_);
  and (_00456_, _00455_, _00454_);
  or (_00457_, _00456_, _00395_);
  and (_00458_, _00457_, _00419_);
  and (_00459_, _00458_, _00450_);
  and (_00460_, _34450_, p1in_reg[3]);
  and (_00461_, _34446_, p1_in[3]);
  or (_00462_, _00461_, _00460_);
  or (_00463_, _00462_, _00389_);
  or (_00464_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_00465_, _00464_, _00463_);
  and (_00466_, _00465_, _00430_);
  or (_00467_, _00466_, _00459_);
  and (_00468_, _34450_, p1in_reg[5]);
  and (_00469_, _34446_, p1_in[5]);
  or (_00470_, _00469_, _00468_);
  or (_00471_, _00470_, _00389_);
  or (_00472_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_00473_, _00472_, _00471_);
  and (_00474_, _00473_, _00395_);
  and (_00475_, _34450_, p1in_reg[1]);
  and (_00476_, _34446_, p1_in[1]);
  or (_00477_, _00476_, _00475_);
  or (_00478_, _00477_, _00389_);
  nand (_00479_, _00389_, _31601_);
  and (_00480_, _00479_, _00478_);
  and (_00481_, _00480_, _32139_);
  or (_00482_, _00481_, _00474_);
  and (_00483_, _00482_, _00425_);
  and (_00484_, _34450_, p1in_reg[6]);
  and (_00485_, _34446_, p1_in[6]);
  or (_00486_, _00485_, _00484_);
  or (_00487_, _00486_, _00389_);
  nand (_00488_, _00389_, _31663_);
  and (_00489_, _00488_, _00487_);
  and (_00490_, _00489_, _00395_);
  and (_00491_, _34450_, p1in_reg[2]);
  and (_00492_, _34446_, p1_in[2]);
  or (_00493_, _00492_, _00491_);
  or (_00494_, _00493_, _00389_);
  nand (_00495_, _00389_, _31614_);
  and (_00496_, _00495_, _00494_);
  and (_00497_, _00496_, _32139_);
  or (_00498_, _00497_, _00490_);
  and (_00499_, _00498_, _00437_);
  and (_00500_, _34450_, p1in_reg[7]);
  and (_00501_, _34446_, p1_in[7]);
  or (_00502_, _00501_, _00500_);
  or (_00503_, _00502_, _00389_);
  nand (_00504_, _00389_, _31447_);
  and (_00505_, _00504_, _00503_);
  and (_00506_, _00505_, _00432_);
  or (_00507_, _00506_, _00499_);
  or (_00508_, _00507_, _00483_);
  or (_00509_, _00508_, _00467_);
  and (_00510_, _32359_, _32037_);
  and (_00511_, _00370_, _00510_);
  and (_00512_, _00511_, _00509_);
  and (_00513_, _34450_, p0in_reg[7]);
  and (_00514_, _34446_, p0_in[7]);
  or (_00515_, _00514_, _00513_);
  or (_00516_, _00515_, _00389_);
  nand (_00517_, _00389_, _31434_);
  and (_00518_, _00517_, _00516_);
  and (_00519_, _00518_, _00432_);
  and (_00520_, _34450_, p0in_reg[3]);
  and (_00521_, _34446_, p0_in[3]);
  or (_00522_, _00521_, _00520_);
  or (_00523_, _00522_, _00389_);
  or (_00524_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_00525_, _00524_, _00523_);
  and (_00526_, _00525_, _00430_);
  or (_00527_, _00526_, _00519_);
  and (_00528_, _34450_, p0in_reg[4]);
  and (_00529_, _34446_, p0_in[4]);
  or (_00530_, _00529_, _00528_);
  or (_00531_, _00530_, _00389_);
  or (_00532_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_00533_, _00532_, _00531_);
  or (_00534_, _00533_, _32139_);
  and (_00535_, _34450_, p0in_reg[0]);
  and (_00536_, _34446_, p0_in[0]);
  or (_00537_, _00536_, _00535_);
  or (_00538_, _00537_, _00389_);
  nand (_00539_, _00389_, _31489_);
  and (_00540_, _00539_, _00538_);
  or (_00541_, _00540_, _00395_);
  and (_00542_, _00541_, _00419_);
  and (_00543_, _00542_, _00534_);
  and (_00544_, _34450_, p0in_reg[6]);
  and (_00545_, _34446_, p0_in[6]);
  or (_00546_, _00545_, _00544_);
  or (_00547_, _00546_, _00389_);
  nand (_00548_, _00389_, _31570_);
  and (_00549_, _00548_, _00547_);
  and (_00550_, _00549_, _00395_);
  and (_00551_, _34450_, p0in_reg[2]);
  and (_00552_, _34446_, p0_in[2]);
  or (_00553_, _00552_, _00551_);
  or (_00554_, _00553_, _00389_);
  nand (_00555_, _00389_, _31525_);
  and (_00556_, _00555_, _00554_);
  and (_00557_, _00556_, _32139_);
  or (_00558_, _00557_, _00550_);
  and (_00559_, _00558_, _00437_);
  or (_00560_, _00559_, _00543_);
  and (_00561_, _34450_, p0in_reg[5]);
  and (_00562_, _34446_, p0_in[5]);
  or (_00563_, _00562_, _00561_);
  or (_00564_, _00563_, _00389_);
  or (_00565_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_00566_, _00565_, _00564_);
  and (_00567_, _00566_, _00395_);
  and (_00568_, _34450_, p0in_reg[1]);
  and (_00569_, _34446_, p0_in[1]);
  or (_00570_, _00569_, _00568_);
  or (_00571_, _00570_, _00389_);
  nand (_00572_, _00389_, _31509_);
  and (_00573_, _00572_, _00571_);
  and (_00574_, _00573_, _32139_);
  or (_00575_, _00574_, _00567_);
  and (_00576_, _00575_, _00425_);
  or (_00577_, _00576_, _00560_);
  or (_00578_, _00577_, _00527_);
  and (_00579_, _32300_, _32191_);
  and (_00580_, _00579_, _00364_);
  and (_00581_, _00580_, _00578_);
  or (_00582_, _00581_, _00512_);
  and (_00583_, _00363_, _32300_);
  and (_00584_, _00395_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_00585_, _32139_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_00586_, _00585_, _00584_);
  and (_00587_, _00586_, _00425_);
  and (_00588_, _00437_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00589_, _00588_, _00395_);
  and (_00590_, _00419_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_00591_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_00592_, _00591_, _00590_);
  or (_00593_, _00592_, _00589_);
  and (_00594_, _00437_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_00595_, _00594_, _32139_);
  and (_00596_, _00419_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_00597_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_00598_, _00597_, _00596_);
  or (_00599_, _00598_, _00595_);
  and (_00600_, _00599_, _00593_);
  or (_00601_, _00600_, _00587_);
  and (_00602_, _00601_, _00366_);
  and (_00603_, _34450_, p2in_reg[7]);
  and (_00604_, _34446_, p2_in[7]);
  or (_00605_, _00604_, _00603_);
  or (_00606_, _00605_, _00389_);
  nand (_00607_, _00389_, _31466_);
  and (_00608_, _00607_, _00606_);
  and (_00609_, _00608_, _00432_);
  and (_00610_, _34450_, p2in_reg[4]);
  and (_00611_, _34446_, p2_in[4]);
  or (_00612_, _00611_, _00610_);
  or (_00613_, _00612_, _00389_);
  or (_00614_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_00615_, _00614_, _00613_);
  or (_00616_, _00615_, _32139_);
  and (_00617_, _34450_, p2in_reg[0]);
  and (_00618_, _34446_, p2_in[0]);
  or (_00619_, _00618_, _00617_);
  or (_00620_, _00619_, _00389_);
  nand (_00621_, _00389_, _31676_);
  and (_00622_, _00621_, _00620_);
  or (_00623_, _00622_, _00395_);
  and (_00624_, _00623_, _00419_);
  and (_00625_, _00624_, _00616_);
  and (_00626_, _34450_, p2in_reg[3]);
  and (_00627_, _34446_, p2_in[3]);
  or (_00628_, _00627_, _00626_);
  or (_00629_, _00628_, _00389_);
  or (_00630_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_00631_, _00630_, _00629_);
  and (_00632_, _00631_, _00430_);
  or (_00633_, _00632_, _00625_);
  or (_00634_, _00633_, _00609_);
  and (_00635_, _34450_, p2in_reg[6]);
  and (_00636_, _34446_, p2_in[6]);
  or (_00637_, _00636_, _00635_);
  or (_00638_, _00637_, _00389_);
  nand (_00639_, _00389_, _31751_);
  and (_00640_, _00639_, _00638_);
  and (_00641_, _00640_, _00395_);
  and (_00642_, _34450_, p2in_reg[2]);
  and (_00643_, _34446_, p2_in[2]);
  or (_00644_, _00643_, _00642_);
  or (_00645_, _00644_, _00389_);
  nand (_00646_, _00389_, _31702_);
  and (_00647_, _00646_, _00645_);
  and (_00648_, _00647_, _32139_);
  or (_00649_, _00648_, _00641_);
  and (_00650_, _00649_, _00437_);
  and (_00651_, _34450_, p2in_reg[5]);
  and (_00652_, _34446_, p2_in[5]);
  or (_00653_, _00652_, _00651_);
  or (_00654_, _00653_, _00389_);
  or (_00655_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_00656_, _00655_, _00654_);
  and (_00657_, _00656_, _00395_);
  and (_00658_, _34450_, p2in_reg[1]);
  and (_00659_, _34446_, p2_in[1]);
  or (_00660_, _00659_, _00658_);
  or (_00661_, _00660_, _00389_);
  nand (_00662_, _00389_, _31689_);
  and (_00663_, _00662_, _00661_);
  and (_00664_, _00663_, _32139_);
  or (_00665_, _00664_, _00657_);
  and (_00666_, _00665_, _00425_);
  or (_00667_, _00666_, _00650_);
  or (_00668_, _00667_, _00634_);
  and (_00669_, _32359_, _32192_);
  and (_00670_, _00669_, _00668_);
  or (_00671_, _00670_, _00602_);
  and (_00672_, _00671_, _00583_);
  and (_00673_, _00367_, _32301_);
  and (_00674_, _00432_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_00675_, _32139_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_00676_, _32139_, _28589_);
  and (_00677_, _00676_, _00419_);
  and (_00678_, _00677_, _00675_);
  and (_00679_, _00430_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_00680_, _00679_, _00678_);
  or (_00681_, _00680_, _00674_);
  nor (_00682_, _32139_, _30312_);
  and (_00683_, _32139_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_00684_, _00683_, _00682_);
  and (_00685_, _00684_, _00437_);
  nor (_00686_, _32139_, _30239_);
  and (_00687_, _32139_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_00688_, _00687_, _00686_);
  and (_00689_, _00688_, _00425_);
  or (_00690_, _00689_, _00685_);
  or (_00691_, _00690_, _00681_);
  and (_00692_, _00691_, _00673_);
  nor (_00693_, _00373_, _27474_);
  and (_00694_, _00693_, _34486_);
  and (_00695_, _34450_, p3in_reg[7]);
  and (_00696_, _34446_, p3_in[7]);
  or (_00697_, _00696_, _00695_);
  or (_00698_, _00697_, _00389_);
  nand (_00699_, _00389_, _31482_);
  and (_00700_, _00699_, _00698_);
  and (_00701_, _00700_, _00432_);
  and (_00702_, _34450_, p3in_reg[4]);
  and (_00703_, _34446_, p3_in[4]);
  or (_00704_, _00703_, _00702_);
  or (_00705_, _00704_, _00389_);
  or (_00706_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_00707_, _00706_, _00705_);
  or (_00708_, _00707_, _32139_);
  and (_00709_, _34450_, p3in_reg[0]);
  and (_00710_, _34446_, p3_in[0]);
  or (_00711_, _00710_, _00709_);
  or (_00712_, _00711_, _00389_);
  nand (_00713_, _00389_, _31764_);
  and (_00714_, _00713_, _00712_);
  or (_00715_, _00714_, _00395_);
  and (_00716_, _00715_, _00419_);
  and (_00717_, _00716_, _00708_);
  and (_00718_, _34450_, p3in_reg[3]);
  and (_00719_, _34446_, p3_in[3]);
  or (_00720_, _00719_, _00718_);
  or (_00721_, _00720_, _00389_);
  or (_00722_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_00723_, _00722_, _00721_);
  and (_00724_, _00723_, _00430_);
  or (_00725_, _00724_, _00717_);
  or (_00726_, _00725_, _00701_);
  and (_00727_, _34450_, p3in_reg[6]);
  and (_00728_, _34446_, p3_in[6]);
  or (_00729_, _00728_, _00727_);
  or (_00730_, _00729_, _00389_);
  nand (_00731_, _00389_, _31839_);
  and (_00732_, _00731_, _00730_);
  and (_00733_, _00732_, _00395_);
  and (_00734_, _34450_, p3in_reg[2]);
  and (_00735_, _34446_, p3_in[2]);
  or (_00736_, _00735_, _00734_);
  or (_00737_, _00736_, _00389_);
  nand (_00738_, _00389_, _31790_);
  and (_00739_, _00738_, _00737_);
  and (_00740_, _00739_, _32139_);
  or (_00741_, _00740_, _00733_);
  and (_00742_, _00741_, _00437_);
  and (_00743_, _34450_, p3in_reg[5]);
  and (_00744_, _34446_, p3_in[5]);
  or (_00745_, _00744_, _00743_);
  or (_00746_, _00745_, _00389_);
  or (_00747_, _00390_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_00748_, _00747_, _00746_);
  and (_00749_, _00748_, _00395_);
  and (_00750_, _34450_, p3in_reg[1]);
  and (_00751_, _34446_, p3_in[1]);
  or (_00752_, _00751_, _00750_);
  or (_00753_, _00752_, _00389_);
  nand (_00754_, _00389_, _31777_);
  and (_00755_, _00754_, _00753_);
  and (_00756_, _00755_, _32139_);
  or (_00757_, _00756_, _00749_);
  and (_00758_, _00757_, _00425_);
  or (_00759_, _00758_, _00742_);
  or (_00760_, _00759_, _00726_);
  and (_00761_, _00669_, _32301_);
  and (_00762_, _00761_, _00363_);
  and (_00763_, _00762_, _00760_);
  or (_00764_, _00763_, _00694_);
  or (_00765_, _00764_, _00692_);
  or (_00766_, _00765_, _00672_);
  or (_00767_, _00766_, _00582_);
  or (_00768_, _00767_, _00443_);
  nand (_00769_, _00694_, _28062_);
  nand (_00770_, _00769_, _00768_);
  and (_00771_, _00583_, _00366_);
  and (_00772_, _00771_, _31316_);
  nor (_00773_, _00772_, _00770_);
  or (_00774_, _32139_, _31412_);
  or (_00775_, _00395_, _31361_);
  and (_00776_, _00775_, _00425_);
  and (_00777_, _00776_, _00774_);
  or (_00778_, _32139_, _31423_);
  nand (_00779_, _32139_, _31376_);
  and (_00780_, _00779_, _00437_);
  and (_00781_, _00780_, _00778_);
  or (_00782_, _00395_, _31350_);
  or (_00783_, _32139_, _31401_);
  and (_00784_, _00783_, _00419_);
  and (_00785_, _00784_, _00782_);
  or (_00786_, _00785_, _00781_);
  and (_00787_, _00432_, _31339_);
  not (_00788_, _31390_);
  and (_00789_, _00430_, _00788_);
  or (_00790_, _00789_, _00787_);
  or (_00791_, _00790_, _00786_);
  or (_00792_, _00791_, _00777_);
  and (_00793_, _00792_, _00772_);
  or (_00794_, _00793_, _00773_);
  or (_00795_, _00794_, _00394_);
  not (_00796_, _00432_);
  nor (_00797_, _00796_, _30808_);
  or (_00798_, _32139_, _32313_);
  or (_00799_, _00395_, _30770_);
  and (_00800_, _00799_, _00437_);
  and (_00801_, _00800_, _00798_);
  or (_00802_, _32139_, _32248_);
  nand (_00803_, _32139_, _30785_);
  and (_00804_, _00803_, _00419_);
  and (_00805_, _00804_, _00802_);
  or (_00806_, _00805_, _00801_);
  and (_00807_, _00430_, _32039_);
  nor (_00808_, _00395_, _30777_);
  nor (_00809_, _32139_, _30749_);
  or (_00810_, _00809_, _00808_);
  and (_00811_, _00810_, _00425_);
  or (_00812_, _00811_, _00807_);
  or (_00813_, _00812_, _00806_);
  nor (_00814_, _00813_, _00797_);
  nand (_00815_, _00814_, _00394_);
  and (_00816_, _00815_, _35583_);
  and (_35961_, _00816_, _00795_);
  and (_00817_, _00579_, _00510_);
  and (_00818_, _32086_, _32139_);
  and (_00819_, _00818_, _00429_);
  and (_00820_, _00819_, _00817_);
  and (_00821_, _00820_, _30860_);
  and (_00822_, _32300_, _32192_);
  and (_00823_, _00818_, _00419_);
  and (_00824_, _00823_, _00368_);
  and (_00825_, _00824_, _00822_);
  and (_00826_, _00825_, _31313_);
  and (_00827_, _00824_, _00369_);
  and (_00828_, _00827_, _31211_);
  or (_00829_, _00828_, _00826_);
  nor (_00830_, _00829_, _00821_);
  nor (_00831_, _00830_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_00832_, _00831_);
  and (_00833_, _00825_, _31316_);
  and (_00834_, _00796_, _31326_);
  and (_00835_, _00834_, _34473_);
  nor (_00836_, _00835_, _00833_);
  and (_00837_, _00836_, _34489_);
  and (_00838_, _00837_, _00832_);
  and (_00839_, _00818_, _00437_);
  and (_00840_, _00839_, _00817_);
  and (_00841_, _00840_, _30860_);
  or (_00842_, _00841_, rst);
  nor (_35962_, _00842_, _00838_);
  not (_00843_, _00841_);
  and (_00844_, _00840_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nor (_00845_, _32300_, _32191_);
  and (_00846_, _00845_, _00824_);
  and (_00847_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_00848_, _00820_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_00849_, _00848_, _00847_);
  and (_00850_, _00818_, _00425_);
  and (_00851_, _00850_, _00817_);
  and (_00852_, _00851_, _30810_);
  and (_00853_, _00845_, _00510_);
  and (_00854_, _00853_, _00823_);
  and (_00855_, _00854_, _00700_);
  or (_00856_, _00855_, _00852_);
  or (_00857_, _00856_, _00849_);
  or (_00858_, _00857_, _00844_);
  and (_00859_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_00860_, _00823_, _00510_);
  and (_00861_, _00860_, _00369_);
  and (_00862_, _00861_, _00505_);
  and (_00863_, _00822_, _00510_);
  and (_00864_, _00863_, _00823_);
  and (_00865_, _00864_, _00608_);
  or (_00866_, _00865_, _00862_);
  and (_00867_, _00827_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_00868_, _00817_, _00823_);
  and (_00869_, _00868_, _00518_);
  or (_00870_, _00869_, _00867_);
  or (_00871_, _00870_, _00866_);
  or (_00872_, _00871_, _00859_);
  or (_00873_, _00872_, _00858_);
  and (_00874_, _00873_, _00838_);
  nor (_00875_, _00838_, _16930_);
  or (_00876_, _00875_, _00874_);
  and (_00877_, _00876_, _00843_);
  nor (_00878_, _00843_, _27441_);
  or (_00879_, _00878_, _00877_);
  and (_35963_[7], _00879_, _35583_);
  and (_00880_, _00827_, _00417_);
  and (_00881_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_00882_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_00883_, _00882_, _00881_);
  and (_00884_, _00861_, _00456_);
  and (_00885_, _00580_, _00430_);
  and (_00886_, _00885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_00887_, _00886_, _00884_);
  or (_00888_, _00887_, _00883_);
  and (_00889_, _00868_, _00540_);
  and (_00890_, _00840_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_00891_, _00851_, _31937_);
  or (_00892_, _00891_, _00890_);
  or (_00893_, _00892_, _00889_);
  and (_00894_, _00860_, _00845_);
  and (_00895_, _00894_, _00714_);
  and (_00896_, _00860_, _00822_);
  and (_00897_, _00896_, _00622_);
  or (_00898_, _00897_, _00895_);
  or (_00899_, _00898_, _00893_);
  nor (_00900_, _00899_, _00888_);
  nand (_00901_, _00900_, _00838_);
  or (_00902_, _00901_, _00880_);
  or (_00903_, _00838_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_00904_, _00903_, _00902_);
  or (_00905_, _00904_, _00841_);
  nand (_00906_, _00841_, _28556_);
  and (_00907_, _00906_, _35583_);
  and (_35963_[0], _00907_, _00905_);
  and (_00908_, _00840_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_00909_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_00910_, _00820_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_00911_, _00910_, _00909_);
  and (_00912_, _00851_, _32200_);
  and (_00913_, _00854_, _00755_);
  or (_00914_, _00913_, _00912_);
  or (_00915_, _00914_, _00911_);
  or (_00916_, _00915_, _00908_);
  and (_00917_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_00918_, _00861_, _00480_);
  and (_00919_, _00864_, _00663_);
  or (_00920_, _00919_, _00918_);
  and (_00921_, _00868_, _00573_);
  and (_00922_, _00827_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_00923_, _00922_, _00921_);
  or (_00924_, _00923_, _00920_);
  or (_00925_, _00924_, _00917_);
  or (_00926_, _00925_, _00916_);
  and (_00927_, _00926_, _00838_);
  nor (_00928_, _00838_, _16756_);
  or (_00929_, _00928_, _00927_);
  and (_00930_, _00929_, _00843_);
  nor (_00931_, _00843_, _29242_);
  or (_00932_, _00931_, _00930_);
  and (_35963_[1], _00932_, _35583_);
  and (_00933_, _00827_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_00934_, _00894_, _00739_);
  and (_00935_, _00885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_00936_, _00935_, _00934_);
  or (_00937_, _00936_, _00933_);
  and (_00938_, _00840_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_00939_, _00851_, _32117_);
  and (_00940_, _00868_, _00556_);
  or (_00941_, _00940_, _00939_);
  or (_00942_, _00941_, _00938_);
  and (_00943_, _00861_, _00496_);
  and (_00944_, _00896_, _00647_);
  or (_00945_, _00944_, _00943_);
  and (_00946_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_00947_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_00948_, _00947_, _00946_);
  or (_00949_, _00948_, _00945_);
  or (_00950_, _00949_, _00942_);
  or (_00951_, _00950_, _00937_);
  and (_00952_, _00951_, _00838_);
  nor (_00953_, _00838_, _15431_);
  or (_00954_, _00953_, _00952_);
  and (_00955_, _00954_, _00843_);
  nor (_00956_, _00843_, _29887_);
  or (_00957_, _00956_, _00955_);
  and (_35963_[2], _00957_, _35583_);
  and (_00958_, _00840_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_00959_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_00960_, _00820_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_00961_, _00960_, _00959_);
  and (_00962_, _00851_, _32063_);
  and (_00963_, _00854_, _00723_);
  or (_00964_, _00963_, _00962_);
  or (_00965_, _00964_, _00961_);
  or (_00966_, _00965_, _00958_);
  and (_00967_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_00968_, _00861_, _00465_);
  and (_00969_, _00864_, _00631_);
  or (_00970_, _00969_, _00968_);
  and (_00971_, _00827_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_00972_, _00868_, _00525_);
  or (_00973_, _00972_, _00971_);
  or (_00974_, _00973_, _00970_);
  or (_00975_, _00974_, _00967_);
  or (_00976_, _00975_, _00966_);
  and (_00977_, _00976_, _00838_);
  nor (_00978_, _00838_, _16454_);
  or (_00979_, _00978_, _00977_);
  and (_00980_, _00979_, _00843_);
  nor (_00981_, _00843_, _30092_);
  or (_00982_, _00981_, _00980_);
  and (_35963_[3], _00982_, _35583_);
  and (_00983_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_00984_, _00894_, _00707_);
  and (_00985_, _00885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_00986_, _00985_, _00984_);
  or (_00987_, _00986_, _00983_);
  and (_00988_, _00840_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_00989_, _00851_, _32274_);
  and (_00990_, _00868_, _00533_);
  or (_00991_, _00990_, _00989_);
  or (_00992_, _00991_, _00988_);
  and (_00993_, _00861_, _00449_);
  and (_00994_, _00896_, _00615_);
  or (_00995_, _00994_, _00993_);
  and (_00996_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_00997_, _00827_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_00998_, _00997_, _00996_);
  or (_00999_, _00998_, _00995_);
  or (_01000_, _00999_, _00992_);
  or (_01001_, _01000_, _00987_);
  and (_01002_, _01001_, _00838_);
  nor (_01003_, _00838_, _15627_);
  or (_01004_, _01003_, _01002_);
  and (_01005_, _01004_, _00843_);
  nor (_01006_, _00843_, _30161_);
  or (_01007_, _01006_, _01005_);
  and (_35963_[4], _01007_, _35583_);
  and (_01008_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01009_, _00894_, _00748_);
  and (_01010_, _00885_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_01011_, _01010_, _01009_);
  or (_01012_, _01011_, _01008_);
  and (_01013_, _00840_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_01014_, _00851_, _32171_);
  and (_01015_, _00868_, _00566_);
  or (_01016_, _01015_, _01014_);
  or (_01017_, _01016_, _01013_);
  and (_01018_, _00861_, _00473_);
  and (_01019_, _00896_, _00656_);
  or (_01020_, _01019_, _01018_);
  and (_01021_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01022_, _00827_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_01023_, _01022_, _01021_);
  or (_01024_, _01023_, _01020_);
  or (_01025_, _01024_, _01017_);
  or (_01026_, _01025_, _01012_);
  and (_01027_, _01026_, _00838_);
  nor (_01028_, _00838_, _16597_);
  or (_01029_, _01028_, _01027_);
  and (_01030_, _01029_, _00843_);
  nor (_01031_, _00843_, _30236_);
  or (_01032_, _01031_, _01030_);
  and (_35963_[5], _01032_, _35583_);
  and (_01033_, _00840_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_01034_, _00846_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01035_, _00820_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_01036_, _01035_, _01034_);
  and (_01037_, _00851_, _32337_);
  and (_01038_, _00854_, _00732_);
  or (_01039_, _01038_, _01037_);
  or (_01040_, _01039_, _01036_);
  or (_01041_, _01040_, _01033_);
  and (_01042_, _00825_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_01043_, _00861_, _00489_);
  and (_01044_, _00864_, _00640_);
  or (_01045_, _01044_, _01043_);
  and (_01046_, _00827_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_01047_, _00868_, _00549_);
  or (_01048_, _01047_, _01046_);
  or (_01049_, _01048_, _01045_);
  or (_01050_, _01049_, _01042_);
  or (_01051_, _01050_, _01041_);
  and (_01052_, _01051_, _00838_);
  nor (_01053_, _00838_, _15964_);
  or (_01054_, _01053_, _01052_);
  and (_01055_, _01054_, _00843_);
  nor (_01056_, _00843_, _30309_);
  or (_01057_, _01056_, _01055_);
  and (_35963_[6], _01057_, _35583_);
  and (_35828_, _32367_, _35583_);
  nor (_35829_[7], _32000_, rst);
  nor (_35831_[2], _32139_, rst);
  and (_35829_[0], _31916_, _35583_);
  nor (_35829_[1], _32213_, rst);
  and (_35829_[2], _32102_, _35583_);
  and (_35829_[3], _32048_, _35583_);
  nor (_35829_[4], _32258_, rst);
  nor (_35829_[5], _32151_, rst);
  nor (_35829_[6], _32331_, rst);
  nor (_35831_[0], _31966_, rst);
  nor (_35831_[1], _32246_, rst);
  not (_01058_, _33622_);
  nor (_01059_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_01060_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01061_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01060_);
  nor (_01062_, _01061_, _01059_);
  not (_01063_, _01062_);
  nor (_01064_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01065_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01060_);
  nor (_01066_, _01065_, _01064_);
  nor (_01067_, _01066_, _01063_);
  nor (_01068_, _01066_, _01062_);
  not (_01069_, _01068_);
  nor (_01070_, _35263_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01071_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01060_);
  nor (_01072_, _01071_, _01070_);
  and (_01073_, _01072_, _01069_);
  nor (_01074_, _01072_, _01069_);
  nor (_01075_, _01074_, _01073_);
  nor (_01076_, _35281_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_01077_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01060_);
  nor (_01078_, _01077_, _01076_);
  and (_01079_, _01078_, _01075_);
  and (_01080_, _01079_, _01067_);
  and (_01081_, _01080_, _01058_);
  not (_01082_, _33663_);
  and (_01083_, _01066_, _01063_);
  and (_01084_, _01079_, _01083_);
  and (_01085_, _01084_, _01082_);
  not (_01086_, _33704_);
  and (_01087_, _01066_, _01062_);
  and (_01088_, _01079_, _01087_);
  and (_01089_, _01088_, _01086_);
  or (_01090_, _01089_, _01085_);
  or (_01091_, _01090_, _01081_);
  not (_01092_, _33417_);
  and (_01093_, _01072_, _01068_);
  not (_01094_, _01078_);
  and (_01095_, _01094_, _01093_);
  and (_01096_, _01095_, _01092_);
  not (_01097_, _33581_);
  and (_01098_, _01078_, _01074_);
  and (_01099_, _01098_, _01097_);
  or (_01100_, _01099_, _01096_);
  or (_01101_, _01100_, _01091_);
  not (_01102_, _33376_);
  nor (_01103_, _01078_, _01073_);
  and (_01104_, _01103_, _01087_);
  and (_01105_, _01104_, _01102_);
  not (_01106_, _33335_);
  and (_01107_, _01083_, _01103_);
  and (_01108_, _01107_, _01106_);
  or (_01109_, _01108_, _01105_);
  not (_01110_, _33294_);
  and (_01111_, _01067_, _01103_);
  and (_01112_, _01111_, _01110_);
  or (_01113_, _01112_, _01109_);
  not (_01114_, _33253_);
  and (_01115_, _01094_, _01074_);
  and (_01116_, _01115_, _01114_);
  not (_01117_, _33171_);
  and (_01118_, _01078_, _01073_);
  nor (_01119_, _01103_, _01118_);
  nor (_01120_, _01119_, _01075_);
  and (_01121_, _01083_, _01120_);
  and (_01122_, _01121_, _01117_);
  or (_01123_, _01122_, _01116_);
  or (_01124_, _01123_, _01113_);
  or (_01125_, _01124_, _01101_);
  not (_01126_, _33458_);
  not (_01127_, _01075_);
  and (_01128_, _01119_, _01127_);
  and (_01129_, _01067_, _01128_);
  and (_01130_, _01129_, _01126_);
  not (_01131_, _33540_);
  and (_01132_, _01128_, _01087_);
  and (_01133_, _01132_, _01131_);
  not (_01134_, _33499_);
  and (_01135_, _01083_, _01128_);
  and (_01136_, _01135_, _01134_);
  or (_01137_, _01136_, _01133_);
  or (_01138_, _01137_, _01130_);
  not (_01139_, _33130_);
  and (_01140_, _01120_, _01067_);
  and (_01141_, _01140_, _01139_);
  not (_01142_, _33212_);
  and (_01143_, _01120_, _01087_);
  and (_01144_, _01143_, _01142_);
  or (_01145_, _01144_, _01141_);
  not (_01146_, _33745_);
  and (_01147_, _01078_, _01093_);
  and (_01148_, _01147_, _01146_);
  or (_01149_, _01148_, _01145_);
  or (_01150_, _01149_, _01138_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _01150_, _01125_);
  and (_01151_, _01132_, _01126_);
  and (_01152_, _01135_, _01092_);
  and (_01153_, _01143_, _01139_);
  or (_01154_, _01153_, _01152_);
  or (_01155_, _01154_, _01151_);
  and (_01156_, _01084_, _01097_);
  and (_01157_, _01098_, _01134_);
  and (_01158_, _01147_, _01082_);
  or (_01159_, _01158_, _01157_);
  and (_01160_, _01095_, _01106_);
  and (_01161_, _01115_, _01117_);
  or (_01162_, _01161_, _01160_);
  or (_01163_, _01162_, _01159_);
  or (_01164_, _01163_, _01156_);
  and (_01165_, _01080_, _01131_);
  and (_01166_, _01088_, _01058_);
  or (_01167_, _01166_, _01165_);
  or (_01168_, _01167_, _01164_);
  and (_01169_, _01121_, _01146_);
  and (_01170_, _01104_, _01110_);
  and (_01171_, _01107_, _01114_);
  and (_01172_, _01111_, _01142_);
  or (_01173_, _01172_, _01171_);
  or (_01174_, _01173_, _01170_);
  or (_01175_, _01174_, _01169_);
  and (_01176_, _01140_, _01086_);
  and (_01177_, _01129_, _01102_);
  or (_01178_, _01177_, _01176_);
  or (_01179_, _01178_, _01175_);
  or (_01180_, _01179_, _01168_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _01180_, _01155_);
  and (_01181_, _01098_, _01131_);
  and (_01182_, _01132_, _01134_);
  or (_01183_, _01182_, _01181_);
  and (_01184_, _01135_, _01126_);
  and (_01185_, _01129_, _01092_);
  or (_01186_, _01185_, _01184_);
  or (_01187_, _01186_, _01183_);
  and (_01188_, _01140_, _01146_);
  and (_01189_, _01088_, _01082_);
  and (_01190_, _01080_, _01097_);
  and (_01191_, _01084_, _01058_);
  or (_01192_, _01191_, _01190_);
  or (_01193_, _01192_, _01189_);
  or (_01194_, _01193_, _01188_);
  or (_01195_, _01194_, _01187_);
  and (_01196_, _01143_, _01117_);
  and (_01197_, _01107_, _01110_);
  and (_01198_, _01111_, _01114_);
  or (_01199_, _01198_, _01197_);
  and (_01200_, _01095_, _01102_);
  and (_01201_, _01104_, _01106_);
  or (_01202_, _01201_, _01200_);
  or (_01203_, _01202_, _01199_);
  or (_01204_, _01203_, _01196_);
  and (_01205_, _01147_, _01086_);
  and (_01206_, _01121_, _01139_);
  and (_01207_, _01115_, _01142_);
  or (_01208_, _01207_, _01206_);
  or (_01209_, _01208_, _01205_);
  or (_01210_, _01209_, _01204_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _01210_, _01195_);
  and (_01211_, _01098_, _01126_);
  and (_01212_, _01080_, _01134_);
  and (_01213_, _01084_, _01131_);
  or (_01214_, _01213_, _01212_);
  or (_01215_, _01214_, _01211_);
  and (_01216_, _01140_, _01082_);
  and (_01217_, _01132_, _01092_);
  or (_01218_, _01217_, _01216_);
  or (_01219_, _01218_, _01215_);
  and (_01220_, _01135_, _01102_);
  and (_01221_, _01115_, _01139_);
  and (_01222_, _01111_, _01117_);
  and (_01223_, _01107_, _01142_);
  or (_01224_, _01223_, _01222_);
  or (_01225_, _01224_, _01221_);
  or (_01226_, _01225_, _01220_);
  or (_01227_, _01226_, _01219_);
  and (_01228_, _01088_, _01097_);
  and (_01229_, _01143_, _01146_);
  and (_01230_, _01121_, _01086_);
  or (_01231_, _01230_, _01229_);
  or (_01232_, _01231_, _01228_);
  and (_01233_, _01147_, _01058_);
  and (_01234_, _01129_, _01106_);
  and (_01235_, _01095_, _01110_);
  and (_01236_, _01104_, _01114_);
  or (_01237_, _01236_, _01235_);
  or (_01238_, _01237_, _01234_);
  or (_01239_, _01238_, _01233_);
  or (_01240_, _01239_, _01232_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _01240_, _01227_);
  not (_01241_, _33545_);
  and (_01242_, _01132_, _01241_);
  not (_01243_, _33463_);
  and (_01244_, _01129_, _01243_);
  not (_01245_, _33176_);
  and (_01246_, _01121_, _01245_);
  or (_01247_, _01246_, _01244_);
  or (_01248_, _01247_, _01242_);
  not (_01249_, _33668_);
  and (_01250_, _01084_, _01249_);
  not (_01251_, _33750_);
  and (_01252_, _01147_, _01251_);
  not (_01253_, _33422_);
  and (_01254_, _01095_, _01253_);
  or (_01255_, _01254_, _01252_);
  not (_01256_, _33586_);
  and (_01257_, _01098_, _01256_);
  not (_01258_, _33258_);
  and (_01259_, _01115_, _01258_);
  or (_01260_, _01259_, _01257_);
  or (_01261_, _01260_, _01255_);
  or (_01262_, _01261_, _01250_);
  not (_01263_, _33709_);
  and (_01264_, _01088_, _01263_);
  not (_01265_, _33627_);
  and (_01266_, _01080_, _01265_);
  or (_01267_, _01266_, _01264_);
  or (_01268_, _01267_, _01262_);
  not (_01269_, _33135_);
  and (_01270_, _01140_, _01269_);
  not (_01271_, _33217_);
  and (_01272_, _01143_, _01271_);
  or (_01273_, _01272_, _01270_);
  not (_01274_, _33504_);
  and (_01275_, _01135_, _01274_);
  not (_01276_, _33381_);
  and (_01277_, _01104_, _01276_);
  not (_01278_, _33340_);
  and (_01279_, _01107_, _01278_);
  or (_01280_, _01279_, _01277_);
  not (_01281_, _33299_);
  and (_01282_, _01111_, _01281_);
  or (_01283_, _01282_, _01280_);
  or (_01284_, _01283_, _01275_);
  or (_01285_, _01284_, _01273_);
  or (_01286_, _01285_, _01268_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _01286_, _01248_);
  not (_01287_, _33550_);
  and (_01288_, _01132_, _01287_);
  not (_01289_, _33509_);
  and (_01290_, _01135_, _01289_);
  or (_01291_, _01290_, _01288_);
  not (_01292_, _33427_);
  and (_01293_, _01095_, _01292_);
  not (_01294_, _33468_);
  and (_01295_, _01129_, _01294_);
  or (_01296_, _01295_, _01293_);
  or (_01297_, _01296_, _01291_);
  not (_01298_, _33345_);
  and (_01299_, _01107_, _01298_);
  not (_01300_, _33386_);
  and (_01301_, _01104_, _01300_);
  or (_01302_, _01301_, _01299_);
  not (_01303_, _33304_);
  and (_01304_, _01111_, _01303_);
  or (_01305_, _01304_, _01302_);
  not (_01306_, _33181_);
  and (_01307_, _01121_, _01306_);
  not (_01308_, _33263_);
  and (_01309_, _01115_, _01308_);
  or (_01310_, _01309_, _01307_);
  or (_01311_, _01310_, _01305_);
  or (_01312_, _01311_, _01297_);
  not (_01313_, _33673_);
  and (_01314_, _01084_, _01313_);
  not (_01315_, _33714_);
  and (_01316_, _01088_, _01315_);
  or (_01317_, _01316_, _01314_);
  not (_01318_, _33591_);
  and (_01319_, _01098_, _01318_);
  not (_01320_, _33632_);
  and (_01321_, _01080_, _01320_);
  or (_01322_, _01321_, _01319_);
  or (_01323_, _01322_, _01317_);
  not (_01324_, _33755_);
  and (_01325_, _01147_, _01324_);
  not (_01326_, _33140_);
  and (_01327_, _01140_, _01326_);
  not (_01328_, _33222_);
  and (_01329_, _01143_, _01328_);
  or (_01330_, _01329_, _01327_);
  or (_01331_, _01330_, _01325_);
  or (_01332_, _01331_, _01323_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _01332_, _01312_);
  not (_01333_, _33514_);
  and (_01334_, _01135_, _01333_);
  not (_01335_, _33186_);
  and (_01336_, _01121_, _01335_);
  not (_01337_, _33227_);
  and (_01338_, _01143_, _01337_);
  or (_01339_, _01338_, _01336_);
  or (_01340_, _01339_, _01334_);
  not (_01341_, _33719_);
  and (_01342_, _01088_, _01341_);
  not (_01343_, _33678_);
  and (_01344_, _01084_, _01343_);
  or (_01345_, _01344_, _01342_);
  not (_01346_, _33637_);
  and (_01347_, _01080_, _01346_);
  not (_01348_, _33760_);
  and (_01349_, _01147_, _01348_);
  not (_01350_, _33432_);
  and (_01351_, _01095_, _01350_);
  or (_01352_, _01351_, _01349_);
  not (_01353_, _33596_);
  and (_01354_, _01098_, _01353_);
  not (_01355_, _33268_);
  and (_01356_, _01115_, _01355_);
  or (_01357_, _01356_, _01354_);
  or (_01358_, _01357_, _01352_);
  or (_01359_, _01358_, _01347_);
  or (_01360_, _01359_, _01345_);
  not (_01361_, _33145_);
  and (_01362_, _01140_, _01361_);
  not (_01363_, _33309_);
  and (_01364_, _01111_, _01363_);
  not (_01365_, _33350_);
  and (_01366_, _01107_, _01365_);
  not (_01367_, _33391_);
  and (_01368_, _01104_, _01367_);
  or (_01369_, _01368_, _01366_);
  or (_01370_, _01369_, _01364_);
  or (_01371_, _01370_, _01362_);
  not (_01372_, _33555_);
  and (_01373_, _01132_, _01372_);
  not (_01374_, _33473_);
  and (_01375_, _01129_, _01374_);
  or (_01376_, _01375_, _01373_);
  or (_01377_, _01376_, _01371_);
  or (_01378_, _01377_, _01360_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _01378_, _01340_);
  not (_01379_, _33232_);
  and (_01380_, _01143_, _01379_);
  not (_01381_, _33150_);
  and (_01382_, _01140_, _01381_);
  not (_01383_, _33560_);
  and (_01384_, _01132_, _01383_);
  or (_01385_, _01384_, _01382_);
  or (_01386_, _01385_, _01380_);
  not (_01387_, _33724_);
  and (_01388_, _01088_, _01387_);
  not (_01389_, _33683_);
  and (_01390_, _01084_, _01389_);
  or (_01391_, _01390_, _01388_);
  not (_01392_, _33642_);
  and (_01393_, _01080_, _01392_);
  not (_01394_, _33765_);
  and (_01395_, _01147_, _01394_);
  not (_01396_, _33273_);
  and (_01397_, _01115_, _01396_);
  or (_01398_, _01397_, _01395_);
  not (_01399_, _33601_);
  and (_01400_, _01098_, _01399_);
  not (_01401_, _33437_);
  and (_01402_, _01095_, _01401_);
  or (_01403_, _01402_, _01400_);
  or (_01404_, _01403_, _01398_);
  or (_01405_, _01404_, _01393_);
  or (_01406_, _01405_, _01391_);
  not (_01407_, _33191_);
  and (_01408_, _01121_, _01407_);
  not (_01409_, _33396_);
  and (_01410_, _01104_, _01409_);
  not (_01411_, _33355_);
  and (_01412_, _01107_, _01411_);
  not (_01413_, _33314_);
  and (_01414_, _01111_, _01413_);
  or (_01415_, _01414_, _01412_);
  or (_01416_, _01415_, _01410_);
  or (_01417_, _01416_, _01408_);
  not (_01418_, _33519_);
  and (_01419_, _01135_, _01418_);
  not (_01420_, _33478_);
  and (_01421_, _01129_, _01420_);
  or (_01422_, _01421_, _01419_);
  or (_01423_, _01422_, _01417_);
  or (_01424_, _01423_, _01406_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _01424_, _01386_);
  not (_01425_, _33565_);
  and (_01426_, _01132_, _01425_);
  not (_01427_, _33483_);
  and (_01428_, _01129_, _01427_);
  not (_01429_, _33196_);
  and (_01430_, _01121_, _01429_);
  or (_01431_, _01430_, _01428_);
  or (_01432_, _01431_, _01426_);
  not (_01433_, _33688_);
  and (_01434_, _01084_, _01433_);
  not (_01435_, _33770_);
  and (_01436_, _01147_, _01435_);
  not (_01437_, _33442_);
  and (_01438_, _01095_, _01437_);
  or (_01439_, _01438_, _01436_);
  not (_01440_, _33606_);
  and (_01441_, _01098_, _01440_);
  not (_01442_, _33278_);
  and (_01443_, _01115_, _01442_);
  or (_01444_, _01443_, _01441_);
  or (_01445_, _01444_, _01439_);
  or (_01446_, _01445_, _01434_);
  not (_01447_, _33729_);
  and (_01448_, _01088_, _01447_);
  not (_01449_, _33647_);
  and (_01450_, _01080_, _01449_);
  or (_01451_, _01450_, _01448_);
  or (_01452_, _01451_, _01446_);
  not (_01453_, _33155_);
  and (_01454_, _01140_, _01453_);
  not (_01455_, _33237_);
  and (_01456_, _01143_, _01455_);
  or (_01457_, _01456_, _01454_);
  not (_01458_, _33524_);
  and (_01459_, _01135_, _01458_);
  not (_01460_, _33401_);
  and (_01461_, _01104_, _01460_);
  not (_01462_, _33360_);
  and (_01463_, _01107_, _01462_);
  not (_01464_, _33319_);
  and (_01465_, _01111_, _01464_);
  or (_01466_, _01465_, _01463_);
  or (_01467_, _01466_, _01461_);
  or (_01468_, _01467_, _01459_);
  or (_01469_, _01468_, _01457_);
  or (_01470_, _01469_, _01452_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _01470_, _01432_);
  not (_01471_, _33570_);
  and (_01472_, _01132_, _01471_);
  not (_01473_, _33488_);
  and (_01474_, _01129_, _01473_);
  not (_01475_, _33201_);
  and (_01476_, _01121_, _01475_);
  or (_01477_, _01476_, _01474_);
  or (_01478_, _01477_, _01472_);
  not (_01479_, _33693_);
  and (_01480_, _01084_, _01479_);
  not (_01481_, _33775_);
  and (_01482_, _01147_, _01481_);
  not (_01483_, _33447_);
  and (_01484_, _01095_, _01483_);
  or (_01485_, _01484_, _01482_);
  not (_01486_, _33611_);
  and (_01487_, _01098_, _01486_);
  not (_01488_, _33283_);
  and (_01489_, _01115_, _01488_);
  or (_01490_, _01489_, _01487_);
  or (_01491_, _01490_, _01485_);
  or (_01492_, _01491_, _01480_);
  not (_01493_, _33734_);
  and (_01494_, _01088_, _01493_);
  not (_01495_, _33652_);
  and (_01496_, _01080_, _01495_);
  or (_01497_, _01496_, _01494_);
  or (_01498_, _01497_, _01492_);
  not (_01499_, _33160_);
  and (_01500_, _01140_, _01499_);
  not (_01501_, _33242_);
  and (_01502_, _01143_, _01501_);
  or (_01503_, _01502_, _01500_);
  not (_01504_, _33529_);
  and (_01505_, _01135_, _01504_);
  not (_01506_, _33365_);
  and (_01507_, _01107_, _01506_);
  not (_01508_, _33406_);
  and (_01509_, _01104_, _01508_);
  or (_01510_, _01509_, _01507_);
  not (_01511_, _33324_);
  and (_01512_, _01111_, _01511_);
  or (_01513_, _01512_, _01510_);
  or (_01514_, _01513_, _01505_);
  or (_01515_, _01514_, _01503_);
  or (_01516_, _01515_, _01498_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _01516_, _01478_);
  not (_01517_, _33657_);
  and (_01518_, _01080_, _01517_);
  not (_01519_, _33698_);
  and (_01520_, _01084_, _01519_);
  not (_01521_, _33739_);
  and (_01522_, _01088_, _01521_);
  or (_01523_, _01522_, _01520_);
  or (_01524_, _01523_, _01518_);
  not (_01525_, _33452_);
  and (_01526_, _01095_, _01525_);
  not (_01527_, _33616_);
  and (_01528_, _01098_, _01527_);
  or (_01529_, _01528_, _01526_);
  or (_01530_, _01529_, _01524_);
  not (_01531_, _33288_);
  and (_01532_, _01115_, _01531_);
  not (_01533_, _33411_);
  and (_01534_, _01104_, _01533_);
  not (_01535_, _33370_);
  and (_01536_, _01107_, _01535_);
  or (_01537_, _01536_, _01534_);
  or (_01538_, _01537_, _01532_);
  not (_01539_, _33329_);
  and (_01540_, _01111_, _01539_);
  not (_01541_, _33206_);
  and (_01542_, _01121_, _01541_);
  or (_01543_, _01542_, _01540_);
  or (_01544_, _01543_, _01538_);
  or (_01545_, _01544_, _01530_);
  not (_01546_, _33493_);
  and (_01547_, _01129_, _01546_);
  not (_01548_, _33575_);
  and (_01549_, _01132_, _01548_);
  not (_01550_, _33534_);
  and (_01551_, _01135_, _01550_);
  or (_01552_, _01551_, _01549_);
  or (_01553_, _01552_, _01547_);
  not (_01554_, _33165_);
  and (_01555_, _01140_, _01554_);
  not (_01556_, _33247_);
  and (_01557_, _01143_, _01556_);
  or (_01558_, _01557_, _01555_);
  not (_01559_, _33780_);
  and (_01560_, _01147_, _01559_);
  or (_01561_, _01560_, _01558_);
  or (_01562_, _01561_, _01553_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _01562_, _01545_);
  and (_01563_, _01121_, _01251_);
  and (_01564_, _01140_, _01263_);
  and (_01565_, _01132_, _01243_);
  or (_01566_, _01565_, _01564_);
  or (_01567_, _01566_, _01563_);
  and (_01568_, _01088_, _01265_);
  and (_01569_, _01084_, _01256_);
  or (_01570_, _01569_, _01568_);
  and (_01571_, _01080_, _01241_);
  and (_01572_, _01147_, _01249_);
  and (_01573_, _01095_, _01278_);
  or (_01574_, _01573_, _01572_);
  and (_01575_, _01098_, _01274_);
  and (_01576_, _01115_, _01245_);
  or (_01577_, _01576_, _01575_);
  or (_01578_, _01577_, _01574_);
  or (_01579_, _01578_, _01571_);
  or (_01580_, _01579_, _01570_);
  and (_01581_, _01129_, _01276_);
  and (_01582_, _01107_, _01258_);
  and (_01583_, _01111_, _01271_);
  and (_01584_, _01104_, _01281_);
  or (_01585_, _01584_, _01583_);
  or (_01586_, _01585_, _01582_);
  or (_01587_, _01586_, _01581_);
  and (_01588_, _01135_, _01253_);
  and (_01589_, _01143_, _01269_);
  or (_01590_, _01589_, _01588_);
  or (_01591_, _01590_, _01587_);
  or (_01592_, _01591_, _01580_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _01592_, _01567_);
  and (_01593_, _01107_, _01308_);
  and (_01594_, _01104_, _01303_);
  or (_01595_, _01594_, _01593_);
  and (_01596_, _01129_, _01300_);
  and (_01597_, _01095_, _01298_);
  or (_01598_, _01597_, _01596_);
  or (_01599_, _01598_, _01595_);
  and (_01600_, _01140_, _01315_);
  and (_01601_, _01084_, _01318_);
  and (_01602_, _01088_, _01320_);
  or (_01603_, _01602_, _01601_);
  or (_01604_, _01603_, _01600_);
  and (_01605_, _01135_, _01292_);
  and (_01606_, _01121_, _01324_);
  or (_01607_, _01606_, _01605_);
  or (_01608_, _01607_, _01604_);
  or (_01609_, _01608_, _01599_);
  and (_01610_, _01143_, _01326_);
  and (_01611_, _01115_, _01306_);
  and (_01612_, _01111_, _01328_);
  or (_01613_, _01612_, _01611_);
  or (_01614_, _01613_, _01610_);
  and (_01615_, _01147_, _01313_);
  and (_01616_, _01132_, _01294_);
  and (_01617_, _01098_, _01289_);
  and (_01618_, _01080_, _01287_);
  or (_01619_, _01618_, _01617_);
  or (_01620_, _01619_, _01616_);
  or (_01621_, _01620_, _01615_);
  or (_01622_, _01621_, _01614_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _01622_, _01609_);
  and (_01623_, _01140_, _01341_);
  and (_01624_, _01084_, _01353_);
  and (_01625_, _01088_, _01346_);
  or (_01626_, _01625_, _01624_);
  or (_01627_, _01626_, _01623_);
  and (_01628_, _01132_, _01374_);
  and (_01629_, _01121_, _01348_);
  or (_01630_, _01629_, _01628_);
  or (_01631_, _01630_, _01627_);
  and (_01632_, _01095_, _01365_);
  and (_01633_, _01107_, _01355_);
  and (_01634_, _01104_, _01363_);
  or (_01635_, _01634_, _01633_);
  or (_01636_, _01635_, _01632_);
  and (_01637_, _01115_, _01335_);
  and (_01638_, _01129_, _01367_);
  or (_01639_, _01638_, _01637_);
  or (_01640_, _01639_, _01636_);
  or (_01641_, _01640_, _01631_);
  and (_01642_, _01147_, _01343_);
  and (_01643_, _01143_, _01361_);
  and (_01644_, _01111_, _01337_);
  or (_01645_, _01644_, _01643_);
  and (_01646_, _01135_, _01350_);
  and (_01647_, _01098_, _01333_);
  and (_01648_, _01080_, _01372_);
  or (_01649_, _01648_, _01647_);
  or (_01650_, _01649_, _01646_);
  or (_01651_, _01650_, _01645_);
  or (_01652_, _01651_, _01642_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _01652_, _01641_);
  and (_01653_, _01121_, _01394_);
  and (_01654_, _01132_, _01420_);
  or (_01655_, _01654_, _01653_);
  and (_01656_, _01140_, _01387_);
  and (_01657_, _01088_, _01392_);
  and (_01658_, _01084_, _01399_);
  or (_01659_, _01658_, _01657_);
  or (_01660_, _01659_, _01656_);
  or (_01661_, _01660_, _01655_);
  and (_01662_, _01095_, _01411_);
  and (_01663_, _01104_, _01413_);
  and (_01664_, _01107_, _01396_);
  or (_01665_, _01664_, _01663_);
  or (_01666_, _01665_, _01662_);
  and (_01667_, _01129_, _01409_);
  and (_01668_, _01115_, _01407_);
  or (_01669_, _01668_, _01667_);
  or (_01670_, _01669_, _01666_);
  or (_01671_, _01670_, _01661_);
  and (_01672_, _01147_, _01389_);
  and (_01673_, _01143_, _01381_);
  and (_01674_, _01111_, _01379_);
  or (_01675_, _01674_, _01673_);
  and (_01676_, _01135_, _01401_);
  and (_01677_, _01080_, _01383_);
  and (_01678_, _01098_, _01418_);
  or (_01679_, _01678_, _01677_);
  or (_01680_, _01679_, _01676_);
  or (_01681_, _01680_, _01675_);
  or (_01682_, _01681_, _01672_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _01682_, _01671_);
  and (_01683_, _01140_, _01447_);
  and (_01684_, _01084_, _01440_);
  and (_01685_, _01088_, _01449_);
  or (_01686_, _01685_, _01684_);
  or (_01687_, _01686_, _01683_);
  and (_01688_, _01132_, _01427_);
  and (_01689_, _01121_, _01435_);
  or (_01690_, _01689_, _01688_);
  or (_01691_, _01690_, _01687_);
  and (_01692_, _01095_, _01462_);
  and (_01693_, _01107_, _01442_);
  and (_01694_, _01104_, _01464_);
  or (_01695_, _01694_, _01693_);
  or (_01696_, _01695_, _01692_);
  and (_01697_, _01115_, _01429_);
  and (_01698_, _01129_, _01460_);
  or (_01699_, _01698_, _01697_);
  or (_01700_, _01699_, _01696_);
  or (_01701_, _01700_, _01691_);
  and (_01702_, _01147_, _01433_);
  and (_01703_, _01143_, _01453_);
  and (_01704_, _01111_, _01455_);
  or (_01705_, _01704_, _01703_);
  and (_01706_, _01135_, _01437_);
  and (_01707_, _01098_, _01458_);
  and (_01708_, _01080_, _01425_);
  or (_01709_, _01708_, _01707_);
  or (_01710_, _01709_, _01706_);
  or (_01711_, _01710_, _01705_);
  or (_01712_, _01711_, _01702_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _01712_, _01701_);
  and (_01713_, _01132_, _01473_);
  and (_01714_, _01135_, _01483_);
  and (_01715_, _01140_, _01493_);
  or (_01716_, _01715_, _01714_);
  or (_01717_, _01716_, _01713_);
  and (_01718_, _01088_, _01495_);
  and (_01719_, _01098_, _01504_);
  and (_01720_, _01095_, _01506_);
  or (_01721_, _01720_, _01719_);
  and (_01722_, _01147_, _01479_);
  and (_01723_, _01115_, _01475_);
  or (_01724_, _01723_, _01722_);
  or (_01725_, _01724_, _01721_);
  or (_01726_, _01725_, _01718_);
  and (_01727_, _01080_, _01471_);
  and (_01728_, _01084_, _01486_);
  or (_01729_, _01728_, _01727_);
  or (_01730_, _01729_, _01726_);
  and (_01731_, _01129_, _01508_);
  and (_01732_, _01107_, _01488_);
  and (_01733_, _01111_, _01501_);
  and (_01734_, _01104_, _01511_);
  or (_01735_, _01734_, _01733_);
  or (_01736_, _01735_, _01732_);
  or (_01737_, _01736_, _01731_);
  and (_01738_, _01121_, _01481_);
  and (_01739_, _01143_, _01499_);
  or (_01740_, _01739_, _01738_);
  or (_01741_, _01740_, _01737_);
  or (_01742_, _01741_, _01730_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _01742_, _01717_);
  and (_01743_, _01098_, _01550_);
  and (_01744_, _01080_, _01548_);
  or (_01745_, _01744_, _01743_);
  and (_01746_, _01135_, _01525_);
  and (_01747_, _01132_, _01546_);
  or (_01748_, _01747_, _01746_);
  or (_01749_, _01748_, _01745_);
  and (_01750_, _01095_, _01535_);
  and (_01751_, _01107_, _01531_);
  and (_01752_, _01104_, _01539_);
  or (_01753_, _01752_, _01751_);
  or (_01754_, _01753_, _01750_);
  and (_01755_, _01129_, _01533_);
  and (_01756_, _01115_, _01541_);
  or (_01757_, _01756_, _01755_);
  or (_01758_, _01757_, _01754_);
  or (_01759_, _01758_, _01749_);
  and (_01760_, _01121_, _01559_);
  and (_01761_, _01140_, _01521_);
  and (_01762_, _01084_, _01527_);
  and (_01763_, _01088_, _01517_);
  or (_01764_, _01763_, _01762_);
  or (_01765_, _01764_, _01761_);
  or (_01766_, _01765_, _01760_);
  and (_01767_, _01147_, _01519_);
  and (_01768_, _01143_, _01554_);
  and (_01769_, _01111_, _01556_);
  or (_01770_, _01769_, _01768_);
  or (_01771_, _01770_, _01767_);
  or (_01772_, _01771_, _01766_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _01772_, _01759_);
  and (_01773_, _01132_, _01274_);
  and (_01774_, _01129_, _01253_);
  and (_01775_, _01143_, _01245_);
  or (_01776_, _01775_, _01774_);
  or (_01777_, _01776_, _01773_);
  and (_01778_, _01080_, _01256_);
  and (_01779_, _01147_, _01263_);
  and (_01780_, _01095_, _01276_);
  or (_01781_, _01780_, _01779_);
  and (_01782_, _01098_, _01241_);
  and (_01783_, _01115_, _01271_);
  or (_01784_, _01783_, _01782_);
  or (_01785_, _01784_, _01781_);
  or (_01786_, _01785_, _01778_);
  and (_01787_, _01084_, _01265_);
  and (_01788_, _01088_, _01249_);
  or (_01789_, _01788_, _01787_);
  or (_01790_, _01789_, _01786_);
  and (_01791_, _01135_, _01243_);
  and (_01792_, _01111_, _01258_);
  and (_01793_, _01104_, _01278_);
  and (_01794_, _01107_, _01281_);
  or (_01795_, _01794_, _01793_);
  or (_01796_, _01795_, _01792_);
  or (_01797_, _01796_, _01791_);
  and (_01798_, _01140_, _01251_);
  and (_01799_, _01121_, _01269_);
  or (_01800_, _01799_, _01798_);
  or (_01801_, _01800_, _01797_);
  or (_01802_, _01801_, _01790_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _01802_, _01777_);
  and (_01803_, _01140_, _01324_);
  and (_01804_, _01129_, _01292_);
  and (_01805_, _01121_, _01326_);
  or (_01806_, _01805_, _01804_);
  or (_01807_, _01806_, _01803_);
  and (_01808_, _01084_, _01320_);
  and (_01809_, _01080_, _01318_);
  or (_01810_, _01809_, _01808_);
  and (_01811_, _01088_, _01313_);
  and (_01812_, _01095_, _01300_);
  and (_01813_, _01115_, _01328_);
  or (_01814_, _01813_, _01812_);
  and (_01815_, _01147_, _01315_);
  and (_01816_, _01098_, _01287_);
  or (_01817_, _01816_, _01815_);
  or (_01818_, _01817_, _01814_);
  or (_01819_, _01818_, _01811_);
  or (_01820_, _01819_, _01810_);
  and (_01821_, _01143_, _01306_);
  and (_01822_, _01111_, _01308_);
  and (_01823_, _01104_, _01298_);
  and (_01824_, _01107_, _01303_);
  or (_01825_, _01824_, _01823_);
  or (_01826_, _01825_, _01822_);
  or (_01827_, _01826_, _01821_);
  and (_01828_, _01132_, _01289_);
  and (_01829_, _01135_, _01294_);
  or (_01830_, _01829_, _01828_);
  or (_01831_, _01830_, _01827_);
  or (_01832_, _01831_, _01820_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _01832_, _01807_);
  and (_01833_, _01143_, _01335_);
  and (_01834_, _01121_, _01361_);
  and (_01835_, _01132_, _01333_);
  or (_01836_, _01835_, _01834_);
  or (_01837_, _01836_, _01833_);
  and (_01838_, _01084_, _01346_);
  and (_01839_, _01115_, _01337_);
  and (_01840_, _01147_, _01341_);
  or (_01841_, _01840_, _01839_);
  and (_01842_, _01095_, _01367_);
  and (_01843_, _01098_, _01372_);
  or (_01844_, _01843_, _01842_);
  or (_01845_, _01844_, _01841_);
  or (_01846_, _01845_, _01838_);
  and (_01847_, _01080_, _01353_);
  and (_01848_, _01088_, _01343_);
  or (_01849_, _01848_, _01847_);
  or (_01850_, _01849_, _01846_);
  and (_01851_, _01129_, _01350_);
  and (_01852_, _01135_, _01374_);
  or (_01853_, _01852_, _01851_);
  and (_01854_, _01140_, _01348_);
  and (_01855_, _01111_, _01355_);
  and (_01856_, _01104_, _01365_);
  and (_01857_, _01107_, _01363_);
  or (_01858_, _01857_, _01856_);
  or (_01859_, _01858_, _01855_);
  or (_01860_, _01859_, _01854_);
  or (_01861_, _01860_, _01853_);
  or (_01862_, _01861_, _01850_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _01862_, _01837_);
  and (_01863_, _01140_, _01394_);
  and (_01864_, _01135_, _01420_);
  and (_01865_, _01121_, _01381_);
  or (_01866_, _01865_, _01864_);
  or (_01867_, _01866_, _01863_);
  and (_01868_, _01084_, _01392_);
  and (_01869_, _01080_, _01399_);
  or (_01870_, _01869_, _01868_);
  and (_01871_, _01088_, _01389_);
  and (_01872_, _01095_, _01409_);
  and (_01873_, _01115_, _01379_);
  or (_01874_, _01873_, _01872_);
  and (_01875_, _01147_, _01387_);
  and (_01876_, _01098_, _01383_);
  or (_01877_, _01876_, _01875_);
  or (_01878_, _01877_, _01874_);
  or (_01879_, _01878_, _01871_);
  or (_01880_, _01879_, _01870_);
  and (_01881_, _01143_, _01407_);
  and (_01882_, _01107_, _01413_);
  and (_01883_, _01104_, _01411_);
  and (_01884_, _01111_, _01396_);
  or (_01885_, _01884_, _01883_);
  or (_01886_, _01885_, _01882_);
  or (_01887_, _01886_, _01881_);
  and (_01888_, _01132_, _01418_);
  and (_01889_, _01129_, _01401_);
  or (_01890_, _01889_, _01888_);
  or (_01891_, _01890_, _01887_);
  or (_01892_, _01891_, _01880_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _01892_, _01867_);
  and (_01893_, _01135_, _01427_);
  and (_01894_, _01140_, _01435_);
  and (_01895_, _01129_, _01437_);
  or (_01896_, _01895_, _01894_);
  or (_01897_, _01896_, _01893_);
  and (_01898_, _01084_, _01449_);
  and (_01899_, _01080_, _01440_);
  or (_01900_, _01899_, _01898_);
  and (_01901_, _01088_, _01433_);
  and (_01902_, _01098_, _01425_);
  and (_01903_, _01095_, _01460_);
  or (_01904_, _01903_, _01902_);
  and (_01905_, _01147_, _01447_);
  and (_01906_, _01115_, _01455_);
  or (_01907_, _01906_, _01905_);
  or (_01908_, _01907_, _01904_);
  or (_01909_, _01908_, _01901_);
  or (_01910_, _01909_, _01900_);
  and (_01911_, _01143_, _01429_);
  and (_01912_, _01107_, _01464_);
  and (_01913_, _01104_, _01462_);
  and (_01914_, _01111_, _01442_);
  or (_01915_, _01914_, _01913_);
  or (_01916_, _01915_, _01912_);
  or (_01917_, _01916_, _01911_);
  and (_01918_, _01132_, _01458_);
  and (_01919_, _01121_, _01453_);
  or (_01920_, _01919_, _01918_);
  or (_01921_, _01920_, _01917_);
  or (_01922_, _01921_, _01910_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _01922_, _01897_);
  and (_01923_, _01098_, _01471_);
  and (_01924_, _01132_, _01504_);
  or (_01925_, _01924_, _01923_);
  and (_01926_, _01135_, _01473_);
  and (_01927_, _01129_, _01483_);
  or (_01928_, _01927_, _01926_);
  or (_01929_, _01928_, _01925_);
  and (_01930_, _01140_, _01481_);
  and (_01931_, _01088_, _01479_);
  and (_01932_, _01080_, _01486_);
  and (_01933_, _01084_, _01495_);
  or (_01934_, _01933_, _01932_);
  or (_01935_, _01934_, _01931_);
  or (_01936_, _01935_, _01930_);
  or (_01937_, _01936_, _01929_);
  and (_01938_, _01143_, _01475_);
  and (_01939_, _01107_, _01511_);
  and (_01940_, _01111_, _01488_);
  or (_01941_, _01940_, _01939_);
  and (_01942_, _01095_, _01508_);
  and (_01943_, _01104_, _01506_);
  or (_01944_, _01943_, _01942_);
  or (_01945_, _01944_, _01941_);
  or (_01946_, _01945_, _01938_);
  and (_01947_, _01147_, _01493_);
  and (_01948_, _01121_, _01499_);
  and (_01949_, _01115_, _01501_);
  or (_01950_, _01949_, _01948_);
  or (_01951_, _01950_, _01947_);
  or (_01952_, _01951_, _01946_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _01952_, _01937_);
  and (_01953_, _01135_, _01546_);
  and (_01954_, _01129_, _01525_);
  and (_01955_, _01121_, _01554_);
  or (_01956_, _01955_, _01954_);
  or (_01957_, _01956_, _01953_);
  and (_01958_, _01084_, _01517_);
  and (_01959_, _01080_, _01527_);
  or (_01960_, _01959_, _01958_);
  and (_01961_, _01088_, _01519_);
  and (_01962_, _01098_, _01548_);
  and (_01963_, _01115_, _01556_);
  or (_01964_, _01963_, _01962_);
  and (_01965_, _01147_, _01521_);
  and (_01966_, _01095_, _01533_);
  or (_01967_, _01966_, _01965_);
  or (_01968_, _01967_, _01964_);
  or (_01969_, _01968_, _01961_);
  or (_01970_, _01969_, _01960_);
  and (_01971_, _01132_, _01550_);
  and (_01972_, _01107_, _01539_);
  and (_01973_, _01111_, _01531_);
  or (_01974_, _01973_, _01972_);
  and (_01975_, _01104_, _01535_);
  or (_01976_, _01975_, _01974_);
  or (_01977_, _01976_, _01971_);
  and (_01978_, _01140_, _01559_);
  and (_01979_, _01143_, _01541_);
  or (_01980_, _01979_, _01978_);
  or (_01981_, _01980_, _01977_);
  or (_01982_, _01981_, _01970_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _01982_, _01957_);
  and (_01983_, _01121_, _01263_);
  and (_01984_, _01132_, _01253_);
  and (_01985_, _01129_, _01278_);
  or (_01986_, _01985_, _01984_);
  or (_01987_, _01986_, _01983_);
  and (_01988_, _01080_, _01274_);
  and (_01989_, _01115_, _01269_);
  and (_01990_, _01095_, _01281_);
  or (_01991_, _01990_, _01989_);
  and (_01992_, _01147_, _01265_);
  and (_01993_, _01098_, _01243_);
  or (_01994_, _01993_, _01992_);
  or (_01995_, _01994_, _01991_);
  or (_01996_, _01995_, _01988_);
  and (_01997_, _01088_, _01256_);
  and (_01998_, _01084_, _01241_);
  or (_01999_, _01998_, _01997_);
  or (_02000_, _01999_, _01996_);
  and (_02001_, _01135_, _01276_);
  and (_02002_, _01111_, _01245_);
  and (_02003_, _01107_, _01271_);
  and (_02004_, _01104_, _01258_);
  or (_02005_, _02004_, _02003_);
  or (_02006_, _02005_, _02002_);
  or (_02007_, _02006_, _02001_);
  and (_02008_, _01143_, _01251_);
  and (_02009_, _01140_, _01249_);
  or (_02010_, _02009_, _02008_);
  or (_02011_, _02010_, _02007_);
  or (_02012_, _02011_, _02000_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _02012_, _01987_);
  and (_02013_, _01129_, _01298_);
  and (_02014_, _01143_, _01324_);
  and (_02015_, _01135_, _01300_);
  or (_02016_, _02015_, _02014_);
  or (_02017_, _02016_, _02013_);
  and (_02018_, _01084_, _01287_);
  and (_02019_, _01080_, _01289_);
  or (_02020_, _02019_, _02018_);
  and (_02021_, _01088_, _01318_);
  and (_02022_, _01095_, _01303_);
  and (_02023_, _01147_, _01320_);
  or (_02024_, _02023_, _02022_);
  and (_02025_, _01115_, _01326_);
  and (_02026_, _01098_, _01294_);
  or (_02027_, _02026_, _02025_);
  or (_02028_, _02027_, _02024_);
  or (_02029_, _02028_, _02021_);
  or (_02030_, _02029_, _02020_);
  and (_02031_, _01140_, _01313_);
  and (_02032_, _01111_, _01306_);
  and (_02033_, _01107_, _01328_);
  and (_02034_, _01104_, _01308_);
  or (_02035_, _02034_, _02033_);
  or (_02036_, _02035_, _02032_);
  or (_02037_, _02036_, _02031_);
  and (_02038_, _01132_, _01292_);
  and (_02039_, _01121_, _01315_);
  or (_02040_, _02039_, _02038_);
  or (_02041_, _02040_, _02037_);
  or (_02042_, _02041_, _02030_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _02042_, _02017_);
  and (_02043_, _01121_, _01341_);
  and (_02044_, _01132_, _01350_);
  and (_02045_, _01140_, _01343_);
  or (_02046_, _02045_, _02044_);
  or (_02047_, _02046_, _02043_);
  and (_02048_, _01080_, _01333_);
  and (_02049_, _01115_, _01361_);
  and (_02050_, _01147_, _01346_);
  or (_02051_, _02050_, _02049_);
  and (_02052_, _01095_, _01363_);
  and (_02053_, _01098_, _01374_);
  or (_02054_, _02053_, _02052_);
  or (_02055_, _02054_, _02051_);
  or (_02056_, _02055_, _02048_);
  and (_02057_, _01084_, _01372_);
  and (_02058_, _01088_, _01353_);
  or (_02059_, _02058_, _02057_);
  or (_02060_, _02059_, _02056_);
  and (_02061_, _01135_, _01367_);
  and (_02062_, _01107_, _01337_);
  and (_02063_, _01111_, _01335_);
  or (_02064_, _02063_, _02062_);
  and (_02065_, _01104_, _01355_);
  or (_02066_, _02065_, _02064_);
  or (_02067_, _02066_, _02061_);
  and (_02068_, _01143_, _01348_);
  and (_02069_, _01129_, _01365_);
  or (_02070_, _02069_, _02068_);
  or (_02071_, _02070_, _02067_);
  or (_02072_, _02071_, _02060_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _02072_, _02047_);
  and (_02073_, _01135_, _01409_);
  and (_02074_, _01129_, _01411_);
  or (_02075_, _02074_, _02073_);
  and (_02076_, _01140_, _01389_);
  or (_02077_, _02076_, _02075_);
  and (_02078_, _01080_, _01418_);
  and (_02079_, _01115_, _01381_);
  and (_02080_, _01095_, _01413_);
  or (_02081_, _02080_, _02079_);
  and (_02082_, _01098_, _01420_);
  and (_02083_, _01147_, _01392_);
  or (_02084_, _02083_, _02082_);
  or (_02085_, _02084_, _02081_);
  or (_02086_, _02085_, _02078_);
  and (_02087_, _01084_, _01383_);
  and (_02088_, _01088_, _01399_);
  or (_02089_, _02088_, _02087_);
  or (_02090_, _02089_, _02086_);
  and (_02091_, _01143_, _01394_);
  and (_02092_, _01121_, _01387_);
  or (_02093_, _02092_, _02091_);
  and (_02094_, _01132_, _01401_);
  and (_02095_, _01111_, _01407_);
  and (_02096_, _01107_, _01379_);
  and (_02097_, _01104_, _01396_);
  or (_02098_, _02097_, _02096_);
  or (_02099_, _02098_, _02095_);
  or (_02100_, _02099_, _02094_);
  or (_02101_, _02100_, _02093_);
  or (_02102_, _02101_, _02090_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _02102_, _02077_);
  and (_02103_, _01135_, _01460_);
  and (_02104_, _01129_, _01462_);
  or (_02105_, _02104_, _02103_);
  and (_02106_, _01140_, _01433_);
  or (_02107_, _02106_, _02105_);
  and (_02108_, _01080_, _01458_);
  and (_02109_, _01115_, _01453_);
  and (_02110_, _01095_, _01464_);
  or (_02111_, _02110_, _02109_);
  and (_02112_, _01098_, _01427_);
  and (_02113_, _01147_, _01449_);
  or (_02114_, _02113_, _02112_);
  or (_02115_, _02114_, _02111_);
  or (_02116_, _02115_, _02108_);
  and (_02117_, _01084_, _01425_);
  and (_02118_, _01088_, _01440_);
  or (_02119_, _02118_, _02117_);
  or (_02120_, _02119_, _02116_);
  and (_02121_, _01143_, _01435_);
  and (_02122_, _01121_, _01447_);
  or (_02123_, _02122_, _02121_);
  and (_02124_, _01132_, _01437_);
  and (_02125_, _01111_, _01429_);
  and (_02126_, _01107_, _01455_);
  and (_02127_, _01104_, _01442_);
  or (_02128_, _02127_, _02126_);
  or (_02129_, _02128_, _02125_);
  or (_02130_, _02129_, _02124_);
  or (_02131_, _02130_, _02123_);
  or (_02132_, _02131_, _02120_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _02132_, _02107_);
  and (_02133_, _01132_, _01483_);
  and (_02134_, _01143_, _01481_);
  and (_02135_, _01129_, _01506_);
  or (_02136_, _02135_, _02134_);
  or (_02137_, _02136_, _02133_);
  and (_02138_, _01084_, _01471_);
  and (_02139_, _01080_, _01504_);
  or (_02140_, _02139_, _02138_);
  and (_02141_, _01088_, _01486_);
  and (_02142_, _01098_, _01473_);
  and (_02143_, _01147_, _01495_);
  or (_02144_, _02143_, _02142_);
  and (_02145_, _01115_, _01499_);
  and (_02146_, _01095_, _01511_);
  or (_02147_, _02146_, _02145_);
  or (_02148_, _02147_, _02144_);
  or (_02149_, _02148_, _02141_);
  or (_02150_, _02149_, _02140_);
  and (_02151_, _01121_, _01493_);
  and (_02152_, _01140_, _01479_);
  or (_02153_, _02152_, _02151_);
  and (_02154_, _01135_, _01508_);
  and (_02155_, _01111_, _01475_);
  and (_02156_, _01107_, _01501_);
  or (_02157_, _02156_, _02155_);
  and (_02158_, _01104_, _01488_);
  or (_02159_, _02158_, _02157_);
  or (_02160_, _02159_, _02154_);
  or (_02161_, _02160_, _02153_);
  or (_02162_, _02161_, _02150_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _02162_, _02137_);
  and (_02163_, _01135_, _01533_);
  and (_02164_, _01129_, _01535_);
  and (_02165_, _01140_, _01519_);
  or (_02166_, _02165_, _02164_);
  or (_02167_, _02166_, _02163_);
  and (_02168_, _01084_, _01548_);
  and (_02169_, _01080_, _01550_);
  or (_02170_, _02169_, _02168_);
  and (_02171_, _01088_, _01527_);
  and (_02172_, _01115_, _01554_);
  and (_02173_, _01147_, _01517_);
  or (_02174_, _02173_, _02172_);
  and (_02175_, _01095_, _01539_);
  and (_02176_, _01098_, _01546_);
  or (_02177_, _02176_, _02175_);
  or (_02178_, _02177_, _02174_);
  or (_02179_, _02178_, _02171_);
  or (_02180_, _02179_, _02170_);
  and (_02181_, _01121_, _01521_);
  and (_02182_, _01111_, _01541_);
  and (_02183_, _01107_, _01556_);
  or (_02184_, _02183_, _02182_);
  and (_02185_, _01104_, _01531_);
  or (_02186_, _02185_, _02184_);
  or (_02187_, _02186_, _02181_);
  and (_02188_, _01143_, _01559_);
  and (_02189_, _01132_, _01525_);
  or (_02190_, _02189_, _02188_);
  or (_02191_, _02190_, _02187_);
  or (_02192_, _02191_, _02180_);
  or (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _02192_, _02167_);
  nand (_02193_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not (_02194_, \oc8051_golden_model_1.PC [3]);
  or (_02195_, \oc8051_golden_model_1.PC [2], _02194_);
  or (_02196_, _02195_, _02193_);
  or (_02197_, _02196_, _33616_);
  not (_02198_, \oc8051_golden_model_1.PC [1]);
  or (_02199_, _02198_, \oc8051_golden_model_1.PC [0]);
  or (_02200_, _02199_, _02195_);
  or (_02201_, _02200_, _33575_);
  and (_02202_, _02201_, _02197_);
  not (_02203_, \oc8051_golden_model_1.PC [2]);
  or (_02204_, _02203_, \oc8051_golden_model_1.PC [3]);
  or (_02205_, _02204_, _02193_);
  or (_02206_, _02205_, _33452_);
  or (_02207_, _02204_, _02199_);
  or (_02208_, _02207_, _33411_);
  and (_02209_, _02208_, _02206_);
  and (_02210_, _02209_, _02202_);
  nand (_02211_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02212_, _02211_, _02193_);
  or (_02213_, _02212_, _33780_);
  or (_02214_, _02211_, _02199_);
  or (_02215_, _02214_, _33739_);
  and (_02216_, _02215_, _02213_);
  or (_02217_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or (_02218_, _02217_, _02193_);
  or (_02219_, _02218_, _33288_);
  or (_02220_, _02217_, _02199_);
  or (_02221_, _02220_, _33247_);
  and (_02222_, _02221_, _02219_);
  and (_02223_, _02222_, _02216_);
  and (_02224_, _02223_, _02210_);
  not (_02225_, \oc8051_golden_model_1.PC [0]);
  or (_02226_, \oc8051_golden_model_1.PC [1], _02225_);
  or (_02227_, _02226_, _02211_);
  or (_02228_, _02227_, _33698_);
  or (_02229_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or (_02230_, _02229_, _02211_);
  or (_02231_, _02230_, _33657_);
  and (_02232_, _02231_, _02228_);
  or (_02233_, _02217_, _02229_);
  or (_02234_, _02233_, _33165_);
  or (_02235_, _02217_, _02226_);
  or (_02236_, _02235_, _33206_);
  and (_02237_, _02236_, _02234_);
  and (_02238_, _02237_, _02232_);
  or (_02239_, _02226_, _02195_);
  or (_02240_, _02239_, _33534_);
  or (_02241_, _02229_, _02195_);
  or (_02242_, _02241_, _33493_);
  and (_02243_, _02242_, _02240_);
  or (_02244_, _02226_, _02204_);
  or (_02245_, _02244_, _33370_);
  or (_02246_, _02229_, _02204_);
  or (_02247_, _02246_, _33329_);
  and (_02248_, _02247_, _02245_);
  and (_02249_, _02248_, _02243_);
  and (_02250_, _02249_, _02238_);
  nand (_02251_, _02250_, _02224_);
  or (_02252_, _02196_, _33581_);
  or (_02253_, _02200_, _33540_);
  and (_02254_, _02253_, _02252_);
  or (_02255_, _02205_, _33417_);
  or (_02256_, _02207_, _33376_);
  and (_02257_, _02256_, _02255_);
  and (_02258_, _02257_, _02254_);
  or (_02259_, _02212_, _33745_);
  or (_02260_, _02214_, _33704_);
  and (_02261_, _02260_, _02259_);
  or (_02262_, _02218_, _33253_);
  or (_02263_, _02220_, _33212_);
  and (_02264_, _02263_, _02262_);
  and (_02265_, _02264_, _02261_);
  and (_02266_, _02265_, _02258_);
  or (_02267_, _02227_, _33663_);
  or (_02268_, _02230_, _33622_);
  and (_02269_, _02268_, _02267_);
  or (_02270_, _02233_, _33130_);
  or (_02271_, _02235_, _33171_);
  and (_02272_, _02271_, _02270_);
  and (_02273_, _02272_, _02269_);
  or (_02274_, _02239_, _33499_);
  or (_02275_, _02241_, _33458_);
  and (_02276_, _02275_, _02274_);
  or (_02277_, _02244_, _33335_);
  or (_02278_, _02246_, _33294_);
  and (_02279_, _02278_, _02277_);
  and (_02280_, _02279_, _02276_);
  and (_02281_, _02280_, _02273_);
  and (_02282_, _02281_, _02266_);
  or (_02283_, _02282_, _02251_);
  or (_02284_, _02196_, _33606_);
  or (_02285_, _02200_, _33565_);
  and (_02286_, _02285_, _02284_);
  or (_02287_, _02205_, _33442_);
  or (_02288_, _02207_, _33401_);
  and (_02289_, _02288_, _02287_);
  and (_02290_, _02289_, _02286_);
  or (_02291_, _02212_, _33770_);
  or (_02292_, _02214_, _33729_);
  and (_02293_, _02292_, _02291_);
  or (_02294_, _02218_, _33278_);
  or (_02295_, _02220_, _33237_);
  and (_02296_, _02295_, _02294_);
  and (_02297_, _02296_, _02293_);
  and (_02298_, _02297_, _02290_);
  or (_02299_, _02227_, _33688_);
  or (_02300_, _02230_, _33647_);
  and (_02301_, _02300_, _02299_);
  or (_02302_, _02233_, _33155_);
  or (_02303_, _02235_, _33196_);
  and (_02304_, _02303_, _02302_);
  and (_02305_, _02304_, _02301_);
  or (_02306_, _02239_, _33524_);
  or (_02307_, _02241_, _33483_);
  and (_02308_, _02307_, _02306_);
  or (_02309_, _02244_, _33360_);
  or (_02310_, _02246_, _33319_);
  and (_02311_, _02310_, _02309_);
  and (_02312_, _02311_, _02308_);
  and (_02313_, _02312_, _02305_);
  nand (_02314_, _02313_, _02298_);
  or (_02315_, _02196_, _33611_);
  or (_02316_, _02200_, _33570_);
  and (_02317_, _02316_, _02315_);
  or (_02318_, _02205_, _33447_);
  or (_02319_, _02207_, _33406_);
  and (_02320_, _02319_, _02318_);
  and (_02321_, _02320_, _02317_);
  or (_02322_, _02212_, _33775_);
  or (_02323_, _02214_, _33734_);
  and (_02324_, _02323_, _02322_);
  or (_02325_, _02218_, _33283_);
  or (_02326_, _02220_, _33242_);
  and (_02327_, _02326_, _02325_);
  and (_02328_, _02327_, _02324_);
  and (_02329_, _02328_, _02321_);
  or (_02330_, _02227_, _33693_);
  or (_02331_, _02230_, _33652_);
  and (_02332_, _02331_, _02330_);
  or (_02333_, _02233_, _33160_);
  or (_02334_, _02235_, _33201_);
  and (_02335_, _02334_, _02333_);
  and (_02336_, _02335_, _02332_);
  or (_02337_, _02239_, _33529_);
  or (_02338_, _02241_, _33488_);
  and (_02339_, _02338_, _02337_);
  or (_02340_, _02244_, _33365_);
  or (_02341_, _02246_, _33324_);
  and (_02342_, _02341_, _02340_);
  and (_02343_, _02342_, _02339_);
  and (_02344_, _02343_, _02336_);
  nand (_02345_, _02344_, _02329_);
  or (_02346_, _02345_, _02314_);
  nor (_02347_, _02346_, _02283_);
  or (_02348_, _02196_, _33596_);
  or (_02349_, _02200_, _33555_);
  and (_02350_, _02349_, _02348_);
  or (_02351_, _02205_, _33432_);
  or (_02352_, _02207_, _33391_);
  and (_02353_, _02352_, _02351_);
  and (_02354_, _02353_, _02350_);
  or (_02355_, _02212_, _33760_);
  or (_02356_, _02214_, _33719_);
  and (_02357_, _02356_, _02355_);
  or (_02358_, _02218_, _33268_);
  or (_02359_, _02220_, _33227_);
  and (_02360_, _02359_, _02358_);
  and (_02361_, _02360_, _02357_);
  and (_02362_, _02361_, _02354_);
  or (_02363_, _02227_, _33678_);
  or (_02364_, _02230_, _33637_);
  and (_02365_, _02364_, _02363_);
  or (_02366_, _02233_, _33145_);
  or (_02367_, _02235_, _33186_);
  and (_02368_, _02367_, _02366_);
  and (_02369_, _02368_, _02365_);
  or (_02370_, _02239_, _33514_);
  or (_02371_, _02241_, _33473_);
  and (_02372_, _02371_, _02370_);
  or (_02373_, _02244_, _33350_);
  or (_02374_, _02246_, _33309_);
  and (_02375_, _02374_, _02373_);
  and (_02376_, _02375_, _02372_);
  and (_02377_, _02376_, _02369_);
  nand (_02378_, _02377_, _02362_);
  or (_02379_, _02196_, _33601_);
  or (_02380_, _02200_, _33560_);
  and (_02381_, _02380_, _02379_);
  or (_02382_, _02205_, _33437_);
  or (_02383_, _02207_, _33396_);
  and (_02384_, _02383_, _02382_);
  and (_02385_, _02384_, _02381_);
  or (_02386_, _02212_, _33765_);
  or (_02387_, _02214_, _33724_);
  and (_02388_, _02387_, _02386_);
  or (_02389_, _02218_, _33273_);
  or (_02390_, _02220_, _33232_);
  and (_02391_, _02390_, _02389_);
  and (_02392_, _02391_, _02388_);
  and (_02393_, _02392_, _02385_);
  or (_02394_, _02227_, _33683_);
  or (_02395_, _02230_, _33642_);
  and (_02396_, _02395_, _02394_);
  or (_02397_, _02233_, _33150_);
  or (_02398_, _02235_, _33191_);
  and (_02399_, _02398_, _02397_);
  and (_02400_, _02399_, _02396_);
  or (_02401_, _02239_, _33519_);
  or (_02402_, _02241_, _33478_);
  and (_02403_, _02402_, _02401_);
  or (_02404_, _02244_, _33355_);
  or (_02405_, _02246_, _33314_);
  and (_02406_, _02405_, _02404_);
  and (_02407_, _02406_, _02403_);
  and (_02408_, _02407_, _02400_);
  nand (_02409_, _02408_, _02393_);
  or (_02410_, _02409_, _02378_);
  or (_02411_, _02196_, _33586_);
  or (_02412_, _02200_, _33545_);
  and (_02413_, _02412_, _02411_);
  or (_02414_, _02205_, _33422_);
  or (_02415_, _02207_, _33381_);
  and (_02416_, _02415_, _02414_);
  and (_02417_, _02416_, _02413_);
  or (_02418_, _02212_, _33750_);
  or (_02419_, _02214_, _33709_);
  and (_02420_, _02419_, _02418_);
  or (_02421_, _02218_, _33258_);
  or (_02422_, _02220_, _33217_);
  and (_02423_, _02422_, _02421_);
  and (_02424_, _02423_, _02420_);
  and (_02425_, _02424_, _02417_);
  or (_02426_, _02227_, _33668_);
  or (_02427_, _02230_, _33627_);
  and (_02428_, _02427_, _02426_);
  or (_02429_, _02233_, _33135_);
  or (_02430_, _02235_, _33176_);
  and (_02431_, _02430_, _02429_);
  and (_02432_, _02431_, _02428_);
  or (_02433_, _02239_, _33504_);
  or (_02434_, _02241_, _33463_);
  and (_02435_, _02434_, _02433_);
  or (_02436_, _02244_, _33340_);
  or (_02437_, _02246_, _33299_);
  and (_02438_, _02437_, _02436_);
  and (_02439_, _02438_, _02435_);
  and (_02440_, _02439_, _02432_);
  and (_02441_, _02440_, _02425_);
  or (_02442_, _02196_, _33591_);
  or (_02443_, _02200_, _33550_);
  and (_02444_, _02443_, _02442_);
  or (_02445_, _02205_, _33427_);
  or (_02446_, _02207_, _33386_);
  and (_02447_, _02446_, _02445_);
  and (_02448_, _02447_, _02444_);
  or (_02449_, _02212_, _33755_);
  or (_02450_, _02214_, _33714_);
  and (_02451_, _02450_, _02449_);
  or (_02452_, _02218_, _33263_);
  or (_02453_, _02220_, _33222_);
  and (_02454_, _02453_, _02452_);
  and (_02455_, _02454_, _02451_);
  and (_02456_, _02455_, _02448_);
  or (_02457_, _02227_, _33673_);
  or (_02458_, _02230_, _33632_);
  and (_02459_, _02458_, _02457_);
  or (_02460_, _02233_, _33140_);
  or (_02461_, _02235_, _33181_);
  and (_02462_, _02461_, _02460_);
  and (_02463_, _02462_, _02459_);
  or (_02464_, _02239_, _33509_);
  or (_02465_, _02241_, _33468_);
  and (_02466_, _02465_, _02464_);
  or (_02467_, _02244_, _33345_);
  or (_02468_, _02246_, _33304_);
  and (_02469_, _02468_, _02467_);
  and (_02470_, _02469_, _02466_);
  and (_02471_, _02470_, _02463_);
  and (_02472_, _02471_, _02456_);
  or (_02473_, _02472_, _02441_);
  or (_02474_, _02473_, _02410_);
  not (_02475_, _02474_);
  and (_02476_, _02475_, _02347_);
  not (_02477_, \oc8051_golden_model_1.ACC [1]);
  and (_02478_, _02226_, _02199_);
  nor (_02479_, _02478_, _02477_);
  and (_02480_, \oc8051_golden_model_1.ACC [0], _02225_);
  and (_02481_, _02478_, _02477_);
  nor (_02482_, _02481_, _02479_);
  and (_02483_, _02482_, _02480_);
  nor (_02484_, _02483_, _02479_);
  nor (_02485_, _02193_, _02203_);
  and (_02486_, _02193_, _02203_);
  nor (_02487_, _02486_, _02485_);
  and (_02488_, _02487_, \oc8051_golden_model_1.ACC [2]);
  nor (_02489_, _02487_, \oc8051_golden_model_1.ACC [2]);
  nor (_02490_, _02489_, _02488_);
  not (_02491_, _02490_);
  and (_02492_, _02491_, _02484_);
  nor (_02493_, _02491_, _02484_);
  nor (_02494_, _02493_, _02492_);
  and (_02495_, _02494_, _02476_);
  and (_02496_, _02313_, _02298_);
  or (_02497_, _02345_, _02496_);
  or (_02498_, _02283_, _02497_);
  or (_02499_, _02474_, _02498_);
  and (_02500_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  and (_02501_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_02502_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor (_02503_, _02502_, _02500_);
  and (_02504_, _02503_, _02501_);
  nor (_02505_, _02504_, _02500_);
  and (_02506_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_02507_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor (_02508_, _02507_, _02506_);
  not (_02509_, _02508_);
  nor (_02510_, _02509_, _02505_);
  and (_02511_, _02509_, _02505_);
  nor (_02512_, _02511_, _02510_);
  not (_02513_, _02512_);
  or (_02514_, _02513_, _02499_);
  nand (_02515_, _02471_, _02456_);
  or (_02516_, _02515_, _02441_);
  or (_02517_, _02516_, _02410_);
  nor (_02518_, _02498_, _02517_);
  nand (_02519_, _02440_, _02425_);
  and (_02520_, _02472_, _02519_);
  and (_02521_, _02408_, _02393_);
  and (_02522_, _02521_, _02378_);
  and (_02523_, _02522_, _02520_);
  and (_02524_, _02523_, _02347_);
  nor (_02525_, _02524_, _02518_);
  and (_02526_, _02525_, _02514_);
  and (_02527_, _02344_, _02329_);
  or (_02528_, _02527_, _02314_);
  or (_02529_, _02528_, _02283_);
  or (_02530_, _02529_, _02517_);
  or (_02531_, _02527_, _02496_);
  or (_02532_, _02531_, _02283_);
  or (_02533_, _02532_, _02517_);
  and (_02534_, _02533_, _02530_);
  and (_02535_, _02250_, _02224_);
  or (_02536_, _02282_, _02535_);
  or (_02537_, _02536_, _02346_);
  or (_02538_, _02537_, _02517_);
  or (_02539_, _02536_, _02497_);
  or (_02540_, _02539_, _02517_);
  and (_02541_, _02540_, _02538_);
  and (_02542_, _02541_, _02534_);
  or (_02543_, _02536_, _02528_);
  or (_02544_, _02543_, _02517_);
  or (_02545_, _02536_, _02531_);
  or (_02546_, _02545_, _02517_);
  and (_02547_, _02546_, _02544_);
  nand (_02548_, _02547_, _02542_);
  or (_02549_, _02548_, _02487_);
  nand (_02550_, _02549_, _02499_);
  nand (_02551_, _02550_, _02526_);
  not (_02552_, _02476_);
  and (_02553_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_02554_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor (_02555_, _02554_, _02553_);
  and (_02556_, _02547_, _02542_);
  and (_02557_, _02556_, _02525_);
  or (_02558_, _02557_, _02555_);
  and (_02559_, _02558_, _02552_);
  and (_02560_, _02559_, _02551_);
  or (_02561_, _02560_, _02495_);
  and (_02562_, _02377_, _02362_);
  and (_02563_, _02521_, _02562_);
  and (_02564_, _02520_, _02563_);
  not (_02565_, _02346_);
  and (_02566_, _02282_, _02535_);
  and (_02567_, _02566_, _02565_);
  and (_02568_, _02567_, _02564_);
  not (_02569_, _02568_);
  not (_02570_, _02497_);
  and (_02571_, _02566_, _02570_);
  and (_02572_, _02571_, _02564_);
  and (_02573_, _02345_, _02496_);
  and (_02574_, _02566_, _02573_);
  and (_02575_, _02574_, _02564_);
  nor (_02576_, _02575_, _02572_);
  and (_02577_, _02576_, _02569_);
  and (_02578_, _02347_, _02564_);
  not (_02579_, _02578_);
  and (_02580_, _02282_, _02251_);
  and (_02581_, _02580_, _02573_);
  and (_02582_, _02581_, _02564_);
  and (_02583_, _02345_, _02314_);
  and (_02584_, _02580_, _02583_);
  and (_02585_, _02584_, _02564_);
  nor (_02586_, _02585_, _02582_);
  and (_02587_, _02586_, _02579_);
  and (_02588_, _02580_, _02565_);
  and (_02589_, _02588_, _02564_);
  not (_02590_, _02589_);
  and (_02591_, _02566_, _02583_);
  and (_02592_, _02591_, _02564_);
  and (_02593_, _02580_, _02570_);
  and (_02594_, _02593_, _02564_);
  nor (_02595_, _02594_, _02592_);
  and (_02596_, _02595_, _02590_);
  and (_02597_, _02596_, _02587_);
  and (_02598_, _02597_, _02577_);
  nand (_02599_, _02598_, _02561_);
  not (_02600_, _02555_);
  nor (_02601_, _02598_, _02600_);
  not (_02602_, _02601_);
  and (_02603_, _02602_, _02599_);
  nor (_02604_, _02493_, _02488_);
  not (_02605_, \oc8051_golden_model_1.ACC [3]);
  not (_02606_, _02205_);
  nor (_02607_, _02485_, _02194_);
  nor (_02608_, _02607_, _02606_);
  nor (_02609_, _02608_, _02605_);
  and (_02610_, _02608_, _02605_);
  nor (_02611_, _02610_, _02609_);
  and (_02612_, _02611_, _02604_);
  nor (_02613_, _02611_, _02604_);
  nor (_02614_, _02613_, _02612_);
  nor (_02615_, _02614_, _02552_);
  not (_02616_, _02608_);
  or (_02617_, _02548_, _02616_);
  nor (_02618_, _02211_, _02198_);
  nor (_02619_, _02553_, \oc8051_golden_model_1.PC [3]);
  nor (_02620_, _02619_, _02618_);
  or (_02621_, _02620_, _02556_);
  and (_02622_, _02621_, _02617_);
  nand (_02623_, _02622_, _02499_);
  nor (_02624_, _02510_, _02506_);
  and (_02625_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_02626_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor (_02627_, _02626_, _02625_);
  not (_02628_, _02627_);
  nor (_02629_, _02628_, _02624_);
  and (_02630_, _02628_, _02624_);
  nor (_02631_, _02630_, _02629_);
  not (_02632_, _02631_);
  or (_02633_, _02632_, _02499_);
  and (_02634_, _02633_, _02525_);
  nand (_02635_, _02634_, _02623_);
  or (_02636_, _02620_, _02525_);
  and (_02637_, _02636_, _02552_);
  and (_02638_, _02637_, _02635_);
  or (_02639_, _02638_, _02615_);
  and (_02640_, _02639_, _02598_);
  not (_02641_, _02620_);
  nor (_02642_, _02641_, _02598_);
  nor (_02643_, _02642_, _02640_);
  or (_02644_, _02643_, _02603_);
  or (_02645_, _02548_, _02225_);
  or (_02646_, _02556_, \oc8051_golden_model_1.PC [0]);
  nand (_02647_, _02646_, _02645_);
  nand (_02648_, _02647_, _02499_);
  nor (_02649_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor (_02650_, _02649_, _02501_);
  or (_02651_, _02650_, _02499_);
  and (_02652_, _02651_, _02525_);
  and (_02653_, _02652_, _02648_);
  nor (_02654_, _02525_, _02225_);
  or (_02655_, _02654_, _02653_);
  nand (_02656_, _02655_, _02552_);
  not (_02657_, _02598_);
  not (_02658_, \oc8051_golden_model_1.ACC [0]);
  and (_02659_, _02658_, \oc8051_golden_model_1.PC [0]);
  nor (_02660_, _02659_, _02480_);
  and (_02661_, _02660_, _02476_);
  nor (_02662_, _02661_, _02657_);
  nand (_02663_, _02662_, _02656_);
  nor (_02664_, _02598_, \oc8051_golden_model_1.PC [0]);
  not (_02665_, _02664_);
  nand (_02666_, _02665_, _02663_);
  and (_02667_, _02499_, _02478_);
  and (_02668_, _02667_, _02547_);
  nand (_02669_, _02668_, _02542_);
  nor (_02670_, _02503_, _02501_);
  nor (_02671_, _02670_, _02504_);
  or (_02672_, _02671_, _02499_);
  nand (_02673_, _02672_, _02669_);
  nand (_02674_, _02673_, _02525_);
  or (_02675_, _02557_, _02198_);
  nand (_02676_, _02675_, _02674_);
  and (_02677_, _02676_, _02552_);
  nor (_02678_, _02482_, _02480_);
  nor (_02679_, _02678_, _02483_);
  nor (_02680_, _02679_, _02552_);
  or (_02681_, _02680_, _02677_);
  nand (_02682_, _02681_, _02598_);
  nor (_02683_, _02598_, _02198_);
  not (_02684_, _02683_);
  nand (_02685_, _02684_, _02682_);
  or (_02686_, _02685_, _02666_);
  or (_02687_, _02686_, _02644_);
  or (_02688_, _02687_, _33745_);
  and (_02689_, _02665_, _02663_);
  or (_02690_, _02685_, _02689_);
  nand (_02691_, _02602_, _02599_);
  or (_02692_, _02643_, _02691_);
  or (_02693_, _02692_, _02690_);
  or (_02694_, _02693_, _33540_);
  and (_02695_, _02694_, _02688_);
  or (_02696_, _02642_, _02640_);
  or (_02697_, _02696_, _02603_);
  or (_02698_, _02697_, _02686_);
  or (_02699_, _02698_, _33417_);
  and (_02700_, _02684_, _02682_);
  or (_02701_, _02700_, _02666_);
  or (_02702_, _02696_, _02691_);
  or (_02703_, _02702_, _02701_);
  or (_02704_, _02703_, _33171_);
  and (_02705_, _02704_, _02699_);
  and (_02706_, _02705_, _02695_);
  or (_02707_, _02692_, _02701_);
  or (_02708_, _02707_, _33499_);
  or (_02709_, _02700_, _02689_);
  or (_02710_, _02692_, _02709_);
  or (_02711_, _02710_, _33458_);
  and (_02712_, _02711_, _02708_);
  or (_02713_, _02690_, _02644_);
  or (_02714_, _02713_, _33704_);
  or (_02715_, _02709_, _02644_);
  or (_02716_, _02715_, _33622_);
  and (_02717_, _02716_, _02714_);
  and (_02718_, _02717_, _02712_);
  and (_02719_, _02718_, _02706_);
  or (_02720_, _02697_, _02701_);
  or (_02721_, _02720_, _33335_);
  or (_02722_, _02702_, _02686_);
  or (_02723_, _02722_, _33253_);
  and (_02724_, _02723_, _02721_);
  or (_02725_, _02697_, _02690_);
  or (_02726_, _02725_, _33376_);
  or (_02727_, _02697_, _02709_);
  or (_02728_, _02727_, _33294_);
  and (_02729_, _02728_, _02726_);
  and (_02730_, _02729_, _02724_);
  or (_02731_, _02701_, _02644_);
  or (_02732_, _02731_, _33663_);
  or (_02733_, _02692_, _02686_);
  or (_02734_, _02733_, _33581_);
  and (_02735_, _02734_, _02732_);
  or (_02736_, _02702_, _02709_);
  or (_02737_, _02736_, _33130_);
  or (_02738_, _02702_, _02690_);
  or (_02739_, _02738_, _33212_);
  and (_02740_, _02739_, _02737_);
  and (_02741_, _02740_, _02735_);
  and (_02742_, _02741_, _02730_);
  and (_02743_, _02742_, _02719_);
  or (_02744_, _02693_, _33560_);
  or (_02745_, _02736_, _33150_);
  and (_02746_, _02745_, _02744_);
  or (_02747_, _02731_, _33683_);
  or (_02748_, _02727_, _33314_);
  and (_02749_, _02748_, _02747_);
  and (_02750_, _02749_, _02746_);
  or (_02751_, _02707_, _33519_);
  or (_02752_, _02710_, _33478_);
  and (_02753_, _02752_, _02751_);
  or (_02754_, _02713_, _33724_);
  or (_02755_, _02722_, _33273_);
  and (_02756_, _02755_, _02754_);
  and (_02757_, _02756_, _02753_);
  and (_02758_, _02757_, _02750_);
  or (_02759_, _02698_, _33437_);
  or (_02760_, _02725_, _33396_);
  and (_02761_, _02760_, _02759_);
  or (_02762_, _02720_, _33355_);
  or (_02763_, _02703_, _33191_);
  and (_02764_, _02763_, _02762_);
  and (_02765_, _02764_, _02761_);
  or (_02766_, _02733_, _33601_);
  or (_02767_, _02738_, _33232_);
  and (_02768_, _02767_, _02766_);
  or (_02769_, _02687_, _33765_);
  or (_02770_, _02715_, _33642_);
  and (_02771_, _02770_, _02769_);
  and (_02772_, _02771_, _02768_);
  and (_02773_, _02772_, _02765_);
  nand (_02774_, _02773_, _02758_);
  and (_02775_, _02774_, _02743_);
  and (_02776_, _02472_, _02441_);
  and (_02777_, _02776_, _02563_);
  and (_02778_, _02777_, _02571_);
  and (_02779_, _02778_, _02775_);
  and (_02780_, _02778_, _02743_);
  not (_02781_, _02780_);
  not (_02782_, _02498_);
  and (_02783_, _02515_, _02441_);
  and (_02784_, _02783_, _02563_);
  and (_02785_, _02784_, _02782_);
  and (_02786_, _02775_, _02785_);
  not (_02787_, \oc8051_golden_model_1.SP [0]);
  nor (_02788_, _02533_, _02787_);
  not (_02789_, _02532_);
  and (_02790_, _02789_, _02784_);
  and (_02791_, _02790_, _02775_);
  and (_02792_, _02790_, _02743_);
  not (_02793_, _02792_);
  not (_02794_, _02537_);
  and (_02795_, _02777_, _02794_);
  and (_02796_, _02794_, _02784_);
  and (_02797_, _02796_, _02775_);
  not (_02798_, _02539_);
  and (_02799_, _02798_, _02784_);
  and (_02800_, _02799_, _02775_);
  nand (_02801_, _02281_, _02266_);
  and (_02802_, _02801_, _02251_);
  and (_02803_, _02802_, _02583_);
  and (_02804_, _02803_, _02564_);
  or (_02805_, _02713_, _33709_);
  or (_02806_, _02731_, _33668_);
  and (_02807_, _02806_, _02805_);
  or (_02808_, _02733_, _33586_);
  or (_02809_, _02693_, _33545_);
  and (_02810_, _02809_, _02808_);
  and (_02811_, _02810_, _02807_);
  or (_02812_, _02720_, _33340_);
  or (_02813_, _02736_, _33135_);
  and (_02814_, _02813_, _02812_);
  or (_02815_, _02722_, _33258_);
  or (_02816_, _02703_, _33176_);
  and (_02817_, _02816_, _02815_);
  and (_02818_, _02817_, _02814_);
  and (_02819_, _02818_, _02811_);
  or (_02820_, _02707_, _33504_);
  or (_02821_, _02710_, _33463_);
  and (_02822_, _02821_, _02820_);
  or (_02823_, _02687_, _33750_);
  or (_02824_, _02715_, _33627_);
  and (_02825_, _02824_, _02823_);
  and (_02826_, _02825_, _02822_);
  or (_02827_, _02698_, _33422_);
  or (_02828_, _02725_, _33381_);
  and (_02829_, _02828_, _02827_);
  or (_02830_, _02727_, _33299_);
  or (_02831_, _02738_, _33217_);
  and (_02832_, _02831_, _02830_);
  and (_02833_, _02832_, _02829_);
  and (_02834_, _02833_, _02826_);
  and (_02835_, _02834_, _02819_);
  not (_02836_, _02835_);
  and (_02837_, _02803_, _02523_);
  and (_02838_, _02837_, _02743_);
  and (_02839_, _02838_, _02836_);
  nor (_02840_, _02839_, _02804_);
  and (_02841_, _02441_, _02409_);
  and (_02842_, _02841_, _02803_);
  nor (_02843_, _02842_, _02838_);
  not (_02844_, _02843_);
  and (_02845_, _02844_, _02840_);
  and (_02846_, _02804_, \oc8051_golden_model_1.SP [0]);
  and (_02847_, _02841_, _02798_);
  nor (_02848_, _02847_, _02846_);
  not (_02849_, _02848_);
  nor (_02850_, _02849_, _02845_);
  not (_02851_, _02850_);
  and (_02852_, _02567_, _02523_);
  not (_02853_, _02852_);
  and (_02854_, _02574_, _02784_);
  not (_02855_, _02854_);
  and (_02856_, _02574_, _02523_);
  not (_02857_, _02856_);
  not (_02858_, _02743_);
  nor (_02859_, _02687_, _33780_);
  nor (_02860_, _02733_, _33616_);
  nor (_02861_, _02860_, _02859_);
  nor (_02862_, _02698_, _33452_);
  nor (_02863_, _02736_, _33165_);
  nor (_02864_, _02863_, _02862_);
  and (_02865_, _02864_, _02861_);
  nor (_02866_, _02713_, _33739_);
  nor (_02867_, _02731_, _33698_);
  nor (_02868_, _02867_, _02866_);
  nor (_02869_, _02693_, _33575_);
  nor (_02870_, _02707_, _33534_);
  nor (_02871_, _02870_, _02869_);
  and (_02872_, _02871_, _02868_);
  and (_02873_, _02872_, _02865_);
  nor (_02874_, _02727_, _33329_);
  nor (_02875_, _02722_, _33288_);
  nor (_02876_, _02875_, _02874_);
  nor (_02877_, _02725_, _33411_);
  nor (_02878_, _02720_, _33370_);
  nor (_02879_, _02878_, _02877_);
  and (_02880_, _02879_, _02876_);
  nor (_02881_, _02738_, _33247_);
  nor (_02882_, _02703_, _33206_);
  nor (_02883_, _02882_, _02881_);
  nor (_02884_, _02715_, _33657_);
  nor (_02885_, _02710_, _33493_);
  nor (_02886_, _02885_, _02884_);
  and (_02887_, _02886_, _02883_);
  and (_02888_, _02887_, _02880_);
  and (_02889_, _02888_, _02873_);
  nor (_02890_, _02889_, _02858_);
  and (_02891_, _02774_, _02858_);
  nor (_02892_, _02891_, _02890_);
  and (_02893_, _02584_, _02784_);
  and (_02894_, _02347_, _02784_);
  nor (_02895_, _02894_, _02893_);
  not (_02896_, _02895_);
  and (_02897_, _02896_, _02892_);
  and (_02898_, _02523_, _02782_);
  not (_02899_, _02898_);
  not (_02900_, _02529_);
  and (_02901_, _02777_, _02900_);
  and (_02902_, _02900_, _02784_);
  nor (_02903_, _02902_, _02901_);
  and (_02904_, _02409_, _02562_);
  and (_02905_, _02904_, _02783_);
  and (_02906_, _02409_, _02378_);
  and (_02907_, _02906_, _02776_);
  nor (_02908_, _02907_, _02905_);
  nor (_02909_, _02908_, _02529_);
  not (_02910_, _02909_);
  not (_02911_, _02776_);
  and (_02912_, _02906_, _02911_);
  and (_02913_, _02912_, _02900_);
  not (_02914_, _02904_);
  nor (_02915_, _02914_, _02529_);
  and (_02916_, _02915_, _02519_);
  nor (_02917_, _02916_, _02913_);
  and (_02918_, _02917_, _02910_);
  and (_02919_, _02904_, _02776_);
  and (_02920_, _02919_, _02900_);
  not (_02921_, _02920_);
  and (_02922_, _02921_, _02918_);
  not (_02923_, _02922_);
  and (_02924_, _02923_, _02774_);
  and (_02925_, _02777_, _02789_);
  nor (_02926_, _02790_, _02925_);
  not (_02927_, _02796_);
  and (_02928_, _02794_, _02523_);
  and (_02929_, _02928_, _02774_);
  and (_02930_, _02777_, _02798_);
  and (_02931_, _02930_, \oc8051_golden_model_1.SP [3]);
  and (_02932_, _02798_, _02523_);
  and (_02933_, _02802_, _02573_);
  and (_02934_, _02933_, _02523_);
  nor (_02935_, _02934_, _02932_);
  or (_02936_, _02935_, _02774_);
  not (_02937_, \oc8051_golden_model_1.PSW [3]);
  nand (_02938_, _02935_, _02937_);
  nor (_02939_, _02799_, _02930_);
  and (_02940_, _02939_, _02938_);
  and (_02941_, _02940_, _02936_);
  or (_02942_, _02941_, _02931_);
  not (_02943_, _02928_);
  and (_02944_, _02789_, _02523_);
  nor (_02945_, _02944_, _02795_);
  and (_02946_, _02945_, _02943_);
  and (_02947_, _02946_, _02922_);
  and (_02948_, _02947_, _02942_);
  or (_02949_, _02948_, _02929_);
  and (_02950_, _02949_, _02927_);
  not (_02951_, _02945_);
  and (_02952_, _02951_, _02774_);
  or (_02953_, _02952_, _02950_);
  and (_02954_, _02953_, _02926_);
  or (_02955_, _02954_, _02924_);
  and (_02956_, _02955_, _02903_);
  nor (_02957_, _02799_, _02796_);
  and (_02958_, _02957_, _02926_);
  and (_02959_, _02958_, _02903_);
  nor (_02960_, _02959_, _02892_);
  or (_02961_, _02960_, _02956_);
  and (_02962_, _02961_, _02899_);
  and (_02963_, _02898_, _02774_);
  nor (_02964_, _02963_, _02962_);
  or (_02965_, _02964_, _02785_);
  not (_02966_, _02785_);
  or (_02967_, _02892_, _02966_);
  and (_02968_, _02967_, _02965_);
  or (_02969_, _02968_, _02524_);
  not (_02970_, _02524_);
  and (_02971_, _02522_, _02515_);
  and (_02972_, _02971_, _02789_);
  nor (_02973_, _02972_, _02944_);
  and (_02974_, _02584_, _02523_);
  and (_02975_, _02777_, _02782_);
  nor (_02976_, _02975_, _02974_);
  and (_02977_, _02581_, _02475_);
  and (_02978_, _02776_, _02522_);
  and (_02979_, _02978_, _02789_);
  nor (_02980_, _02979_, _02977_);
  and (_02981_, _02980_, _02976_);
  and (_02982_, _02567_, _02784_);
  and (_02983_, _02906_, _02783_);
  and (_02984_, _02983_, _02789_);
  nor (_02985_, _02984_, _02982_);
  and (_02986_, _02985_, _02981_);
  and (_02987_, _02986_, _02973_);
  and (_02988_, _02571_, _02784_);
  nor (_02989_, _02988_, _02778_);
  and (_02990_, _02777_, _02574_);
  and (_02991_, _02593_, _02475_);
  nor (_02992_, _02991_, _02990_);
  and (_02993_, _02777_, _02591_);
  and (_02994_, _02588_, _02475_);
  nor (_02995_, _02994_, _02993_);
  and (_02996_, _02995_, _02992_);
  and (_02997_, _02996_, _02989_);
  and (_02998_, _02919_, _02789_);
  and (_02999_, _02906_, _02520_);
  and (_03000_, _02999_, _02789_);
  or (_03001_, _03000_, _02998_);
  not (_03002_, _03001_);
  not (_03003_, _02473_);
  and (_03004_, _02906_, _03003_);
  and (_03005_, _03004_, _02789_);
  nor (_03006_, _03005_, _02932_);
  and (_03007_, _03006_, _03002_);
  and (_03008_, _02904_, _02520_);
  or (_03009_, _03008_, _02905_);
  not (_03010_, _03009_);
  and (_03011_, _02904_, _03003_);
  nor (_03012_, _03011_, _02907_);
  nand (_03013_, _03012_, _03010_);
  and (_03014_, _03013_, _02789_);
  not (_03015_, _03014_);
  and (_03016_, _03015_, _03007_);
  and (_03017_, _03016_, _02997_);
  and (_03018_, _03017_, _02987_);
  or (_03019_, _03018_, _02225_);
  nand (_03020_, _03018_, _02225_);
  nand (_03021_, _03020_, _03019_);
  and (_03022_, _03020_, \oc8051_golden_model_1.PC [1]);
  nor (_03023_, _03020_, \oc8051_golden_model_1.PC [1]);
  nor (_03024_, _03023_, _03022_);
  not (_03025_, _03024_);
  nor (_03026_, _03025_, _03021_);
  nor (_03027_, _03018_, _02600_);
  and (_03028_, _03018_, _02487_);
  nor (_03029_, _03028_, _03027_);
  nor (_03030_, _03018_, _02641_);
  and (_03031_, _03018_, _02616_);
  nor (_03032_, _03031_, _03030_);
  nor (_03033_, _03032_, _03029_);
  and (_03034_, _03033_, _03026_);
  and (_03035_, _03034_, _01387_);
  and (_03036_, _03025_, _03021_);
  and (_03037_, _03036_, _03033_);
  and (_03038_, _03037_, _01389_);
  nor (_03039_, _03038_, _03035_);
  and (_03040_, _03024_, _03021_);
  not (_03041_, _03032_);
  nor (_03042_, _03041_, _03029_);
  and (_03043_, _03042_, _03040_);
  and (_03044_, _03043_, _01401_);
  and (_03045_, _03032_, _03029_);
  and (_03046_, _03045_, _03040_);
  and (_03047_, _03046_, _01396_);
  nor (_03048_, _03047_, _03044_);
  and (_03049_, _03048_, _03039_);
  and (_03050_, _03042_, _03026_);
  and (_03051_, _03050_, _01409_);
  and (_03052_, _03042_, _03036_);
  and (_03053_, _03052_, _01411_);
  nor (_03054_, _03053_, _03051_);
  and (_03055_, _03045_, _03026_);
  and (_03056_, _03055_, _01379_);
  and (_03057_, _03045_, _03036_);
  and (_03058_, _03057_, _01407_);
  nor (_03059_, _03058_, _03056_);
  and (_03060_, _03059_, _03054_);
  and (_03061_, _03060_, _03049_);
  and (_03062_, _03041_, _03029_);
  and (_03063_, _03062_, _03026_);
  and (_03064_, _03063_, _01383_);
  nor (_03065_, _03024_, _03021_);
  and (_03066_, _03065_, _03062_);
  and (_03067_, _03066_, _01420_);
  nor (_03068_, _03067_, _03064_);
  and (_03069_, _03040_, _03033_);
  and (_03070_, _03069_, _01394_);
  and (_03071_, _03065_, _03033_);
  and (_03072_, _03071_, _01392_);
  nor (_03073_, _03072_, _03070_);
  and (_03074_, _03073_, _03068_);
  and (_03075_, _03065_, _03042_);
  and (_03076_, _03075_, _01413_);
  and (_03077_, _03065_, _03045_);
  and (_03078_, _03077_, _01381_);
  nor (_03079_, _03078_, _03076_);
  and (_03080_, _03062_, _03040_);
  and (_03081_, _03080_, _01399_);
  and (_03082_, _03062_, _03036_);
  and (_03083_, _03082_, _01418_);
  nor (_03084_, _03083_, _03081_);
  and (_03085_, _03084_, _03079_);
  and (_03086_, _03085_, _03074_);
  and (_03087_, _03086_, _03061_);
  nor (_03088_, _03087_, _02970_);
  nor (_03089_, _03088_, _02896_);
  and (_03090_, _03089_, _02969_);
  or (_03091_, _03090_, _02897_);
  and (_03092_, _02593_, _02523_);
  not (_03093_, _03092_);
  and (_03094_, _02593_, _02784_);
  nor (_03095_, _03094_, _02991_);
  and (_03096_, _03095_, _03093_);
  and (_03097_, _02588_, _02523_);
  not (_03098_, _03097_);
  and (_03099_, _02588_, _02784_);
  nor (_03100_, _03099_, _02994_);
  and (_03101_, _03100_, _03098_);
  and (_03102_, _03101_, _03096_);
  and (_03103_, _02591_, _02523_);
  not (_03104_, _03103_);
  and (_03105_, _02581_, _02523_);
  not (_03106_, _03105_);
  and (_03107_, _02581_, _02784_);
  nor (_03108_, _03107_, _02977_);
  and (_03109_, _03108_, _03106_);
  and (_03110_, _03109_, _03104_);
  and (_03111_, _03110_, _03102_);
  nand (_03112_, _03111_, _03091_);
  and (_03113_, _02591_, _02784_);
  nor (_03114_, _03111_, _02774_);
  nor (_03115_, _03114_, _03113_);
  and (_03116_, _03115_, _03112_);
  and (_03117_, _03113_, \oc8051_golden_model_1.SP [3]);
  or (_03118_, _03117_, _02993_);
  nor (_03119_, _03118_, _03116_);
  and (_03120_, _02892_, _02993_);
  or (_03121_, _03120_, _03119_);
  nand (_03122_, _03121_, _02857_);
  and (_03123_, _02574_, _02522_);
  and (_03124_, _03123_, _02520_);
  not (_03125_, _03124_);
  or (_03126_, _03125_, _02774_);
  nand (_03127_, _03126_, _03122_);
  nand (_03128_, _03127_, _02855_);
  not (_03129_, \oc8051_golden_model_1.SP [3]);
  and (_03130_, _02854_, _03129_);
  nor (_03131_, _03130_, _02990_);
  nand (_03132_, _03131_, _03128_);
  and (_03133_, _02571_, _02523_);
  not (_03134_, _02990_);
  nor (_03135_, _03134_, _02892_);
  nor (_03136_, _03135_, _03133_);
  nand (_03137_, _03136_, _03132_);
  not (_03138_, _03133_);
  nor (_03139_, _03138_, _02774_);
  nor (_03140_, _03139_, _02778_);
  and (_03141_, _03140_, _03137_);
  not (_03142_, _02778_);
  nor (_03143_, _03142_, _02892_);
  or (_03144_, _03143_, _03141_);
  nand (_03145_, _03144_, _02853_);
  and (_03146_, _02852_, _02774_);
  not (_03147_, _03146_);
  and (_03148_, _03147_, _03145_);
  nor (_03149_, _02703_, _33201_);
  nor (_03150_, _02738_, _33242_);
  nor (_03151_, _03150_, _03149_);
  nor (_03152_, _02715_, _33652_);
  nor (_03153_, _02725_, _33406_);
  nor (_03154_, _03153_, _03152_);
  and (_03155_, _03154_, _03151_);
  nor (_03156_, _02733_, _33611_);
  nor (_03157_, _02710_, _33488_);
  nor (_03158_, _03157_, _03156_);
  nor (_03159_, _02720_, _33365_);
  nor (_03160_, _02736_, _33160_);
  nor (_03161_, _03160_, _03159_);
  and (_03162_, _03161_, _03158_);
  and (_03163_, _03162_, _03155_);
  nor (_03164_, _02687_, _33775_);
  nor (_03165_, _02713_, _33734_);
  nor (_03166_, _03165_, _03164_);
  nor (_03167_, _02731_, _33693_);
  nor (_03168_, _02707_, _33529_);
  nor (_03169_, _03168_, _03167_);
  and (_03170_, _03169_, _03166_);
  nor (_03171_, _02693_, _33570_);
  nor (_03172_, _02722_, _33283_);
  nor (_03173_, _03172_, _03171_);
  nor (_03174_, _02698_, _33447_);
  nor (_03175_, _02727_, _33324_);
  nor (_03176_, _03175_, _03174_);
  and (_03177_, _03176_, _03173_);
  and (_03178_, _03177_, _03170_);
  and (_03179_, _03178_, _03163_);
  nor (_03180_, _03179_, _02858_);
  not (_03181_, _03180_);
  nor (_03182_, _02778_, _02796_);
  nor (_03183_, _02990_, _02993_);
  and (_03184_, _03183_, _02966_);
  and (_03185_, _03184_, _03182_);
  not (_03186_, _02799_);
  and (_03187_, _03186_, _02895_);
  and (_03188_, _02926_, _02903_);
  and (_03189_, _03188_, _03187_);
  and (_03190_, _03189_, _03185_);
  nor (_03191_, _03190_, _03181_);
  not (_03192_, _03191_);
  and (_03193_, _03071_, _01346_);
  and (_03194_, _03080_, _01353_);
  nor (_03195_, _03194_, _03193_);
  and (_03196_, _03050_, _01367_);
  and (_03197_, _03077_, _01361_);
  nor (_03198_, _03197_, _03196_);
  and (_03199_, _03198_, _03195_);
  and (_03200_, _03063_, _01372_);
  and (_03201_, _03082_, _01333_);
  nor (_03202_, _03201_, _03200_);
  and (_03203_, _03069_, _01348_);
  and (_03204_, _03037_, _01343_);
  nor (_03205_, _03204_, _03203_);
  and (_03206_, _03205_, _03202_);
  and (_03207_, _03206_, _03199_);
  and (_03208_, _03075_, _01363_);
  and (_03209_, _03046_, _01355_);
  nor (_03210_, _03209_, _03208_);
  and (_03211_, _03043_, _01350_);
  and (_03212_, _03052_, _01365_);
  nor (_03213_, _03212_, _03211_);
  and (_03214_, _03213_, _03210_);
  and (_03215_, _03055_, _01337_);
  and (_03216_, _03057_, _01335_);
  nor (_03217_, _03216_, _03215_);
  and (_03218_, _03034_, _01341_);
  and (_03219_, _03066_, _01374_);
  nor (_03220_, _03219_, _03218_);
  and (_03221_, _03220_, _03217_);
  and (_03222_, _03221_, _03214_);
  and (_03223_, _03222_, _03207_);
  nor (_03224_, _03223_, _02970_);
  and (_03225_, _02907_, _02593_);
  and (_03226_, _02999_, _02593_);
  nor (_03227_, _03226_, _03225_);
  and (_03228_, _02907_, _02571_);
  and (_03229_, _02999_, _02571_);
  nor (_03230_, _03229_, _03228_);
  and (_03231_, _02906_, _02515_);
  and (_03232_, _03231_, _02789_);
  and (_03233_, _03231_, _02782_);
  nor (_03234_, _03233_, _03232_);
  and (_03235_, _03231_, _02591_);
  and (_03236_, _03231_, _02571_);
  nor (_03237_, _03236_, _03235_);
  and (_03238_, _03237_, _03234_);
  and (_03239_, _03238_, _03230_);
  and (_03240_, _03239_, _03227_);
  and (_03241_, _03231_, _02794_);
  and (_03242_, _02906_, _02588_);
  nor (_03243_, _03242_, _03241_);
  and (_03244_, _02906_, _02472_);
  and (_03245_, _03244_, _02581_);
  and (_03246_, _03231_, _02347_);
  nor (_03247_, _03246_, _03245_);
  and (_03248_, _03247_, _03243_);
  and (_03249_, _03244_, _02574_);
  not (_03250_, _03249_);
  and (_03251_, _03244_, _02591_);
  and (_03252_, _03244_, _02789_);
  nor (_03253_, _03252_, _03251_);
  and (_03254_, _03253_, _03250_);
  and (_03255_, _03254_, _03248_);
  not (_03256_, \oc8051_golden_model_1.SP [2]);
  nor (_03257_, _02930_, _03113_);
  nor (_03258_, _03257_, _03256_);
  and (_03259_, _03231_, _02581_);
  and (_03260_, _03231_, _02574_);
  nor (_03261_, _03260_, _03259_);
  not (_03262_, _03261_);
  nor (_03263_, _03262_, _03258_);
  and (_03264_, _03263_, _03255_);
  and (_03265_, _02907_, _02347_);
  and (_03266_, _02999_, _02782_);
  nor (_03267_, _03266_, _03265_);
  and (_03268_, _02907_, _02782_);
  not (_03269_, _02906_);
  nor (_03270_, _02567_, _02933_);
  nor (_03271_, _03270_, _03269_);
  nor (_03272_, _03271_, _03268_);
  and (_03273_, _03272_, _03267_);
  and (_03274_, _03244_, _02794_);
  and (_03275_, _03244_, _02798_);
  nor (_03276_, _03275_, _03274_);
  and (_03277_, _03231_, _02798_);
  and (_03278_, _03231_, _02593_);
  nor (_03279_, _03278_, _03277_);
  and (_03280_, _03279_, _03276_);
  and (_03281_, _02854_, \oc8051_golden_model_1.SP [2]);
  and (_03282_, _02999_, _02347_);
  nor (_03283_, _03282_, _03281_);
  and (_03284_, _03283_, _03280_);
  and (_03285_, _03284_, _03273_);
  and (_03286_, _03285_, _03264_);
  and (_03287_, _03286_, _03240_);
  not (_03288_, _03287_);
  nor (_03289_, _03288_, _03224_);
  nor (_03290_, _02687_, _33760_);
  nor (_03291_, _02736_, _33145_);
  nor (_03292_, _03291_, _03290_);
  nor (_03293_, _02733_, _33596_);
  nor (_03294_, _02703_, _33186_);
  nor (_03295_, _03294_, _03293_);
  and (_03296_, _03295_, _03292_);
  nor (_03297_, _02707_, _33514_);
  nor (_03298_, _02738_, _33227_);
  nor (_03299_, _03298_, _03297_);
  nor (_03300_, _02698_, _33432_);
  nor (_03301_, _02720_, _33350_);
  nor (_03302_, _03301_, _03300_);
  and (_03303_, _03302_, _03299_);
  and (_03304_, _03303_, _03296_);
  nor (_03305_, _02722_, _33268_);
  nor (_03306_, _02727_, _33309_);
  nor (_03307_, _03306_, _03305_);
  nor (_03308_, _02713_, _33719_);
  nor (_03309_, _02693_, _33555_);
  nor (_03310_, _03309_, _03308_);
  and (_03311_, _03310_, _03307_);
  nor (_03312_, _02731_, _33678_);
  nor (_03313_, _02710_, _33473_);
  nor (_03314_, _03313_, _03312_);
  nor (_03315_, _02715_, _33637_);
  nor (_03316_, _02725_, _33391_);
  nor (_03317_, _03316_, _03315_);
  and (_03318_, _03317_, _03314_);
  and (_03319_, _03318_, _03311_);
  and (_03320_, _03319_, _03304_);
  not (_03321_, _03320_);
  and (_03322_, _02945_, _02935_);
  and (_03323_, _03322_, _03125_);
  nor (_03324_, _02928_, _02898_);
  and (_03325_, _03324_, _03104_);
  and (_03326_, _03325_, _03101_);
  and (_03327_, _03326_, _03323_);
  nand (_03328_, _03327_, _02922_);
  not (_03329_, _03109_);
  nor (_03330_, _03133_, _02852_);
  nand (_03331_, _03330_, _03096_);
  or (_03332_, _03331_, _03329_);
  or (_03333_, _03332_, _03328_);
  and (_03334_, _03333_, _03321_);
  not (_03335_, _03334_);
  and (_03336_, _03335_, _03289_);
  and (_03337_, _03336_, _03192_);
  not (_03338_, \oc8051_golden_model_1.IRAM[0] [0]);
  not (_03339_, _02775_);
  nor (_03340_, _02903_, _03339_);
  or (_03341_, _02943_, _02835_);
  nor (_03342_, _02935_, _02835_);
  and (_03343_, _02971_, _02933_);
  and (_03344_, _02906_, _02933_);
  and (_03345_, _02971_, _02803_);
  or (_03346_, _03345_, _03344_);
  or (_03347_, _03346_, _03343_);
  and (_03348_, _03347_, _02441_);
  and (_03349_, _02919_, _02933_);
  and (_03350_, _02905_, _02933_);
  and (_03351_, _02803_, _02784_);
  or (_03352_, _03351_, _02934_);
  or (_03353_, _03352_, _03350_);
  or (_03354_, _03353_, _03349_);
  nor (_03355_, _03354_, _03348_);
  and (_03356_, _02904_, _02441_);
  nor (_03357_, _02983_, _03356_);
  or (_03358_, _03357_, _02539_);
  and (_03359_, _02522_, _02783_);
  and (_03360_, _03359_, _02798_);
  not (_03361_, _03360_);
  and (_03362_, _02907_, _02798_);
  and (_03363_, _02933_, _02784_);
  or (_03364_, _03363_, _02932_);
  nor (_03365_, _03364_, _03362_);
  and (_03366_, _03365_, _03361_);
  and (_03367_, _03366_, _03358_);
  and (_03368_, _03367_, _03355_);
  or (_03369_, _03368_, _03342_);
  nand (_03370_, _03369_, _02939_);
  and (_03371_, _02930_, \oc8051_golden_model_1.SP [0]);
  nor (_03372_, _03371_, _02800_);
  nand (_03373_, _03372_, _03370_);
  and (_03374_, _02971_, _02794_);
  not (_03375_, _03374_);
  nor (_03376_, _02914_, _02537_);
  nor (_03377_, _03376_, _03241_);
  and (_03378_, _03377_, _03375_);
  nor (_03379_, _03378_, _02519_);
  and (_03380_, _02907_, _02794_);
  nor (_03381_, _03380_, _02928_);
  not (_03382_, _03381_);
  nor (_03383_, _03382_, _03379_);
  nand (_03384_, _03383_, _03373_);
  nand (_03385_, _03384_, _03341_);
  and (_03386_, _03385_, _02927_);
  or (_03387_, _02797_, _03386_);
  and (_03388_, _02835_, _02795_);
  nor (_03389_, _02984_, _02944_);
  or (_03390_, _02907_, _03356_);
  nor (_03391_, _03390_, _03359_);
  or (_03392_, _03391_, _02532_);
  and (_03393_, _03392_, _03389_);
  not (_03394_, _03393_);
  nor (_03395_, _03394_, _03388_);
  and (_03396_, _03395_, _03387_);
  not (_03397_, _02944_);
  nor (_03398_, _03397_, _02835_);
  or (_03399_, _03398_, _03396_);
  nand (_03400_, _03399_, _02926_);
  nor (_03401_, _02926_, _03339_);
  nor (_03402_, _03401_, _02923_);
  nand (_03403_, _03402_, _03400_);
  and (_03404_, _02923_, _02835_);
  and (_03405_, _03359_, _02900_);
  not (_03406_, _03405_);
  and (_03407_, _03406_, _02903_);
  not (_03408_, _03407_);
  nor (_03409_, _03408_, _03404_);
  and (_03410_, _03409_, _03403_);
  or (_03411_, _03410_, _03340_);
  nor (_03412_, _02983_, _02523_);
  nor (_03413_, _03412_, _02498_);
  not (_03414_, _03413_);
  not (_03415_, _03268_);
  and (_03416_, _02905_, _02782_);
  not (_03417_, _03416_);
  and (_03418_, _03359_, _02782_);
  and (_03419_, _02919_, _02782_);
  nor (_03420_, _03419_, _03418_);
  and (_03421_, _03420_, _03417_);
  and (_03422_, _03421_, _03415_);
  and (_03423_, _03422_, _03414_);
  and (_03424_, _03423_, _03411_);
  nor (_03425_, _02899_, _02835_);
  or (_03426_, _03425_, _03424_);
  and (_03427_, _03426_, _02966_);
  or (_03428_, _03427_, _02786_);
  or (_03429_, _02983_, _02919_);
  and (_03430_, _03429_, _02347_);
  not (_03431_, _03430_);
  and (_03432_, _03359_, _02347_);
  not (_03433_, _03432_);
  not (_03434_, _03265_);
  and (_03435_, _02905_, _02347_);
  nor (_03436_, _03435_, _02524_);
  and (_03437_, _03436_, _03434_);
  and (_03438_, _03437_, _03433_);
  and (_03439_, _03438_, _03431_);
  and (_03440_, _03439_, _03428_);
  and (_03441_, _03046_, _01258_);
  and (_03442_, _03055_, _01271_);
  nor (_03443_, _03442_, _03441_);
  and (_03444_, _03075_, _01281_);
  and (_03445_, _03057_, _01245_);
  nor (_03446_, _03445_, _03444_);
  and (_03447_, _03446_, _03443_);
  and (_03448_, _03069_, _01251_);
  and (_03449_, _03034_, _01263_);
  nor (_03450_, _03449_, _03448_);
  and (_03451_, _03037_, _01249_);
  and (_03452_, _03063_, _01241_);
  nor (_03453_, _03452_, _03451_);
  and (_03454_, _03453_, _03450_);
  and (_03455_, _03454_, _03447_);
  and (_03456_, _03082_, _01274_);
  and (_03457_, _03052_, _01278_);
  nor (_03458_, _03457_, _03456_);
  and (_03459_, _03080_, _01256_);
  and (_03460_, _03077_, _01269_);
  nor (_03461_, _03460_, _03459_);
  and (_03462_, _03461_, _03458_);
  and (_03463_, _03066_, _01243_);
  and (_03464_, _03050_, _01276_);
  nor (_03465_, _03464_, _03463_);
  and (_03466_, _03071_, _01265_);
  and (_03467_, _03043_, _01253_);
  nor (_03468_, _03467_, _03466_);
  and (_03469_, _03468_, _03465_);
  and (_03470_, _03469_, _03462_);
  and (_03471_, _03470_, _03455_);
  nor (_03472_, _03471_, _02970_);
  or (_03473_, _03472_, _03440_);
  not (_03474_, _02894_);
  nor (_03475_, _03474_, _02775_);
  and (_03476_, _03359_, _02584_);
  nor (_03477_, _03476_, _02893_);
  not (_03478_, _03477_);
  nor (_03479_, _03478_, _03475_);
  and (_03480_, _03479_, _03473_);
  and (_03481_, _02893_, _02775_);
  or (_03482_, _03481_, _03480_);
  and (_03483_, _02905_, _02581_);
  and (_03484_, _02919_, _02581_);
  nor (_03485_, _03484_, _03483_);
  and (_03486_, _03359_, _02581_);
  not (_03487_, _03486_);
  and (_03488_, _02907_, _02581_);
  and (_03489_, _02983_, _02581_);
  nor (_03490_, _03489_, _03488_);
  and (_03491_, _03490_, _03487_);
  and (_03492_, _03491_, _03485_);
  and (_03493_, _03492_, _03482_);
  and (_03494_, _03329_, _02835_);
  and (_03495_, _02904_, _02472_);
  and (_03496_, _03495_, _02593_);
  and (_03497_, _03496_, _02441_);
  not (_03498_, _03497_);
  and (_03499_, _02971_, _02593_);
  and (_03500_, _03499_, _02441_);
  not (_03501_, _03500_);
  and (_03502_, _02906_, _02441_);
  and (_03503_, _03502_, _02593_);
  and (_03504_, _02905_, _02593_);
  nor (_03505_, _03504_, _03503_);
  and (_03506_, _03505_, _03501_);
  and (_03507_, _03506_, _03498_);
  not (_03508_, _03507_);
  nor (_03509_, _03508_, _03494_);
  and (_03510_, _03509_, _03493_);
  nor (_03511_, _03102_, _02836_);
  and (_03512_, _03359_, _02591_);
  and (_03513_, _02919_, _02591_);
  nor (_03514_, _03513_, _03512_);
  and (_03515_, _02907_, _02591_);
  nor (_03516_, _03515_, _03103_);
  and (_03517_, _02983_, _02591_);
  and (_03518_, _02905_, _02591_);
  nor (_03519_, _03518_, _03517_);
  and (_03520_, _03519_, _03516_);
  and (_03521_, _03520_, _03514_);
  and (_03522_, _03359_, _02588_);
  not (_03523_, _03522_);
  and (_03524_, _02919_, _02588_);
  not (_03525_, _03524_);
  and (_03526_, _02905_, _02588_);
  and (_03527_, _03502_, _02588_);
  nor (_03528_, _03527_, _03526_);
  and (_03529_, _03528_, _03525_);
  and (_03530_, _03529_, _03523_);
  and (_03531_, _03530_, _03521_);
  not (_03532_, _03531_);
  nor (_03533_, _03532_, _03511_);
  and (_03534_, _03533_, _03510_);
  nor (_03535_, _03104_, _02835_);
  nor (_03536_, _03535_, _03534_);
  and (_03537_, _03113_, _02787_);
  nor (_03538_, _03537_, _03536_);
  and (_03539_, _02905_, _02574_);
  nor (_03540_, _03539_, _03124_);
  and (_03541_, _03359_, _02574_);
  and (_03542_, _02919_, _02574_);
  nor (_03543_, _03542_, _03541_);
  nand (_03544_, _02906_, _02574_);
  or (_03545_, _03544_, _02519_);
  and (_03546_, _03545_, _03543_);
  and (_03547_, _03546_, _03540_);
  not (_03548_, _03547_);
  not (_03549_, _02993_);
  nor (_03550_, _03549_, _02775_);
  nor (_03551_, _03550_, _03548_);
  and (_03552_, _03551_, _03538_);
  nor (_03553_, _02857_, _02835_);
  nor (_03554_, _03553_, _03552_);
  and (_03555_, _02854_, _02787_);
  nor (_03556_, _03555_, _03554_);
  and (_03557_, _02919_, _02571_);
  nor (_03558_, _03557_, _03133_);
  and (_03559_, _03359_, _02571_);
  not (_03560_, _03559_);
  and (_03561_, _02983_, _02571_);
  not (_03562_, _02571_);
  nor (_03563_, _02908_, _03562_);
  nor (_03564_, _03563_, _03561_);
  and (_03565_, _03564_, _03560_);
  and (_03566_, _03565_, _03558_);
  not (_03567_, _03566_);
  nor (_03568_, _03134_, _02775_);
  nor (_03569_, _03568_, _03567_);
  and (_03570_, _03569_, _03556_);
  nor (_03571_, _03138_, _02835_);
  or (_03572_, _03571_, _03570_);
  and (_03573_, _03572_, _03142_);
  or (_03574_, _02779_, _03573_);
  not (_03575_, _02567_);
  nor (_03576_, _02908_, _03575_);
  not (_03577_, _03576_);
  and (_03578_, _02983_, _02567_);
  and (_03579_, _03359_, _02567_);
  nor (_03580_, _03579_, _03578_);
  and (_03581_, _02919_, _02567_);
  nor (_03582_, _03581_, _02852_);
  and (_03583_, _03582_, _03580_);
  and (_03584_, _03583_, _03577_);
  nand (_03585_, _03584_, _03574_);
  nor (_03586_, _02853_, _02835_);
  not (_03587_, _03586_);
  nand (_03588_, _03587_, _03585_);
  or (_03589_, _03588_, _03338_);
  nor (_03590_, _02687_, _33770_);
  nor (_03591_, _02710_, _33483_);
  nor (_03592_, _03591_, _03590_);
  nor (_03593_, _02727_, _33319_);
  nor (_03594_, _02703_, _33196_);
  nor (_03595_, _03594_, _03593_);
  and (_03596_, _03595_, _03592_);
  nor (_03597_, _02698_, _33442_);
  nor (_03598_, _02720_, _33360_);
  nor (_03599_, _03598_, _03597_);
  nor (_03600_, _02731_, _33688_);
  nor (_03601_, _02715_, _33647_);
  nor (_03602_, _03601_, _03600_);
  and (_03603_, _03602_, _03599_);
  and (_03604_, _03603_, _03596_);
  nor (_03605_, _02693_, _33565_);
  nor (_03606_, _02707_, _33524_);
  nor (_03607_, _03606_, _03605_);
  nor (_03608_, _02722_, _33278_);
  nor (_03609_, _02736_, _33155_);
  nor (_03610_, _03609_, _03608_);
  and (_03611_, _03610_, _03607_);
  nor (_03612_, _02713_, _33729_);
  nor (_03613_, _02725_, _33401_);
  nor (_03614_, _03613_, _03612_);
  nor (_03615_, _02733_, _33606_);
  nor (_03616_, _02738_, _33237_);
  nor (_03617_, _03616_, _03615_);
  and (_03618_, _03617_, _03614_);
  and (_03619_, _03618_, _03611_);
  and (_03620_, _03619_, _03604_);
  nor (_03621_, _03620_, _02858_);
  and (_03622_, _03182_, _03183_);
  and (_03623_, _03622_, _03188_);
  and (_03624_, _03623_, _03187_);
  not (_03625_, _03624_);
  and (_03626_, _03625_, _03621_);
  not (_03627_, _03626_);
  and (_03628_, _03621_, _02785_);
  not (_03629_, _03628_);
  and (_03630_, _03080_, _01318_);
  and (_03631_, _03043_, _01292_);
  nor (_03632_, _03631_, _03630_);
  and (_03633_, _03052_, _01298_);
  and (_03634_, _03057_, _01306_);
  nor (_03635_, _03634_, _03633_);
  and (_03636_, _03635_, _03632_);
  and (_03637_, _03069_, _01324_);
  and (_03638_, _03046_, _01308_);
  nor (_03639_, _03638_, _03637_);
  and (_03640_, _03034_, _01315_);
  and (_03641_, _03082_, _01289_);
  nor (_03642_, _03641_, _03640_);
  and (_03643_, _03642_, _03639_);
  and (_03644_, _03643_, _03636_);
  and (_03645_, _03050_, _01300_);
  and (_03646_, _03075_, _01303_);
  nor (_03647_, _03646_, _03645_);
  and (_03648_, _03063_, _01287_);
  and (_03649_, _03077_, _01326_);
  nor (_03650_, _03649_, _03648_);
  and (_03651_, _03650_, _03647_);
  and (_03652_, _03037_, _01313_);
  and (_03653_, _03055_, _01328_);
  nor (_03654_, _03653_, _03652_);
  and (_03655_, _03071_, _01320_);
  and (_03656_, _03066_, _01294_);
  nor (_03657_, _03656_, _03655_);
  and (_03658_, _03657_, _03654_);
  and (_03659_, _03658_, _03651_);
  and (_03660_, _03659_, _03644_);
  nor (_03661_, _03660_, _02970_);
  not (_03662_, _02581_);
  not (_03663_, _02347_);
  and (_03664_, _02539_, _03663_);
  and (_03665_, _03664_, _03662_);
  nor (_03666_, _03665_, _02441_);
  not (_03667_, _03666_);
  and (_03668_, _02532_, _02498_);
  nor (_03669_, _02593_, _02794_);
  nor (_03670_, _02567_, _02588_);
  and (_03671_, _03670_, _03669_);
  and (_03672_, _03671_, _03668_);
  and (_03673_, _03672_, _03667_);
  nor (_03674_, _03673_, _02914_);
  nor (_03675_, _03344_, _03242_);
  not (_03676_, _03675_);
  nor (_03677_, _03676_, _03674_);
  nor (_03678_, _03677_, _02472_);
  nor (_03679_, _03246_, _03241_);
  and (_03680_, _02904_, _02515_);
  and (_03681_, _03680_, _02591_);
  nor (_03682_, _03681_, _03483_);
  and (_03683_, _03682_, _03679_);
  and (_03684_, _03683_, _03261_);
  not (_03685_, _02905_);
  nor (_03686_, _02574_, _02933_);
  and (_03687_, _03686_, _03664_);
  nor (_03688_, _03687_, _03685_);
  not (_03689_, _03688_);
  and (_03690_, _03689_, _03238_);
  and (_03691_, _03690_, _03684_);
  not (_03692_, \oc8051_golden_model_1.SP [1]);
  not (_03693_, _02930_);
  nor (_03694_, _03113_, _02854_);
  and (_03695_, _03694_, _03693_);
  nor (_03696_, _03695_, _03692_);
  not (_03697_, _03696_);
  and (_03698_, _03231_, _02567_);
  and (_03699_, _03680_, _02571_);
  nor (_03700_, _03699_, _03698_);
  and (_03701_, _03700_, _03279_);
  and (_03702_, _03011_, _02574_);
  and (_03703_, _03011_, _02933_);
  nor (_03704_, _03703_, _03702_);
  and (_03705_, _03704_, _03701_);
  and (_03706_, _03705_, _03697_);
  and (_03707_, _03706_, _03691_);
  not (_03708_, _03707_);
  nor (_03709_, _03708_, _03678_);
  not (_03710_, _03709_);
  nor (_03711_, _03710_, _03661_);
  nor (_03712_, _02687_, _33755_);
  nor (_03713_, _02710_, _33468_);
  nor (_03714_, _03713_, _03712_);
  nor (_03715_, _02693_, _33550_);
  nor (_03716_, _02736_, _33140_);
  nor (_03717_, _03716_, _03715_);
  and (_03718_, _03717_, _03714_);
  nor (_03719_, _02698_, _33427_);
  nor (_03720_, _02720_, _33345_);
  nor (_03721_, _03720_, _03719_);
  nor (_03722_, _02731_, _33673_);
  nor (_03723_, _02715_, _33632_);
  nor (_03724_, _03723_, _03722_);
  and (_03725_, _03724_, _03721_);
  and (_03726_, _03725_, _03718_);
  nor (_03727_, _02727_, _33304_);
  nor (_03728_, _02738_, _33222_);
  nor (_03729_, _03728_, _03727_);
  nor (_03730_, _02722_, _33263_);
  nor (_03731_, _02703_, _33181_);
  nor (_03732_, _03731_, _03730_);
  and (_03733_, _03732_, _03729_);
  nor (_03734_, _02713_, _33714_);
  nor (_03735_, _02725_, _33386_);
  nor (_03736_, _03735_, _03734_);
  nor (_03737_, _02733_, _33591_);
  nor (_03738_, _02707_, _33509_);
  nor (_03739_, _03738_, _03737_);
  and (_03740_, _03739_, _03736_);
  and (_03741_, _03740_, _03733_);
  and (_03742_, _03741_, _03726_);
  not (_03743_, _03742_);
  and (_03744_, _03743_, _03333_);
  not (_03745_, _03744_);
  and (_03746_, _03745_, _03711_);
  and (_03747_, _03746_, _03629_);
  and (_03748_, _03747_, _03627_);
  nand (_03749_, _03588_, \oc8051_golden_model_1.IRAM[1] [0]);
  and (_03750_, _03749_, _03748_);
  nand (_03751_, _03750_, _03589_);
  not (_03752_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_03753_, _03587_, _03585_);
  or (_03754_, _03753_, _03752_);
  not (_03755_, _03748_);
  nand (_03756_, _03753_, \oc8051_golden_model_1.IRAM[2] [0]);
  and (_03757_, _03756_, _03755_);
  nand (_03758_, _03757_, _03754_);
  nand (_03759_, _03758_, _03751_);
  nand (_03760_, _03759_, _03337_);
  not (_03761_, _03337_);
  not (_03762_, \oc8051_golden_model_1.IRAM[7] [0]);
  or (_03763_, _03753_, _03762_);
  not (_03764_, \oc8051_golden_model_1.IRAM[6] [0]);
  or (_03765_, _03588_, _03764_);
  and (_03766_, _03765_, _03755_);
  nand (_03767_, _03766_, _03763_);
  not (_03768_, \oc8051_golden_model_1.IRAM[4] [0]);
  or (_03769_, _03588_, _03768_);
  not (_03770_, \oc8051_golden_model_1.IRAM[5] [0]);
  or (_03771_, _03753_, _03770_);
  and (_03772_, _03771_, _03748_);
  nand (_03773_, _03772_, _03769_);
  nand (_03774_, _03773_, _03767_);
  nand (_03775_, _03774_, _03761_);
  nand (_03776_, _03775_, _03760_);
  nand (_03777_, _03776_, _03148_);
  not (_03778_, _03148_);
  not (_03779_, \oc8051_golden_model_1.IRAM[11] [0]);
  or (_03780_, _03753_, _03779_);
  nand (_03781_, _03753_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_03782_, _03781_, _03755_);
  nand (_03783_, _03782_, _03780_);
  not (_03784_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_03785_, _03588_, _03784_);
  nand (_03786_, _03588_, \oc8051_golden_model_1.IRAM[9] [0]);
  and (_03787_, _03786_, _03748_);
  nand (_03788_, _03787_, _03785_);
  nand (_03789_, _03788_, _03783_);
  nand (_03790_, _03789_, _03337_);
  not (_03791_, \oc8051_golden_model_1.IRAM[15] [0]);
  or (_03792_, _03753_, _03791_);
  nand (_03793_, _03753_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_03794_, _03793_, _03755_);
  nand (_03795_, _03794_, _03792_);
  not (_03796_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_03797_, _03588_, _03796_);
  nand (_03798_, _03588_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_03799_, _03798_, _03748_);
  nand (_03800_, _03799_, _03797_);
  nand (_03801_, _03800_, _03795_);
  nand (_03802_, _03801_, _03761_);
  nand (_03803_, _03802_, _03790_);
  nand (_03804_, _03803_, _03778_);
  and (_03805_, _03804_, _03777_);
  and (_03806_, _02971_, _02798_);
  nor (_03807_, _03806_, _03345_);
  nor (_03808_, _03807_, _03805_);
  nor (_03809_, _03808_, _02851_);
  and (_03810_, _02799_, _02743_);
  and (_03811_, _02932_, _02743_);
  and (_03812_, _03811_, _02835_);
  nor (_03813_, _03812_, _03810_);
  and (_03814_, _03813_, _03809_);
  nor (_03815_, _03814_, _02800_);
  nor (_03816_, _02540_, _02787_);
  nor (_03817_, _03816_, _03815_);
  and (_03818_, _02930_, _02743_);
  and (_03819_, _03818_, _02835_);
  and (_03820_, _02841_, _02794_);
  nor (_03821_, _03820_, _03819_);
  and (_03822_, _03821_, _03817_);
  nand (_03823_, _03804_, _03777_);
  and (_03824_, _03823_, _03374_);
  not (_03825_, _03824_);
  and (_03826_, _03825_, _03822_);
  and (_03827_, _02796_, _02743_);
  and (_03828_, _02928_, _02743_);
  and (_03829_, _03828_, _02835_);
  nor (_03830_, _03829_, _03827_);
  and (_03831_, _03830_, _03826_);
  nor (_03832_, _03831_, _02797_);
  or (_03833_, _03832_, _02795_);
  nand (_03834_, _02795_, _02787_);
  nand (_03835_, _03834_, _03833_);
  and (_03836_, _03835_, _02793_);
  nor (_03837_, _03836_, _02791_);
  and (_03838_, _02841_, _02900_);
  or (_03839_, _03838_, _03837_);
  nor (_03840_, _03839_, _02788_);
  and (_03841_, _02743_, _02785_);
  and (_03842_, _02971_, _02900_);
  and (_03843_, _03823_, _03842_);
  nor (_03844_, _03843_, _03841_);
  and (_03845_, _03844_, _03840_);
  nor (_03846_, _03845_, _02786_);
  nor (_03847_, _03846_, _02518_);
  and (_03848_, _02518_, _02787_);
  nor (_03849_, _03848_, _03847_);
  and (_03850_, _02971_, _02347_);
  and (_03851_, _03850_, _02743_);
  not (_03852_, _03851_);
  and (_03853_, _02743_, _02524_);
  or (_03854_, _03282_, _03246_);
  nor (_03855_, _03012_, _03663_);
  nor (_03856_, _03855_, _03854_);
  and (_03857_, _02904_, _02473_);
  and (_03858_, _03857_, _02347_);
  not (_03859_, _03858_);
  and (_03860_, _03859_, _03856_);
  not (_03861_, _03860_);
  and (_03862_, _03861_, _02743_);
  nor (_03863_, _03862_, _03853_);
  and (_03864_, _03863_, _03852_);
  nor (_03865_, _03864_, _02836_);
  and (_03866_, _02841_, _02584_);
  nor (_03867_, _03866_, _03865_);
  not (_03868_, _03867_);
  nor (_03869_, _03868_, _03849_);
  and (_03870_, _02971_, _02584_);
  and (_03871_, _03823_, _03870_);
  not (_03872_, _03871_);
  and (_03873_, _03872_, _03869_);
  and (_03874_, _02974_, _02743_);
  and (_03875_, _03874_, _02835_);
  nor (_03876_, _03875_, _02585_);
  and (_03877_, _03876_, _03873_);
  and (_03878_, _02585_, _02787_);
  nor (_03879_, _03878_, _03877_);
  and (_03880_, _03094_, _02743_);
  not (_03881_, _02991_);
  and (_03882_, _03108_, _03881_);
  nor (_03883_, _03882_, _02858_);
  nor (_03884_, _03883_, _03880_);
  nor (_03885_, _03884_, _02836_);
  nor (_03886_, _03885_, _02594_);
  not (_03887_, _03886_);
  nor (_03888_, _03887_, _03879_);
  and (_03889_, _02594_, _02787_);
  nor (_03890_, _03889_, _03888_);
  nor (_03891_, _03100_, _02858_);
  and (_03892_, _03891_, _02835_);
  nor (_03893_, _03892_, _02592_);
  not (_03894_, _03893_);
  nor (_03895_, _03894_, _03890_);
  and (_03896_, _02592_, _02787_);
  nor (_03897_, _03896_, _03895_);
  and (_03898_, _02971_, _02571_);
  and (_03899_, _03823_, _03898_);
  and (_03900_, _03133_, _02743_);
  and (_03901_, _02841_, _02571_);
  or (_03902_, _03901_, _03900_);
  or (_03903_, _03902_, _03899_);
  nor (_03904_, _03903_, _03897_);
  and (_03905_, _03900_, _02836_);
  nor (_03906_, _03905_, _03904_);
  nor (_03907_, _02988_, _02572_);
  nor (_03908_, _03907_, _02787_);
  nor (_03909_, _03908_, _03906_);
  and (_03910_, _03909_, _02781_);
  nor (_03911_, _03910_, _02779_);
  and (_03912_, _02971_, _02567_);
  and (_03913_, _03823_, _03912_);
  and (_03914_, _02852_, _02743_);
  and (_03915_, _02841_, _02567_);
  or (_03916_, _03915_, _03914_);
  or (_03917_, _03916_, _03913_);
  nor (_03918_, _03917_, _03911_);
  and (_03919_, _03914_, _02836_);
  nor (_03920_, _03919_, _03918_);
  not (_03921_, _03920_);
  and (_03922_, _03914_, _03743_);
  and (_03923_, _03621_, _02778_);
  and (_03924_, _03692_, \oc8051_golden_model_1.SP [0]);
  and (_03925_, \oc8051_golden_model_1.SP [1], _02787_);
  nor (_03926_, _03925_, _03924_);
  not (_03927_, _03926_);
  and (_03928_, _03927_, _02592_);
  and (_03929_, _03874_, _03743_);
  nor (_03930_, _03864_, _03743_);
  and (_03931_, _03927_, _02795_);
  not (_03932_, _02795_);
  not (_03933_, \oc8051_golden_model_1.IRAM[0] [1]);
  or (_03934_, _03588_, _03933_);
  nand (_03935_, _03588_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_03936_, _03935_, _03748_);
  nand (_03937_, _03936_, _03934_);
  not (_03938_, \oc8051_golden_model_1.IRAM[3] [1]);
  or (_03939_, _03753_, _03938_);
  nand (_03940_, _03753_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_03941_, _03940_, _03755_);
  nand (_03942_, _03941_, _03939_);
  nand (_03943_, _03942_, _03937_);
  nand (_03944_, _03943_, _03337_);
  not (_03945_, \oc8051_golden_model_1.IRAM[7] [1]);
  or (_03946_, _03753_, _03945_);
  not (_03947_, \oc8051_golden_model_1.IRAM[6] [1]);
  or (_03948_, _03588_, _03947_);
  and (_03949_, _03948_, _03755_);
  nand (_03950_, _03949_, _03946_);
  not (_03951_, \oc8051_golden_model_1.IRAM[4] [1]);
  or (_03952_, _03588_, _03951_);
  not (_03953_, \oc8051_golden_model_1.IRAM[5] [1]);
  or (_03954_, _03753_, _03953_);
  and (_03955_, _03954_, _03748_);
  nand (_03956_, _03955_, _03952_);
  nand (_03957_, _03956_, _03950_);
  nand (_03958_, _03957_, _03761_);
  nand (_03959_, _03958_, _03944_);
  nand (_03960_, _03959_, _03148_);
  not (_03961_, \oc8051_golden_model_1.IRAM[11] [1]);
  or (_03962_, _03753_, _03961_);
  nand (_03963_, _03753_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_03964_, _03963_, _03755_);
  nand (_03965_, _03964_, _03962_);
  not (_03966_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_03967_, _03588_, _03966_);
  nand (_03968_, _03588_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_03969_, _03968_, _03748_);
  nand (_03970_, _03969_, _03967_);
  nand (_03971_, _03970_, _03965_);
  nand (_03972_, _03971_, _03337_);
  not (_03973_, \oc8051_golden_model_1.IRAM[15] [1]);
  or (_03974_, _03753_, _03973_);
  not (_03975_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_03976_, _03588_, _03975_);
  and (_03977_, _03976_, _03755_);
  nand (_03978_, _03977_, _03974_);
  not (_03979_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_03980_, _03588_, _03979_);
  not (_03981_, \oc8051_golden_model_1.IRAM[13] [1]);
  or (_03982_, _03753_, _03981_);
  and (_03983_, _03982_, _03748_);
  nand (_03984_, _03983_, _03980_);
  nand (_03985_, _03984_, _03978_);
  nand (_03986_, _03985_, _03761_);
  nand (_03987_, _03986_, _03972_);
  nand (_03988_, _03987_, _03778_);
  nand (_03989_, _03988_, _03960_);
  not (_03990_, _03989_);
  or (_03991_, _03990_, _03807_);
  not (_03992_, _03811_);
  and (_03993_, _02472_, _02409_);
  and (_03994_, _03993_, _02803_);
  nor (_03995_, _03994_, _02838_);
  and (_03996_, _03743_, _02838_);
  or (_03997_, _03996_, _02804_);
  or (_03998_, _03997_, _03995_);
  and (_03999_, _03926_, _02804_);
  and (_04000_, _03993_, _02798_);
  nor (_04001_, _04000_, _03999_);
  and (_04002_, _04001_, _03998_);
  and (_04003_, _04002_, _03992_);
  and (_04004_, _04003_, _03991_);
  and (_04005_, _03811_, _03743_);
  nor (_04006_, _04005_, _04004_);
  and (_04007_, _03620_, _03810_);
  nor (_04008_, _04007_, _04006_);
  or (_04009_, _03927_, _02540_);
  nand (_04010_, _04009_, _04008_);
  and (_04011_, _03818_, _03742_);
  and (_04012_, _03993_, _02794_);
  nor (_04013_, _04012_, _04011_);
  not (_04014_, _04013_);
  nor (_04015_, _04014_, _04010_);
  and (_04016_, _03989_, _03374_);
  nor (_04017_, _04016_, _03828_);
  and (_04018_, _04017_, _04015_);
  and (_04019_, _03828_, _03743_);
  nor (_04020_, _04019_, _04018_);
  and (_04021_, _03620_, _03827_);
  nor (_04022_, _04021_, _04020_);
  and (_04023_, _04022_, _03932_);
  nor (_04024_, _04023_, _03931_);
  and (_04025_, _03620_, _02792_);
  or (_04026_, _04025_, _04024_);
  nor (_04027_, _03927_, _02533_);
  and (_04028_, _03993_, _02900_);
  nor (_04029_, _04028_, _04027_);
  not (_04030_, _04029_);
  nor (_04031_, _04030_, _04026_);
  and (_04032_, _03989_, _03842_);
  nor (_04033_, _04032_, _03841_);
  and (_04034_, _04033_, _04031_);
  nor (_04035_, _04034_, _03628_);
  nor (_04036_, _04035_, _02518_);
  and (_04037_, _03927_, _02518_);
  nor (_04038_, _04037_, _04036_);
  and (_04039_, _03993_, _02584_);
  or (_04040_, _04039_, _04038_);
  nor (_04041_, _04040_, _03930_);
  and (_04042_, _03989_, _03870_);
  nor (_04043_, _04042_, _03874_);
  and (_04044_, _04043_, _04041_);
  nor (_04045_, _04044_, _03929_);
  nor (_04046_, _04045_, _02585_);
  and (_04047_, _03927_, _02585_);
  nor (_04048_, _04047_, _04046_);
  nor (_04049_, _03884_, _03743_);
  nor (_04050_, _04049_, _02594_);
  not (_04051_, _04050_);
  nor (_04052_, _04051_, _04048_);
  and (_04053_, _03927_, _02594_);
  nor (_04054_, _04053_, _04052_);
  and (_04055_, _03891_, _03742_);
  nor (_04056_, _04055_, _02592_);
  not (_04057_, _04056_);
  nor (_04058_, _04057_, _04054_);
  nor (_04059_, _04058_, _03928_);
  and (_04060_, _03495_, _02571_);
  not (_04061_, _04060_);
  nand (_04062_, _04061_, _03230_);
  nor (_04063_, _04062_, _04059_);
  and (_04064_, _03989_, _03898_);
  nor (_04065_, _04064_, _03900_);
  and (_04066_, _04065_, _04063_);
  and (_04067_, _03900_, _03743_);
  nor (_04068_, _04067_, _04066_);
  nor (_04069_, _03927_, _03907_);
  nor (_04070_, _04069_, _02780_);
  not (_04071_, _04070_);
  nor (_04072_, _04071_, _04068_);
  nor (_04073_, _04072_, _03923_);
  and (_04074_, _03993_, _02567_);
  nor (_04075_, _04074_, _04073_);
  and (_04076_, _03989_, _03912_);
  nor (_04077_, _04076_, _03914_);
  and (_04078_, _04077_, _04075_);
  nor (_04079_, _04078_, _03922_);
  not (_04080_, _00000_);
  nor (_04081_, _03828_, _03818_);
  nor (_04082_, _03811_, _03810_);
  and (_04083_, _04082_, _04081_);
  nor (_04084_, _03874_, _03827_);
  and (_04085_, _03244_, _02584_);
  not (_04086_, _04085_);
  and (_04087_, _02919_, _02798_);
  and (_04088_, _03011_, _02900_);
  nor (_04089_, _04088_, _04087_);
  and (_04090_, _04089_, _04086_);
  and (_04091_, _03011_, _02584_);
  and (_04092_, _03376_, _02776_);
  nor (_04093_, _04092_, _04091_);
  and (_04094_, _03231_, _02584_);
  not (_04095_, _04094_);
  and (_04096_, _04095_, _04093_);
  not (_04097_, _03579_);
  and (_04098_, _03700_, _04097_);
  and (_04099_, _02904_, _02584_);
  and (_04100_, _04099_, _02776_);
  and (_04101_, _03912_, _02519_);
  nor (_04102_, _04101_, _04100_);
  and (_04103_, _04102_, _04098_);
  and (_04104_, _04103_, _04096_);
  and (_04105_, _04104_, _04090_);
  and (_04106_, _03009_, _02584_);
  not (_04107_, _04106_);
  and (_04108_, _02912_, _02571_);
  nor (_04109_, _04108_, _03228_);
  and (_04110_, _04109_, _04107_);
  and (_04111_, _03011_, _02567_);
  and (_04112_, _03244_, _02567_);
  nor (_04113_, _04112_, _04111_);
  and (_04114_, _02915_, _02472_);
  nor (_04115_, _04114_, _03842_);
  and (_04116_, _04115_, _04113_);
  and (_04117_, _04116_, _04110_);
  and (_04118_, _02906_, _02803_);
  not (_04119_, _04118_);
  and (_04120_, _02904_, _02911_);
  and (_04121_, _04120_, _02798_);
  and (_04122_, _02904_, _02803_);
  nor (_04123_, _04122_, _04121_);
  and (_04124_, _04123_, _04119_);
  and (_04125_, _03857_, _02567_);
  nor (_04126_, _04125_, _03374_);
  and (_04127_, _04120_, _02794_);
  nor (_04128_, _04127_, _04060_);
  and (_04129_, _04128_, _04126_);
  and (_04130_, _04129_, _04124_);
  not (_04131_, _02585_);
  not (_04132_, _02518_);
  and (_04133_, _02533_, _04132_);
  and (_04134_, _04133_, _04131_);
  and (_04135_, _04134_, _02910_);
  and (_04136_, _04135_, _04130_);
  and (_04137_, _03907_, _02595_);
  and (_04138_, _02546_, _02540_);
  and (_04139_, _03276_, _04138_);
  and (_04140_, _04139_, _04137_);
  nor (_04141_, _03277_, _03241_);
  and (_04142_, _04141_, _03807_);
  nor (_04143_, _03898_, _03870_);
  nor (_04144_, _02913_, _02795_);
  and (_04145_, _04144_, _04143_);
  and (_04146_, _04145_, _04142_);
  and (_04147_, _04146_, _04140_);
  and (_04148_, _04147_, _04136_);
  and (_04149_, _04148_, _04117_);
  and (_04150_, _04149_, _04105_);
  not (_04151_, _04150_);
  nor (_04152_, _04151_, _03891_);
  and (_04153_, _04152_, _04084_);
  and (_04154_, _04153_, _04083_);
  nor (_04155_, _03914_, _02780_);
  not (_04156_, _03855_);
  not (_04157_, _03854_);
  and (_04158_, _03495_, _02347_);
  nor (_04159_, _04158_, _02837_);
  and (_04160_, _04159_, _04157_);
  nor (_04161_, _03850_, _03094_);
  and (_04162_, _04161_, _03436_);
  and (_04163_, _04162_, _04160_);
  and (_04164_, _04163_, _04156_);
  nor (_04165_, _04164_, _02858_);
  not (_04166_, _04165_);
  and (_04167_, _04166_, _04155_);
  nor (_04168_, _03841_, _02792_);
  nor (_04169_, _03900_, _03883_);
  and (_04170_, _04169_, _04168_);
  and (_04171_, _04170_, _04167_);
  and (_04172_, _04171_, _04154_);
  nor (_04173_, _04172_, _04080_);
  not (_04174_, _04173_);
  nor (_04175_, _04174_, _04079_);
  and (_04176_, _04175_, _03921_);
  nand (_04177_, _03753_, \oc8051_golden_model_1.IRAM[0] [3]);
  nand (_04178_, _03588_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_04179_, _04178_, _03748_);
  nand (_04180_, _04179_, _04177_);
  nand (_04181_, _03588_, \oc8051_golden_model_1.IRAM[3] [3]);
  nand (_04182_, _03753_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_04183_, _04182_, _03755_);
  nand (_04184_, _04183_, _04181_);
  nand (_04185_, _04184_, _04180_);
  nand (_04186_, _04185_, _03337_);
  not (_04187_, \oc8051_golden_model_1.IRAM[7] [3]);
  or (_04188_, _03753_, _04187_);
  not (_04189_, \oc8051_golden_model_1.IRAM[6] [3]);
  or (_04190_, _03588_, _04189_);
  and (_04191_, _04190_, _03755_);
  nand (_04192_, _04191_, _04188_);
  not (_04193_, \oc8051_golden_model_1.IRAM[4] [3]);
  or (_04194_, _03588_, _04193_);
  not (_04195_, \oc8051_golden_model_1.IRAM[5] [3]);
  or (_04196_, _03753_, _04195_);
  and (_04197_, _04196_, _03748_);
  nand (_04198_, _04197_, _04194_);
  nand (_04199_, _04198_, _04192_);
  nand (_04200_, _04199_, _03761_);
  nand (_04201_, _04200_, _04186_);
  nand (_04202_, _04201_, _03148_);
  nand (_04203_, _03588_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_04204_, _03753_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_04205_, _04204_, _03755_);
  nand (_04206_, _04205_, _04203_);
  nand (_04207_, _03753_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand (_04208_, _03588_, \oc8051_golden_model_1.IRAM[9] [3]);
  and (_04209_, _04208_, _03748_);
  nand (_04210_, _04209_, _04207_);
  nand (_04211_, _04210_, _04206_);
  nand (_04212_, _04211_, _03337_);
  nand (_04213_, _03588_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_04214_, _03753_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_04215_, _04214_, _03755_);
  nand (_04216_, _04215_, _04213_);
  not (_04217_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_04218_, _03588_, _04217_);
  nand (_04219_, _03588_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_04220_, _04219_, _03748_);
  nand (_04221_, _04220_, _04218_);
  nand (_04222_, _04221_, _04216_);
  nand (_04223_, _04222_, _03761_);
  nand (_04224_, _04223_, _04212_);
  nand (_04225_, _04224_, _03778_);
  nand (_04226_, _04225_, _04202_);
  and (_04227_, _04226_, _03912_);
  and (_04228_, _02974_, _02775_);
  and (_04229_, _04226_, _03870_);
  not (_04230_, _02533_);
  and (_04231_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_04232_, _04231_, \oc8051_golden_model_1.SP [2]);
  or (_04233_, _04232_, \oc8051_golden_model_1.SP [3]);
  and (_04234_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_04235_, _04234_, \oc8051_golden_model_1.SP [3]);
  nand (_04236_, _04235_, \oc8051_golden_model_1.SP [0]);
  and (_04237_, _04236_, _04233_);
  and (_04238_, _04237_, _04230_);
  not (_04239_, _02540_);
  and (_04240_, _03810_, _02889_);
  and (_04241_, _04226_, _03806_);
  and (_04242_, _04237_, _02804_);
  and (_04243_, _04226_, _03345_);
  nor (_04244_, _03345_, \oc8051_golden_model_1.PSW [3]);
  nor (_04245_, _04244_, _02838_);
  not (_04246_, _04245_);
  nor (_04247_, _04246_, _04243_);
  and (_04248_, _02837_, _02775_);
  nor (_04249_, _04248_, _04247_);
  nor (_04250_, _04249_, _02804_);
  or (_04251_, _04250_, _03806_);
  nor (_04252_, _04251_, _04242_);
  or (_04253_, _04252_, _03811_);
  nor (_04254_, _04253_, _04241_);
  and (_04255_, _03811_, _02774_);
  or (_04256_, _04255_, _03810_);
  nor (_04257_, _04256_, _04254_);
  nor (_04258_, _04257_, _04240_);
  nor (_04259_, _04258_, _04239_);
  nor (_04260_, _04237_, _02540_);
  nor (_04261_, _04260_, _03818_);
  not (_04262_, _04261_);
  nor (_04263_, _04262_, _04259_);
  and (_04264_, _03818_, _02774_);
  or (_04265_, _04264_, _03374_);
  nor (_04266_, _04265_, _04263_);
  and (_04267_, _04226_, _03374_);
  nor (_04268_, _04267_, _03828_);
  not (_04269_, _04268_);
  nor (_04270_, _04269_, _04266_);
  and (_04271_, _02928_, _02775_);
  or (_04272_, _04271_, _03827_);
  nor (_04273_, _04272_, _04270_);
  and (_04274_, _02889_, _03827_);
  nor (_04275_, _04274_, _04273_);
  and (_04276_, _04275_, _03932_);
  and (_04277_, _04237_, _02795_);
  nor (_04278_, _04277_, _04276_);
  nor (_04279_, _04278_, _02792_);
  nor (_04280_, _02793_, _02892_);
  or (_04281_, _04280_, _04279_);
  and (_04282_, _04281_, _02533_);
  or (_04283_, _04282_, _03842_);
  nor (_04284_, _04283_, _04238_);
  and (_04285_, _04226_, _03842_);
  nor (_04286_, _04285_, _03841_);
  not (_04287_, _04286_);
  nor (_04288_, _04287_, _04284_);
  not (_04289_, _03841_);
  nor (_04290_, _04289_, _02892_);
  nor (_04291_, _04290_, _04288_);
  nor (_04292_, _04291_, _02518_);
  and (_04293_, _04237_, _02518_);
  not (_04294_, _04293_);
  and (_04295_, _04294_, _03864_);
  not (_04296_, _04295_);
  nor (_04297_, _04296_, _04292_);
  nor (_04298_, _03864_, _02774_);
  nor (_04299_, _04298_, _04297_);
  nor (_04300_, _04299_, _03870_);
  or (_04301_, _04300_, _03874_);
  nor (_04302_, _04301_, _04229_);
  nor (_04303_, _04302_, _04228_);
  nor (_04304_, _04303_, _02585_);
  and (_04305_, _04237_, _02585_);
  not (_04306_, _04305_);
  and (_04307_, _04306_, _03884_);
  not (_04308_, _04307_);
  nor (_04309_, _04308_, _04304_);
  nor (_04310_, _03884_, _02774_);
  nor (_04311_, _04310_, _02594_);
  not (_04312_, _04311_);
  nor (_04313_, _04312_, _04309_);
  and (_04314_, _04237_, _02594_);
  nor (_04315_, _04314_, _03891_);
  not (_04316_, _04315_);
  nor (_04317_, _04316_, _04313_);
  not (_04318_, _02774_);
  and (_04319_, _03891_, _04318_);
  nor (_04320_, _04319_, _02592_);
  not (_04321_, _04320_);
  nor (_04322_, _04321_, _04317_);
  and (_04323_, _04237_, _02592_);
  nor (_04324_, _04323_, _03898_);
  not (_04325_, _04324_);
  nor (_04326_, _04325_, _04322_);
  and (_04327_, _04226_, _03898_);
  nor (_04328_, _04327_, _03900_);
  not (_04329_, _04328_);
  nor (_04330_, _04329_, _04326_);
  not (_04331_, _03907_);
  and (_04332_, _03133_, _02775_);
  nor (_04333_, _04332_, _04331_);
  not (_04334_, _04333_);
  nor (_04335_, _04334_, _04330_);
  nor (_04336_, _04237_, _03907_);
  nor (_04337_, _04336_, _02780_);
  not (_04338_, _04337_);
  nor (_04339_, _04338_, _04335_);
  not (_04340_, _02889_);
  and (_04341_, _02780_, _04340_);
  nor (_04342_, _04341_, _03912_);
  not (_04343_, _04342_);
  nor (_04344_, _04343_, _04339_);
  or (_04345_, _04344_, _03914_);
  nor (_04346_, _04345_, _04227_);
  and (_04347_, _03914_, _02774_);
  nor (_04348_, _04347_, _04346_);
  and (_04349_, _02904_, _02567_);
  and (_04350_, _03180_, _02778_);
  nor (_04351_, _04231_, \oc8051_golden_model_1.SP [2]);
  nor (_04352_, _04351_, _04232_);
  and (_04353_, _04352_, _02592_);
  and (_04354_, _03874_, _03321_);
  nor (_04355_, _03864_, _03321_);
  and (_04356_, _03180_, _02785_);
  and (_04357_, _04352_, _02795_);
  and (_04358_, _03811_, _03321_);
  nand (_04359_, _03753_, \oc8051_golden_model_1.IRAM[0] [2]);
  nand (_04360_, _03588_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_04361_, _04360_, _03748_);
  nand (_04362_, _04361_, _04359_);
  not (_04363_, \oc8051_golden_model_1.IRAM[3] [2]);
  or (_04364_, _03753_, _04363_);
  not (_04365_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_04366_, _03588_, _04365_);
  and (_04367_, _04366_, _03755_);
  nand (_04368_, _04367_, _04364_);
  nand (_04369_, _04368_, _04362_);
  nand (_04370_, _04369_, _03337_);
  not (_04371_, \oc8051_golden_model_1.IRAM[7] [2]);
  or (_04372_, _03753_, _04371_);
  not (_04373_, \oc8051_golden_model_1.IRAM[6] [2]);
  or (_04374_, _03588_, _04373_);
  and (_04375_, _04374_, _03755_);
  nand (_04376_, _04375_, _04372_);
  not (_04377_, \oc8051_golden_model_1.IRAM[4] [2]);
  or (_04378_, _03588_, _04377_);
  not (_04379_, \oc8051_golden_model_1.IRAM[5] [2]);
  or (_04380_, _03753_, _04379_);
  and (_04381_, _04380_, _03748_);
  nand (_04382_, _04381_, _04378_);
  nand (_04383_, _04382_, _04376_);
  nand (_04384_, _04383_, _03761_);
  nand (_04385_, _04384_, _04370_);
  nand (_04386_, _04385_, _03148_);
  not (_04387_, \oc8051_golden_model_1.IRAM[11] [2]);
  or (_04388_, _03753_, _04387_);
  not (_04389_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_04390_, _03588_, _04389_);
  and (_04391_, _04390_, _03755_);
  nand (_04392_, _04391_, _04388_);
  nand (_04393_, _03753_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand (_04394_, _03588_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_04395_, _04394_, _03748_);
  nand (_04396_, _04395_, _04393_);
  nand (_04397_, _04396_, _04392_);
  nand (_04398_, _04397_, _03337_);
  not (_04399_, \oc8051_golden_model_1.IRAM[15] [2]);
  or (_04400_, _03753_, _04399_);
  not (_04401_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_04402_, _03588_, _04401_);
  and (_04403_, _04402_, _03755_);
  nand (_04404_, _04403_, _04400_);
  nand (_04405_, _03753_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand (_04406_, _03588_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_04407_, _04406_, _03748_);
  nand (_04408_, _04407_, _04405_);
  nand (_04409_, _04408_, _04404_);
  nand (_04410_, _04409_, _03761_);
  nand (_04411_, _04410_, _04398_);
  nand (_04412_, _04411_, _03778_);
  nand (_04413_, _04412_, _04386_);
  not (_04414_, _04413_);
  or (_04415_, _04414_, _03807_);
  nor (_04416_, _04122_, _02838_);
  and (_04417_, _03321_, _02838_);
  or (_04418_, _04417_, _02804_);
  or (_04419_, _04418_, _04416_);
  not (_04420_, _04352_);
  and (_04421_, _04420_, _02804_);
  not (_04422_, _04421_);
  nor (_04423_, _04121_, _04087_);
  and (_04424_, _04423_, _04422_);
  and (_04425_, _04424_, _04419_);
  and (_04426_, _04425_, _03992_);
  and (_04427_, _04426_, _04415_);
  nor (_04428_, _04427_, _04358_);
  and (_04429_, _03810_, _03179_);
  or (_04430_, _04429_, _04428_);
  nor (_04431_, _04352_, _02540_);
  nor (_04432_, _04431_, _03818_);
  not (_04433_, _04432_);
  nor (_04434_, _04433_, _04430_);
  and (_04435_, _03818_, _03321_);
  nor (_04436_, _04435_, _04434_);
  nor (_04437_, _04436_, _03376_);
  and (_04438_, _04413_, _03374_);
  nor (_04439_, _04438_, _03828_);
  and (_04440_, _04439_, _04437_);
  and (_04441_, _03828_, _03321_);
  nor (_04442_, _04441_, _04440_);
  and (_04443_, _03179_, _03827_);
  nor (_04444_, _04443_, _04442_);
  and (_04445_, _04444_, _03932_);
  nor (_04446_, _04445_, _04357_);
  and (_04447_, _02792_, _03179_);
  or (_04448_, _04447_, _04446_);
  nor (_04449_, _04352_, _02533_);
  nor (_04450_, _04449_, _02915_);
  not (_04451_, _04450_);
  nor (_04452_, _04451_, _04448_);
  and (_04453_, _04413_, _03842_);
  nor (_04454_, _04453_, _03841_);
  and (_04455_, _04454_, _04452_);
  nor (_04456_, _04455_, _04356_);
  nor (_04457_, _04456_, _02518_);
  and (_04458_, _04352_, _02518_);
  nor (_04459_, _04458_, _04457_);
  or (_04460_, _04459_, _04099_);
  nor (_04461_, _04460_, _04355_);
  and (_04462_, _04413_, _03870_);
  nor (_04463_, _04462_, _03874_);
  and (_04464_, _04463_, _04461_);
  nor (_04465_, _04464_, _04354_);
  nor (_04466_, _04465_, _02585_);
  and (_04467_, _04352_, _02585_);
  nor (_04468_, _04467_, _04466_);
  nor (_04469_, _03884_, _03321_);
  nor (_04470_, _04469_, _02594_);
  not (_04471_, _04470_);
  nor (_04472_, _04471_, _04468_);
  and (_04473_, _04352_, _02594_);
  nor (_04474_, _04473_, _04472_);
  and (_04475_, _03891_, _03320_);
  nor (_04476_, _04475_, _02592_);
  not (_04477_, _04476_);
  nor (_04478_, _04477_, _04474_);
  nor (_04479_, _04478_, _04353_);
  and (_04480_, _02904_, _02571_);
  nor (_04481_, _04480_, _04479_);
  and (_04482_, _04413_, _03898_);
  nor (_04483_, _04482_, _03900_);
  and (_04484_, _04483_, _04481_);
  and (_04485_, _03900_, _03321_);
  nor (_04486_, _04485_, _04484_);
  nor (_04487_, _04352_, _03907_);
  nor (_04488_, _04487_, _02780_);
  not (_04489_, _04488_);
  nor (_04490_, _04489_, _04486_);
  nor (_04491_, _04490_, _04350_);
  nor (_04492_, _04491_, _04349_);
  and (_04493_, _04413_, _03912_);
  nor (_04494_, _04493_, _03914_);
  and (_04495_, _04494_, _04492_);
  and (_04496_, _03914_, _03321_);
  nor (_04497_, _04496_, _04495_);
  nor (_04498_, _04497_, _04174_);
  not (_04499_, _04498_);
  nor (_04500_, _04499_, _04348_);
  and (_04501_, _04500_, _04176_);
  or (_04502_, _04501_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_04503_, _04234_, _02787_);
  nor (_04504_, _04352_, _03925_);
  nor (_04505_, _04504_, _04503_);
  and (_04506_, _04235_, _02787_);
  nor (_04507_, _04503_, _04237_);
  nor (_04508_, _04507_, _04506_);
  and (_04509_, _34976_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  not (_04510_, _04509_);
  and (_04511_, _04137_, _04138_);
  and (_04512_, _04511_, _04134_);
  nor (_04513_, _04512_, _04510_);
  and (_04514_, _04513_, _04508_);
  and (_04515_, _04514_, _04505_);
  and (_04516_, _04515_, _03924_);
  not (_04517_, _04516_);
  and (_04518_, _04517_, _04502_);
  nor (_04519_, _04510_, _04172_);
  not (_04520_, _04519_);
  nor (_04521_, _04520_, _03920_);
  not (_04522_, _04521_);
  nor (_04523_, _04522_, _04079_);
  not (_04524_, _04497_);
  nor (_04525_, _04520_, _04348_);
  and (_04526_, _04525_, _04524_);
  and (_04527_, _04526_, _04523_);
  not (_04528_, _04527_);
  not (_04529_, \oc8051_golden_model_1.IRAM[0] [7]);
  or (_04530_, _03588_, _04529_);
  not (_04531_, \oc8051_golden_model_1.IRAM[1] [7]);
  or (_04532_, _03753_, _04531_);
  and (_04533_, _04532_, _03748_);
  nand (_04534_, _04533_, _04530_);
  not (_04535_, \oc8051_golden_model_1.IRAM[3] [7]);
  or (_04536_, _03753_, _04535_);
  not (_04537_, \oc8051_golden_model_1.IRAM[2] [7]);
  or (_04538_, _03588_, _04537_);
  and (_04539_, _04538_, _03755_);
  nand (_04540_, _04539_, _04536_);
  nand (_04541_, _04540_, _04534_);
  nand (_04542_, _04541_, _03337_);
  not (_04543_, \oc8051_golden_model_1.IRAM[7] [7]);
  or (_04544_, _03753_, _04543_);
  not (_04545_, \oc8051_golden_model_1.IRAM[6] [7]);
  or (_04546_, _03588_, _04545_);
  and (_04547_, _04546_, _03755_);
  nand (_04548_, _04547_, _04544_);
  not (_04549_, \oc8051_golden_model_1.IRAM[4] [7]);
  or (_04550_, _03588_, _04549_);
  not (_04551_, \oc8051_golden_model_1.IRAM[5] [7]);
  or (_04552_, _03753_, _04551_);
  and (_04553_, _04552_, _03748_);
  nand (_04554_, _04553_, _04550_);
  nand (_04555_, _04554_, _04548_);
  nand (_04556_, _04555_, _03761_);
  nand (_04557_, _04556_, _04542_);
  nand (_04558_, _04557_, _03148_);
  not (_04559_, \oc8051_golden_model_1.IRAM[11] [7]);
  or (_04560_, _03753_, _04559_);
  not (_04561_, \oc8051_golden_model_1.IRAM[10] [7]);
  or (_04562_, _03588_, _04561_);
  and (_04563_, _04562_, _03755_);
  nand (_04564_, _04563_, _04560_);
  nand (_04565_, _03753_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand (_04566_, _03588_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_04567_, _04566_, _03748_);
  nand (_04568_, _04567_, _04565_);
  nand (_04569_, _04568_, _04564_);
  nand (_04570_, _04569_, _03337_);
  not (_04571_, \oc8051_golden_model_1.IRAM[15] [7]);
  or (_04572_, _03753_, _04571_);
  not (_04573_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_04574_, _03588_, _04573_);
  and (_04575_, _04574_, _03755_);
  nand (_04576_, _04575_, _04572_);
  nand (_04577_, _03753_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand (_04578_, _03588_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_04579_, _04578_, _03748_);
  nand (_04580_, _04579_, _04577_);
  nand (_04581_, _04580_, _04576_);
  nand (_04582_, _04581_, _03761_);
  nand (_04583_, _04582_, _04570_);
  nand (_04584_, _04583_, _03778_);
  nand (_04585_, _04584_, _04558_);
  or (_04586_, _04585_, _02858_);
  and (_04587_, _02889_, _02858_);
  and (_04588_, _04587_, _03179_);
  and (_04589_, _04588_, _03620_);
  and (_04590_, _03742_, _02836_);
  nor (_04591_, _03320_, _04318_);
  and (_04592_, _04591_, _04590_);
  and (_04593_, _04592_, _04589_);
  and (_04594_, _04593_, \oc8051_golden_model_1.TH1 [7]);
  and (_04595_, _04590_, _03320_);
  and (_04596_, _04595_, _02774_);
  not (_04597_, _03620_);
  and (_04598_, _04597_, _03179_);
  and (_04599_, _04598_, _04587_);
  and (_04600_, _04599_, _04596_);
  and (_04601_, _04600_, \oc8051_golden_model_1.SBUF [7]);
  nor (_04602_, _04601_, _04594_);
  and (_04603_, _03742_, _02835_);
  and (_04604_, _04603_, _04591_);
  and (_04605_, _04604_, _04589_);
  and (_04606_, _04605_, \oc8051_golden_model_1.TH0 [7]);
  and (_04607_, _04603_, _03320_);
  and (_04608_, _04607_, _02774_);
  and (_04609_, _04608_, _04599_);
  and (_04610_, _04609_, \oc8051_golden_model_1.SCON [7]);
  nor (_04611_, _04610_, _04606_);
  and (_04612_, _04611_, _04602_);
  and (_04613_, _04589_, _04318_);
  nor (_04614_, _03742_, _02835_);
  and (_04615_, _04614_, _03320_);
  and (_04616_, _04615_, _04613_);
  and (_04617_, _04616_, \oc8051_golden_model_1.DPH [7]);
  not (_04618_, _04617_);
  and (_04619_, _04596_, _04589_);
  and (_04620_, _04619_, \oc8051_golden_model_1.TMOD [7]);
  not (_04621_, _03179_);
  and (_04622_, _03620_, _04621_);
  and (_04623_, _04622_, _04587_);
  and (_04624_, _04623_, _04608_);
  and (_04625_, _04624_, \oc8051_golden_model_1.IE [7]);
  nor (_04626_, _04625_, _04620_);
  and (_04627_, _04626_, _04618_);
  nor (_04628_, _03742_, _02836_);
  not (_04629_, _04589_);
  nand (_04630_, _03320_, _02774_);
  nor (_04631_, _04630_, _04629_);
  and (_04632_, _04631_, _04628_);
  and (_04633_, _04632_, \oc8051_golden_model_1.TL0 [7]);
  and (_04634_, _04631_, _04614_);
  and (_04635_, _04634_, \oc8051_golden_model_1.TL1 [7]);
  nor (_04636_, _04635_, _04633_);
  and (_04637_, _04636_, _04627_);
  and (_04638_, _04637_, _04612_);
  and (_04639_, _04614_, _03321_);
  and (_04640_, _04639_, _04613_);
  and (_04641_, _04640_, \oc8051_golden_model_1.PCON [7]);
  not (_04642_, _04641_);
  and (_04643_, _04608_, _04589_);
  and (_04644_, _04643_, \oc8051_golden_model_1.TCON [7]);
  not (_04645_, _04644_);
  nor (_04646_, _03620_, _03179_);
  and (_04647_, _04646_, _04587_);
  and (_04648_, _04647_, _04608_);
  and (_04649_, _04648_, \oc8051_golden_model_1.IP [7]);
  and (_04650_, _03320_, _04318_);
  and (_04651_, _04650_, _04603_);
  nor (_04652_, _02889_, _02743_);
  and (_04653_, _04652_, _04622_);
  and (_04654_, _04653_, _04651_);
  and (_04655_, _04654_, \oc8051_golden_model_1.ACC [7]);
  nor (_04656_, _04655_, _04649_);
  and (_04657_, _04652_, _04598_);
  and (_04658_, _04657_, _04651_);
  and (_04659_, _04658_, \oc8051_golden_model_1.PSW [7]);
  and (_04660_, _04652_, _04646_);
  and (_04661_, _04660_, _04651_);
  and (_04662_, _04661_, \oc8051_golden_model_1.B [7]);
  nor (_04663_, _04662_, _04659_);
  and (_04664_, _04663_, _04656_);
  and (_04665_, _04664_, _04645_);
  and (_04666_, _04665_, _04642_);
  and (_04667_, _04613_, _04595_);
  and (_04668_, _04667_, \oc8051_golden_model_1.SP [7]);
  and (_04669_, _04628_, _03320_);
  and (_04670_, _04669_, _04613_);
  and (_04671_, _04670_, \oc8051_golden_model_1.DPL [7]);
  nor (_04672_, _04671_, _04668_);
  and (_04673_, _04651_, _04589_);
  and (_04674_, _04673_, \oc8051_golden_model_1.P0 [7]);
  not (_04675_, _04674_);
  and (_04676_, _04651_, _04599_);
  and (_04677_, _04676_, \oc8051_golden_model_1.P1 [7]);
  not (_04678_, _04677_);
  and (_04679_, _04651_, _04623_);
  and (_04680_, _04679_, \oc8051_golden_model_1.P2 [7]);
  and (_04681_, _04651_, _04647_);
  and (_04682_, _04681_, \oc8051_golden_model_1.P3 [7]);
  nor (_04683_, _04682_, _04680_);
  and (_04684_, _04683_, _04678_);
  and (_04685_, _04684_, _04675_);
  and (_04686_, _04685_, _04672_);
  and (_04687_, _04686_, _04666_);
  and (_04688_, _04687_, _04638_);
  and (_04689_, _04688_, _04586_);
  not (_04690_, _04689_);
  nand (_04691_, _03753_, \oc8051_golden_model_1.IRAM[0] [6]);
  nand (_04692_, _03588_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_04693_, _04692_, _03748_);
  nand (_04694_, _04693_, _04691_);
  nand (_04695_, _03588_, \oc8051_golden_model_1.IRAM[3] [6]);
  nand (_04696_, _03753_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_04697_, _04696_, _03755_);
  nand (_04698_, _04697_, _04695_);
  nand (_04699_, _04698_, _04694_);
  nand (_04700_, _04699_, _03337_);
  nand (_04701_, _03588_, \oc8051_golden_model_1.IRAM[7] [6]);
  nand (_04702_, _03753_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_04703_, _04702_, _03755_);
  nand (_04704_, _04703_, _04701_);
  nand (_04705_, _03753_, \oc8051_golden_model_1.IRAM[4] [6]);
  nand (_04706_, _03588_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_04707_, _04706_, _03748_);
  nand (_04708_, _04707_, _04705_);
  nand (_04709_, _04708_, _04704_);
  nand (_04710_, _04709_, _03761_);
  nand (_04711_, _04710_, _04700_);
  nand (_04712_, _04711_, _03148_);
  nand (_04713_, _03588_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_04714_, _03753_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_04715_, _04714_, _03755_);
  nand (_04716_, _04715_, _04713_);
  nand (_04717_, _03753_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand (_04718_, _03588_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_04719_, _04718_, _03748_);
  nand (_04720_, _04719_, _04717_);
  nand (_04721_, _04720_, _04716_);
  nand (_04722_, _04721_, _03337_);
  nand (_04723_, _03588_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_04724_, _03753_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_04725_, _04724_, _03755_);
  nand (_04726_, _04725_, _04723_);
  nand (_04727_, _03753_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand (_04728_, _03588_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_04729_, _04728_, _03748_);
  nand (_04730_, _04729_, _04727_);
  nand (_04731_, _04730_, _04726_);
  nand (_04732_, _04731_, _03761_);
  nand (_04733_, _04732_, _04722_);
  nand (_04734_, _04733_, _03778_);
  nand (_04735_, _04734_, _04712_);
  or (_04736_, _04735_, _02858_);
  and (_04737_, _04593_, \oc8051_golden_model_1.TH1 [6]);
  and (_04738_, _04600_, \oc8051_golden_model_1.SBUF [6]);
  nor (_04739_, _04738_, _04737_);
  and (_04740_, _04605_, \oc8051_golden_model_1.TH0 [6]);
  and (_04741_, _04609_, \oc8051_golden_model_1.SCON [6]);
  nor (_04742_, _04741_, _04740_);
  and (_04743_, _04742_, _04739_);
  and (_04744_, _04616_, \oc8051_golden_model_1.DPH [6]);
  not (_04745_, _04744_);
  and (_04746_, _04619_, \oc8051_golden_model_1.TMOD [6]);
  and (_04747_, _04624_, \oc8051_golden_model_1.IE [6]);
  nor (_04748_, _04747_, _04746_);
  and (_04749_, _04748_, _04745_);
  and (_04750_, _04632_, \oc8051_golden_model_1.TL0 [6]);
  and (_04751_, _04634_, \oc8051_golden_model_1.TL1 [6]);
  nor (_04752_, _04751_, _04750_);
  and (_04753_, _04752_, _04749_);
  and (_04754_, _04753_, _04743_);
  and (_04755_, _04640_, \oc8051_golden_model_1.PCON [6]);
  not (_04756_, _04755_);
  and (_04757_, _04643_, \oc8051_golden_model_1.TCON [6]);
  not (_04758_, _04757_);
  and (_04759_, _04648_, \oc8051_golden_model_1.IP [6]);
  and (_04760_, _04654_, \oc8051_golden_model_1.ACC [6]);
  nor (_04761_, _04760_, _04759_);
  and (_04762_, _04658_, \oc8051_golden_model_1.PSW [6]);
  and (_04763_, _04661_, \oc8051_golden_model_1.B [6]);
  nor (_04764_, _04763_, _04762_);
  and (_04765_, _04764_, _04761_);
  and (_04766_, _04765_, _04758_);
  and (_04767_, _04766_, _04756_);
  and (_04768_, _04667_, \oc8051_golden_model_1.SP [6]);
  and (_04769_, _04670_, \oc8051_golden_model_1.DPL [6]);
  nor (_04770_, _04769_, _04768_);
  and (_04771_, _04673_, \oc8051_golden_model_1.P0 [6]);
  not (_04772_, _04771_);
  and (_04773_, _04676_, \oc8051_golden_model_1.P1 [6]);
  not (_04774_, _04773_);
  and (_04775_, _04679_, \oc8051_golden_model_1.P2 [6]);
  and (_04776_, _04681_, \oc8051_golden_model_1.P3 [6]);
  nor (_04777_, _04776_, _04775_);
  and (_04778_, _04777_, _04774_);
  and (_04779_, _04778_, _04772_);
  and (_04780_, _04779_, _04770_);
  and (_04781_, _04780_, _04767_);
  and (_04782_, _04781_, _04754_);
  and (_04783_, _04782_, _04736_);
  not (_04784_, _04783_);
  nand (_04785_, _03753_, \oc8051_golden_model_1.IRAM[0] [5]);
  not (_04786_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_04787_, _03753_, _04786_);
  and (_04788_, _04787_, _03748_);
  nand (_04789_, _04788_, _04785_);
  nand (_04790_, _03588_, \oc8051_golden_model_1.IRAM[3] [5]);
  not (_04791_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_04792_, _03588_, _04791_);
  and (_04793_, _04792_, _03755_);
  nand (_04794_, _04793_, _04790_);
  nand (_04795_, _04794_, _04789_);
  nand (_04796_, _04795_, _03337_);
  not (_04797_, \oc8051_golden_model_1.IRAM[7] [5]);
  or (_04798_, _03753_, _04797_);
  not (_04799_, \oc8051_golden_model_1.IRAM[6] [5]);
  or (_04800_, _03588_, _04799_);
  and (_04801_, _04800_, _03755_);
  nand (_04802_, _04801_, _04798_);
  not (_04803_, \oc8051_golden_model_1.IRAM[4] [5]);
  or (_04804_, _03588_, _04803_);
  not (_04805_, \oc8051_golden_model_1.IRAM[5] [5]);
  or (_04806_, _03753_, _04805_);
  and (_04807_, _04806_, _03748_);
  nand (_04808_, _04807_, _04804_);
  nand (_04809_, _04808_, _04802_);
  nand (_04810_, _04809_, _03761_);
  nand (_04811_, _04810_, _04796_);
  nand (_04812_, _04811_, _03148_);
  nand (_04813_, _03588_, \oc8051_golden_model_1.IRAM[11] [5]);
  not (_04814_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_04815_, _03588_, _04814_);
  and (_04816_, _04815_, _03755_);
  nand (_04817_, _04816_, _04813_);
  nand (_04818_, _03753_, \oc8051_golden_model_1.IRAM[8] [5]);
  not (_04819_, \oc8051_golden_model_1.IRAM[9] [5]);
  or (_04820_, _03753_, _04819_);
  and (_04821_, _04820_, _03748_);
  nand (_04822_, _04821_, _04818_);
  nand (_04823_, _04822_, _04817_);
  nand (_04824_, _04823_, _03337_);
  nand (_04825_, _03588_, \oc8051_golden_model_1.IRAM[15] [5]);
  not (_04826_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_04827_, _03588_, _04826_);
  and (_04828_, _04827_, _03755_);
  nand (_04829_, _04828_, _04825_);
  nand (_04830_, _03753_, \oc8051_golden_model_1.IRAM[12] [5]);
  not (_04831_, \oc8051_golden_model_1.IRAM[13] [5]);
  or (_04832_, _03753_, _04831_);
  and (_04833_, _04832_, _03748_);
  nand (_04834_, _04833_, _04830_);
  nand (_04835_, _04834_, _04829_);
  nand (_04836_, _04835_, _03761_);
  nand (_04837_, _04836_, _04824_);
  nand (_04838_, _04837_, _03778_);
  nand (_04839_, _04838_, _04812_);
  or (_04840_, _04839_, _02858_);
  and (_04841_, _04605_, \oc8051_golden_model_1.TH0 [5]);
  and (_04842_, _04609_, \oc8051_golden_model_1.SCON [5]);
  nor (_04843_, _04842_, _04841_);
  and (_04844_, _04619_, \oc8051_golden_model_1.TMOD [5]);
  and (_04845_, _04593_, \oc8051_golden_model_1.TH1 [5]);
  nor (_04846_, _04845_, _04844_);
  and (_04847_, _04846_, _04843_);
  and (_04848_, _04634_, \oc8051_golden_model_1.TL1 [5]);
  not (_04849_, _04848_);
  and (_04850_, _04632_, \oc8051_golden_model_1.TL0 [5]);
  and (_04851_, _04616_, \oc8051_golden_model_1.DPH [5]);
  nor (_04852_, _04851_, _04850_);
  and (_04853_, _04852_, _04849_);
  and (_04854_, _04853_, _04847_);
  and (_04855_, _04640_, \oc8051_golden_model_1.PCON [5]);
  not (_04856_, _04855_);
  and (_04857_, _04648_, \oc8051_golden_model_1.IP [5]);
  not (_04858_, _04857_);
  and (_04859_, _04658_, \oc8051_golden_model_1.PSW [5]);
  and (_04860_, _04654_, \oc8051_golden_model_1.ACC [5]);
  nor (_04861_, _04860_, _04859_);
  and (_04862_, _04861_, _04858_);
  and (_04863_, _04600_, \oc8051_golden_model_1.SBUF [5]);
  not (_04864_, _04863_);
  and (_04865_, _04624_, \oc8051_golden_model_1.IE [5]);
  and (_04866_, _04661_, \oc8051_golden_model_1.B [5]);
  nor (_04867_, _04866_, _04865_);
  and (_04868_, _04867_, _04864_);
  and (_04869_, _04868_, _04862_);
  and (_04870_, _04869_, _04856_);
  and (_04871_, _04667_, \oc8051_golden_model_1.SP [5]);
  not (_04872_, _04871_);
  and (_04873_, _04670_, \oc8051_golden_model_1.DPL [5]);
  and (_04874_, _04643_, \oc8051_golden_model_1.TCON [5]);
  nor (_04875_, _04874_, _04873_);
  and (_04876_, _04875_, _04872_);
  and (_04877_, _04673_, \oc8051_golden_model_1.P0 [5]);
  not (_04878_, _04877_);
  and (_04879_, _04676_, \oc8051_golden_model_1.P1 [5]);
  not (_04880_, _04879_);
  and (_04881_, _04679_, \oc8051_golden_model_1.P2 [5]);
  and (_04882_, _04681_, \oc8051_golden_model_1.P3 [5]);
  nor (_04883_, _04882_, _04881_);
  and (_04884_, _04883_, _04880_);
  and (_04885_, _04884_, _04878_);
  and (_04886_, _04885_, _04876_);
  and (_04887_, _04886_, _04870_);
  and (_04888_, _04887_, _04854_);
  and (_04889_, _04888_, _04840_);
  not (_04890_, _04889_);
  or (_04891_, _04226_, _02858_);
  and (_04892_, _04640_, \oc8051_golden_model_1.PCON [3]);
  not (_04893_, _04892_);
  and (_04894_, _04600_, \oc8051_golden_model_1.SBUF [3]);
  and (_04895_, _04624_, \oc8051_golden_model_1.IE [3]);
  nor (_04896_, _04895_, _04894_);
  and (_04897_, _04896_, _04893_);
  and (_04898_, _04679_, \oc8051_golden_model_1.P2 [3]);
  and (_04899_, _04681_, \oc8051_golden_model_1.P3 [3]);
  nor (_04900_, _04899_, _04898_);
  and (_04901_, _04900_, _04897_);
  and (_04902_, _04658_, \oc8051_golden_model_1.PSW [3]);
  and (_04903_, _04654_, \oc8051_golden_model_1.ACC [3]);
  nor (_04904_, _04903_, _04902_);
  and (_04905_, _04648_, \oc8051_golden_model_1.IP [3]);
  and (_04906_, _04661_, \oc8051_golden_model_1.B [3]);
  nor (_04907_, _04906_, _04905_);
  and (_04908_, _04907_, _04904_);
  and (_04909_, _04643_, \oc8051_golden_model_1.TCON [3]);
  and (_04910_, _04605_, \oc8051_golden_model_1.TH0 [3]);
  nor (_04911_, _04910_, _04909_);
  and (_04912_, _04676_, \oc8051_golden_model_1.P1 [3]);
  not (_04913_, _04614_);
  nor (_04914_, _04913_, _04630_);
  and (_04915_, _04914_, _04589_);
  and (_04916_, _04915_, \oc8051_golden_model_1.TL1 [3]);
  nor (_04917_, _04916_, _04912_);
  and (_04918_, _04917_, _04911_);
  and (_04919_, _04609_, \oc8051_golden_model_1.SCON [3]);
  and (_04920_, _04593_, \oc8051_golden_model_1.TH1 [3]);
  nor (_04921_, _04920_, _04919_);
  and (_04922_, _04619_, \oc8051_golden_model_1.TMOD [3]);
  and (_04923_, _04632_, \oc8051_golden_model_1.TL0 [3]);
  nor (_04924_, _04923_, _04922_);
  and (_04925_, _04924_, _04921_);
  and (_04926_, _04925_, _04918_);
  and (_04927_, _04926_, _04908_);
  and (_04928_, _04927_, _04901_);
  and (_04929_, _04673_, \oc8051_golden_model_1.P0 [3]);
  not (_04930_, _04929_);
  and (_04931_, _04667_, \oc8051_golden_model_1.SP [3]);
  and (_04932_, _04670_, \oc8051_golden_model_1.DPL [3]);
  nor (_04933_, _04932_, _04931_);
  nand (_04934_, _04616_, \oc8051_golden_model_1.DPH [3]);
  and (_04935_, _04934_, _04933_);
  and (_04936_, _04935_, _04930_);
  and (_04937_, _04936_, _04928_);
  and (_04938_, _04937_, _04891_);
  not (_04939_, _04938_);
  or (_04940_, _03989_, _02858_);
  and (_04941_, _04605_, \oc8051_golden_model_1.TH0 [1]);
  and (_04942_, _04600_, \oc8051_golden_model_1.SBUF [1]);
  nor (_04943_, _04942_, _04941_);
  and (_04944_, _04619_, \oc8051_golden_model_1.TMOD [1]);
  and (_04945_, _04609_, \oc8051_golden_model_1.SCON [1]);
  nor (_04946_, _04945_, _04944_);
  and (_04947_, _04946_, _04943_);
  and (_04948_, _04632_, \oc8051_golden_model_1.TL0 [1]);
  and (_04949_, _04593_, \oc8051_golden_model_1.TH1 [1]);
  and (_04950_, _04624_, \oc8051_golden_model_1.IE [1]);
  nor (_04951_, _04950_, _04949_);
  not (_04952_, _04951_);
  nor (_04953_, _04952_, _04948_);
  and (_04954_, _04616_, \oc8051_golden_model_1.DPH [1]);
  and (_04955_, _04634_, \oc8051_golden_model_1.TL1 [1]);
  nor (_04956_, _04955_, _04954_);
  and (_04957_, _04956_, _04953_);
  and (_04958_, _04957_, _04947_);
  and (_04959_, _04640_, \oc8051_golden_model_1.PCON [1]);
  not (_04960_, _04959_);
  and (_04961_, _04643_, \oc8051_golden_model_1.TCON [1]);
  not (_04962_, _04961_);
  and (_04963_, _04658_, \oc8051_golden_model_1.PSW [1]);
  and (_04964_, _04654_, \oc8051_golden_model_1.ACC [1]);
  nor (_04965_, _04964_, _04963_);
  and (_04966_, _04648_, \oc8051_golden_model_1.IP [1]);
  and (_04967_, _04661_, \oc8051_golden_model_1.B [1]);
  nor (_04968_, _04967_, _04966_);
  and (_04969_, _04968_, _04965_);
  and (_04970_, _04969_, _04962_);
  and (_04971_, _04970_, _04960_);
  and (_04972_, _04667_, \oc8051_golden_model_1.SP [1]);
  and (_04973_, _04670_, \oc8051_golden_model_1.DPL [1]);
  nor (_04974_, _04973_, _04972_);
  and (_04975_, _04673_, \oc8051_golden_model_1.P0 [1]);
  not (_04976_, _04975_);
  and (_04977_, _04676_, \oc8051_golden_model_1.P1 [1]);
  not (_04978_, _04977_);
  and (_04979_, _04679_, \oc8051_golden_model_1.P2 [1]);
  and (_04980_, _04681_, \oc8051_golden_model_1.P3 [1]);
  nor (_04981_, _04980_, _04979_);
  and (_04982_, _04981_, _04978_);
  and (_04983_, _04982_, _04976_);
  and (_04984_, _04983_, _04974_);
  and (_04985_, _04984_, _04971_);
  and (_04986_, _04985_, _04958_);
  and (_04987_, _04986_, _04940_);
  not (_04988_, _04987_);
  or (_04989_, _03823_, _02858_);
  and (_04990_, _04673_, \oc8051_golden_model_1.P0 [0]);
  not (_04991_, _04990_);
  and (_04992_, _04648_, \oc8051_golden_model_1.IP [0]);
  and (_04993_, _04654_, \oc8051_golden_model_1.ACC [0]);
  nor (_04994_, _04993_, _04992_);
  and (_04995_, _04658_, \oc8051_golden_model_1.PSW [0]);
  and (_04996_, _04661_, \oc8051_golden_model_1.B [0]);
  nor (_04997_, _04996_, _04995_);
  and (_04998_, _04997_, _04994_);
  and (_04999_, _04676_, \oc8051_golden_model_1.P1 [0]);
  not (_05000_, _04999_);
  and (_05001_, _04679_, \oc8051_golden_model_1.P2 [0]);
  and (_05002_, _04681_, \oc8051_golden_model_1.P3 [0]);
  nor (_05003_, _05002_, _05001_);
  and (_05004_, _05003_, _05000_);
  and (_05005_, _05004_, _04998_);
  and (_05006_, _05005_, _04991_);
  and (_05007_, _04667_, \oc8051_golden_model_1.SP [0]);
  and (_05008_, _04670_, \oc8051_golden_model_1.DPL [0]);
  nor (_05009_, _05008_, _05007_);
  and (_05010_, _04640_, \oc8051_golden_model_1.PCON [0]);
  not (_05011_, _05010_);
  and (_05012_, _04600_, \oc8051_golden_model_1.SBUF [0]);
  and (_05013_, _04624_, \oc8051_golden_model_1.IE [0]);
  nor (_05014_, _05013_, _05012_);
  and (_05015_, _05014_, _05011_);
  and (_05016_, _05015_, _05009_);
  and (_05017_, _05016_, _05006_);
  and (_05018_, _04632_, \oc8051_golden_model_1.TL0 [0]);
  not (_05019_, _05018_);
  and (_05020_, _04619_, \oc8051_golden_model_1.TMOD [0]);
  and (_05021_, _04609_, \oc8051_golden_model_1.SCON [0]);
  nor (_05022_, _05021_, _05020_);
  and (_05023_, _04643_, \oc8051_golden_model_1.TCON [0]);
  and (_05024_, _04593_, \oc8051_golden_model_1.TH1 [0]);
  nor (_05025_, _05024_, _05023_);
  and (_05026_, _05025_, _05022_);
  and (_05027_, _05026_, _05019_);
  and (_05028_, _04634_, \oc8051_golden_model_1.TL1 [0]);
  not (_05029_, _05028_);
  and (_05030_, _04605_, \oc8051_golden_model_1.TH0 [0]);
  and (_05031_, _04616_, \oc8051_golden_model_1.DPH [0]);
  nor (_05032_, _05031_, _05030_);
  and (_05033_, _05032_, _05029_);
  and (_05034_, _05033_, _05027_);
  and (_05035_, _05034_, _05017_);
  nand (_05036_, _05035_, _04989_);
  and (_05037_, _05036_, _04988_);
  or (_05038_, _04413_, _02858_);
  and (_05039_, _04605_, \oc8051_golden_model_1.TH0 [2]);
  and (_05040_, _04600_, \oc8051_golden_model_1.SBUF [2]);
  nor (_05041_, _05040_, _05039_);
  and (_05042_, _04619_, \oc8051_golden_model_1.TMOD [2]);
  and (_05043_, _04609_, \oc8051_golden_model_1.SCON [2]);
  nor (_05044_, _05043_, _05042_);
  and (_05045_, _05044_, _05041_);
  and (_05046_, _04632_, \oc8051_golden_model_1.TL0 [2]);
  and (_05047_, _04593_, \oc8051_golden_model_1.TH1 [2]);
  and (_05048_, _04624_, \oc8051_golden_model_1.IE [2]);
  nor (_05049_, _05048_, _05047_);
  not (_05050_, _05049_);
  nor (_05051_, _05050_, _05046_);
  and (_05052_, _04616_, \oc8051_golden_model_1.DPH [2]);
  and (_05053_, _04634_, \oc8051_golden_model_1.TL1 [2]);
  nor (_05054_, _05053_, _05052_);
  and (_05055_, _05054_, _05051_);
  and (_05056_, _05055_, _05045_);
  and (_05057_, _04640_, \oc8051_golden_model_1.PCON [2]);
  not (_05058_, _05057_);
  and (_05059_, _04643_, \oc8051_golden_model_1.TCON [2]);
  not (_05060_, _05059_);
  and (_05061_, _04648_, \oc8051_golden_model_1.IP [2]);
  and (_05062_, _04661_, \oc8051_golden_model_1.B [2]);
  nor (_05063_, _05062_, _05061_);
  and (_05064_, _04658_, \oc8051_golden_model_1.PSW [2]);
  and (_05065_, _04654_, \oc8051_golden_model_1.ACC [2]);
  nor (_05066_, _05065_, _05064_);
  and (_05067_, _05066_, _05063_);
  and (_05068_, _05067_, _05060_);
  and (_05069_, _05068_, _05058_);
  and (_05070_, _04667_, \oc8051_golden_model_1.SP [2]);
  and (_05071_, _04670_, \oc8051_golden_model_1.DPL [2]);
  nor (_05072_, _05071_, _05070_);
  and (_05073_, _04673_, \oc8051_golden_model_1.P0 [2]);
  not (_05074_, _05073_);
  and (_05075_, _04676_, \oc8051_golden_model_1.P1 [2]);
  not (_05076_, _05075_);
  and (_05077_, _04679_, \oc8051_golden_model_1.P2 [2]);
  and (_05078_, _04681_, \oc8051_golden_model_1.P3 [2]);
  nor (_05079_, _05078_, _05077_);
  and (_05080_, _05079_, _05076_);
  and (_05081_, _05080_, _05074_);
  and (_05082_, _05081_, _05072_);
  and (_05083_, _05082_, _05069_);
  and (_05084_, _05083_, _05056_);
  and (_05085_, _05084_, _05038_);
  not (_05086_, _05085_);
  and (_05087_, _05086_, _05037_);
  and (_05088_, _05087_, _04939_);
  nand (_05089_, _03753_, \oc8051_golden_model_1.IRAM[0] [4]);
  not (_05090_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_05091_, _03753_, _05090_);
  and (_05092_, _05091_, _03748_);
  nand (_05093_, _05092_, _05089_);
  nand (_05094_, _03588_, \oc8051_golden_model_1.IRAM[3] [4]);
  not (_05095_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_05096_, _03588_, _05095_);
  and (_05097_, _05096_, _03755_);
  nand (_05098_, _05097_, _05094_);
  nand (_05099_, _05098_, _05093_);
  nand (_05100_, _05099_, _03337_);
  not (_05101_, \oc8051_golden_model_1.IRAM[7] [4]);
  or (_05102_, _03753_, _05101_);
  not (_05103_, \oc8051_golden_model_1.IRAM[6] [4]);
  or (_05104_, _03588_, _05103_);
  and (_05105_, _05104_, _03755_);
  nand (_05106_, _05105_, _05102_);
  not (_05107_, \oc8051_golden_model_1.IRAM[4] [4]);
  or (_05108_, _03588_, _05107_);
  not (_05109_, \oc8051_golden_model_1.IRAM[5] [4]);
  or (_05110_, _03753_, _05109_);
  and (_05111_, _05110_, _03748_);
  nand (_05112_, _05111_, _05108_);
  nand (_05113_, _05112_, _05106_);
  nand (_05114_, _05113_, _03761_);
  nand (_05115_, _05114_, _05100_);
  nand (_05116_, _05115_, _03148_);
  nand (_05117_, _03588_, \oc8051_golden_model_1.IRAM[11] [4]);
  not (_05118_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_05119_, _03588_, _05118_);
  and (_05120_, _05119_, _03755_);
  nand (_05121_, _05120_, _05117_);
  nand (_05122_, _03753_, \oc8051_golden_model_1.IRAM[8] [4]);
  not (_05123_, \oc8051_golden_model_1.IRAM[9] [4]);
  or (_05124_, _03753_, _05123_);
  and (_05125_, _05124_, _03748_);
  nand (_05126_, _05125_, _05122_);
  nand (_05127_, _05126_, _05121_);
  nand (_05128_, _05127_, _03337_);
  nand (_05129_, _03588_, \oc8051_golden_model_1.IRAM[15] [4]);
  not (_05130_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_05131_, _03588_, _05130_);
  and (_05132_, _05131_, _03755_);
  nand (_05133_, _05132_, _05129_);
  nand (_05134_, _03753_, \oc8051_golden_model_1.IRAM[12] [4]);
  not (_05135_, \oc8051_golden_model_1.IRAM[13] [4]);
  or (_05136_, _03753_, _05135_);
  and (_05137_, _05136_, _03748_);
  nand (_05138_, _05137_, _05134_);
  nand (_05139_, _05138_, _05133_);
  nand (_05140_, _05139_, _03761_);
  nand (_05141_, _05140_, _05128_);
  nand (_05142_, _05141_, _03778_);
  nand (_05143_, _05142_, _05116_);
  or (_05144_, _05143_, _02858_);
  and (_05145_, _04667_, \oc8051_golden_model_1.SP [4]);
  and (_05146_, _04670_, \oc8051_golden_model_1.DPL [4]);
  nor (_05147_, _05146_, _05145_);
  and (_05148_, _04643_, \oc8051_golden_model_1.TCON [4]);
  and (_05149_, _04605_, \oc8051_golden_model_1.TH0 [4]);
  nor (_05150_, _05149_, _05148_);
  and (_05151_, _04676_, \oc8051_golden_model_1.P1 [4]);
  and (_05152_, _04915_, \oc8051_golden_model_1.TL1 [4]);
  nor (_05153_, _05152_, _05151_);
  and (_05154_, _05153_, _05150_);
  and (_05155_, _04609_, \oc8051_golden_model_1.SCON [4]);
  and (_05156_, _04593_, \oc8051_golden_model_1.TH1 [4]);
  nor (_05157_, _05156_, _05155_);
  and (_05158_, _04632_, \oc8051_golden_model_1.TL0 [4]);
  and (_05159_, _04619_, \oc8051_golden_model_1.TMOD [4]);
  nor (_05160_, _05159_, _05158_);
  and (_05161_, _05160_, _05157_);
  and (_05162_, _05161_, _05154_);
  and (_05163_, _05162_, _05147_);
  and (_05164_, _04679_, \oc8051_golden_model_1.P2 [4]);
  and (_05165_, _04681_, \oc8051_golden_model_1.P3 [4]);
  nor (_05166_, _05165_, _05164_);
  and (_05167_, _04640_, \oc8051_golden_model_1.PCON [4]);
  not (_05168_, _05167_);
  and (_05169_, _04600_, \oc8051_golden_model_1.SBUF [4]);
  and (_05170_, _04624_, \oc8051_golden_model_1.IE [4]);
  nor (_05171_, _05170_, _05169_);
  and (_05172_, _05171_, _05168_);
  and (_05173_, _05172_, _05166_);
  and (_05174_, _04658_, \oc8051_golden_model_1.PSW [4]);
  and (_05175_, _04654_, \oc8051_golden_model_1.ACC [4]);
  nor (_05176_, _05175_, _05174_);
  and (_05177_, _04648_, \oc8051_golden_model_1.IP [4]);
  and (_05178_, _04661_, \oc8051_golden_model_1.B [4]);
  nor (_05179_, _05178_, _05177_);
  and (_05180_, _05179_, _05176_);
  and (_05181_, _04673_, \oc8051_golden_model_1.P0 [4]);
  and (_05182_, _04650_, _04614_);
  and (_05183_, _05182_, _04589_);
  and (_05184_, _05183_, \oc8051_golden_model_1.DPH [4]);
  nor (_05185_, _05184_, _05181_);
  and (_05186_, _05185_, _05180_);
  and (_05187_, _05186_, _05173_);
  and (_05188_, _05187_, _05163_);
  and (_05189_, _05188_, _05144_);
  not (_05190_, _05189_);
  and (_05191_, _05190_, _05088_);
  and (_05192_, _05191_, _04890_);
  and (_05193_, _05192_, _04784_);
  nor (_05194_, _05193_, _04690_);
  and (_05195_, _05193_, _04690_);
  nor (_05196_, _05195_, _05194_);
  and (_05197_, _05196_, _03914_);
  not (_05198_, _04585_);
  not (_05199_, _04839_);
  not (_05200_, _05143_);
  nor (_05201_, _03989_, _03823_);
  nor (_05202_, _04413_, _04226_);
  and (_05203_, _05202_, _05201_);
  and (_05204_, _05203_, _05200_);
  and (_05205_, _05204_, _05199_);
  nor (_05206_, _05205_, _05198_);
  and (_05207_, _04735_, _04585_);
  nor (_05208_, _04735_, _04585_);
  nor (_05209_, _05208_, _05207_);
  not (_05210_, _05209_);
  and (_05211_, _05210_, _05205_);
  nor (_05212_, _05211_, _05206_);
  not (_05213_, _04125_);
  not (_05214_, _03698_);
  and (_05215_, _04113_, _05214_);
  and (_05216_, _05215_, _05213_);
  nor (_05217_, _05216_, _05212_);
  not (_05218_, _02572_);
  not (_05219_, _02988_);
  not (_05220_, _03880_);
  and (_05221_, _02991_, _02743_);
  not (_05222_, _05221_);
  and (_05223_, _03107_, _02743_);
  not (_05224_, _05223_);
  and (_05225_, _02977_, _02743_);
  and (_05226_, _03069_, _01146_);
  and (_05227_, _03075_, _01110_);
  nor (_05228_, _05227_, _05226_);
  and (_05229_, _03034_, _01086_);
  and (_05230_, _03082_, _01134_);
  nor (_05231_, _05230_, _05229_);
  and (_05232_, _05231_, _05228_);
  and (_05233_, _03080_, _01097_);
  and (_05234_, _03046_, _01114_);
  nor (_05235_, _05234_, _05233_);
  and (_05236_, _03077_, _01139_);
  and (_05237_, _03055_, _01142_);
  nor (_05238_, _05237_, _05236_);
  and (_05239_, _05238_, _05235_);
  and (_05240_, _05239_, _05232_);
  and (_05241_, _03037_, _01082_);
  and (_05242_, _03071_, _01058_);
  nor (_05243_, _05242_, _05241_);
  and (_05244_, _03066_, _01126_);
  and (_05245_, _03050_, _01102_);
  nor (_05246_, _05245_, _05244_);
  and (_05247_, _05246_, _05243_);
  and (_05248_, _03063_, _01131_);
  and (_05249_, _03043_, _01092_);
  nor (_05250_, _05249_, _05248_);
  and (_05251_, _03052_, _01106_);
  and (_05252_, _03057_, _01117_);
  nor (_05253_, _05252_, _05251_);
  and (_05254_, _05253_, _05250_);
  and (_05255_, _05254_, _05247_);
  and (_05256_, _05255_, _05240_);
  and (_05257_, _05256_, _04689_);
  nor (_05258_, _05256_, _04689_);
  nor (_05259_, _05258_, _05257_);
  and (_05260_, _05259_, _05225_);
  not (_05261_, _02974_);
  not (_05262_, _03870_);
  nor (_05263_, _04091_, _04085_);
  and (_05264_, _03857_, _02584_);
  nor (_05265_, _05264_, _04094_);
  and (_05266_, _05265_, _05263_);
  and (_05267_, _05266_, _05262_);
  and (_05268_, _05267_, _05261_);
  or (_05269_, _05268_, _02858_);
  not (_05270_, _03827_);
  not (_05271_, _02892_);
  nor (_05272_, _03621_, _02775_);
  and (_05273_, _05272_, _03181_);
  and (_05274_, _05273_, _05271_);
  and (_05275_, _05274_, _04589_);
  and (_05276_, _05275_, \oc8051_golden_model_1.TCON [7]);
  and (_05277_, _05273_, _02892_);
  and (_05278_, _04623_, _05277_);
  and (_05279_, _05278_, \oc8051_golden_model_1.P2 [7]);
  and (_05280_, _04647_, _05277_);
  and (_05281_, _05280_, \oc8051_golden_model_1.P3 [7]);
  or (_05282_, _05281_, _05279_);
  nor (_05283_, _05282_, _05276_);
  and (_05284_, _05274_, _04647_);
  and (_05285_, _05284_, \oc8051_golden_model_1.IP [7]);
  and (_05286_, _04660_, _05277_);
  and (_05287_, _05286_, \oc8051_golden_model_1.B [7]);
  nor (_05288_, _05287_, _05285_);
  and (_05289_, _04657_, _05277_);
  and (_05290_, _05289_, \oc8051_golden_model_1.PSW [7]);
  and (_05291_, _04653_, _05277_);
  and (_05292_, _05291_, \oc8051_golden_model_1.ACC [7]);
  nor (_05293_, _05292_, _05290_);
  and (_05294_, _05293_, _05288_);
  and (_05295_, _05274_, _04599_);
  and (_05296_, _05295_, \oc8051_golden_model_1.SCON [7]);
  and (_05297_, _05274_, _04623_);
  and (_05298_, _05297_, \oc8051_golden_model_1.IE [7]);
  nor (_05299_, _05298_, _05296_);
  and (_05300_, _05277_, _04599_);
  and (_05301_, _05300_, \oc8051_golden_model_1.P1 [7]);
  and (_05302_, _04613_, \oc8051_golden_model_1.P0 [7]);
  nor (_05303_, _05302_, _05301_);
  and (_05304_, _05303_, _05299_);
  and (_05305_, _05304_, _05294_);
  and (_05306_, _05305_, _05283_);
  and (_05307_, _05306_, _04586_);
  nor (_05308_, _05307_, _04639_);
  or (_05309_, _05308_, _05270_);
  not (_05310_, _03810_);
  not (_05311_, _03806_);
  and (_05312_, _02546_, \oc8051_golden_model_1.ACC [7]);
  and (_05313_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and (_05314_, _05313_, \oc8051_golden_model_1.PC [6]);
  and (_05315_, _05314_, _02618_);
  and (_05316_, _05315_, \oc8051_golden_model_1.PC [7]);
  nor (_05317_, _05315_, \oc8051_golden_model_1.PC [7]);
  nor (_05318_, _05317_, _05316_);
  and (_05319_, _05318_, _02804_);
  or (_05320_, _05319_, _05312_);
  not (_05321_, _04087_);
  and (_05322_, _02912_, _02798_);
  or (_05323_, _05322_, _04121_);
  nor (_05324_, _05323_, _03362_);
  and (_05325_, _05324_, _05321_);
  and (_05326_, _05325_, _05320_);
  not (_05327_, _05325_);
  and (_05328_, _05143_, _04839_);
  and (_05329_, _03989_, _03823_);
  and (_05330_, _04413_, _04226_);
  and (_05331_, _05330_, _05329_);
  and (_05332_, _05331_, _05328_);
  and (_05333_, _05332_, _04735_);
  or (_05334_, _05333_, _05198_);
  nand (_05335_, _05333_, _05198_);
  and (_05336_, _05335_, _05334_);
  and (_05337_, _05336_, _05327_);
  or (_05338_, _05337_, _05326_);
  and (_05339_, _05338_, _05311_);
  nor (_05340_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and (_05341_, _05340_, _03256_);
  nor (_05342_, _05341_, _03129_);
  nor (_05343_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and (_05344_, _05343_, _03129_);
  and (_05345_, _05344_, _02787_);
  nor (_05346_, _05345_, _05342_);
  nor (_05347_, _05346_, _03694_);
  not (_05348_, _05347_);
  not (_05349_, _03842_);
  nand (_05350_, _04226_, _05349_);
  not (_05351_, _03694_);
  nor (_05352_, _05349_, _02774_);
  nor (_05353_, _05352_, _05351_);
  nand (_05354_, _05353_, _05350_);
  and (_05355_, _05354_, _05348_);
  not (_05356_, _05355_);
  nor (_05357_, _05340_, _03256_);
  nor (_05358_, _05357_, _05341_);
  nor (_05359_, _05358_, _03694_);
  not (_05360_, _05359_);
  nand (_05361_, _04413_, _05349_);
  and (_05362_, _03842_, _03320_);
  nor (_05363_, _05362_, _05351_);
  nand (_05364_, _05363_, _05361_);
  and (_05365_, _05364_, _05360_);
  or (_05366_, _03805_, _03842_);
  and (_05367_, _03842_, _02835_);
  nor (_05368_, _05367_, _05351_);
  nand (_05369_, _05368_, _05366_);
  or (_05370_, _03694_, \oc8051_golden_model_1.SP [0]);
  and (_05371_, _05370_, _05369_);
  or (_05372_, _05371_, \oc8051_golden_model_1.IRAM[9] [7]);
  nor (_05373_, _03742_, _05349_);
  nor (_05374_, _03989_, _03842_);
  or (_05375_, _05374_, _05373_);
  nand (_05376_, _05375_, _03694_);
  nor (_05377_, _03927_, _03694_);
  not (_05378_, _05377_);
  and (_05379_, _05378_, _05376_);
  nand (_05380_, _05370_, _05369_);
  or (_05381_, _05380_, \oc8051_golden_model_1.IRAM[8] [7]);
  and (_05382_, _05381_, _05379_);
  and (_05383_, _05382_, _05372_);
  or (_05384_, _05380_, \oc8051_golden_model_1.IRAM[10] [7]);
  nand (_05385_, _05378_, _05376_);
  or (_05386_, _05371_, \oc8051_golden_model_1.IRAM[11] [7]);
  and (_05387_, _05386_, _05385_);
  and (_05388_, _05387_, _05384_);
  nor (_05389_, _05388_, _05383_);
  nand (_05390_, _05389_, _05365_);
  not (_05391_, _05365_);
  or (_05392_, _05371_, \oc8051_golden_model_1.IRAM[13] [7]);
  or (_05393_, _05380_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_05394_, _05393_, _05379_);
  and (_05395_, _05394_, _05392_);
  or (_05396_, _05380_, \oc8051_golden_model_1.IRAM[14] [7]);
  or (_05397_, _05371_, \oc8051_golden_model_1.IRAM[15] [7]);
  and (_05398_, _05397_, _05385_);
  and (_05399_, _05398_, _05396_);
  nor (_05400_, _05399_, _05395_);
  nand (_05401_, _05400_, _05391_);
  nand (_05402_, _05401_, _05390_);
  nand (_05403_, _05402_, _05356_);
  or (_05404_, _05380_, _04537_);
  or (_05405_, _05371_, _04535_);
  and (_05406_, _05405_, _05385_);
  nand (_05407_, _05406_, _05404_);
  or (_05408_, _05380_, _04529_);
  or (_05409_, _05371_, _04531_);
  and (_05410_, _05409_, _05379_);
  nand (_05411_, _05410_, _05408_);
  nand (_05412_, _05411_, _05407_);
  nand (_05413_, _05412_, _05365_);
  or (_05414_, _05380_, _04545_);
  or (_05415_, _05371_, _04543_);
  and (_05416_, _05415_, _05385_);
  nand (_05417_, _05416_, _05414_);
  or (_05418_, _05380_, _04549_);
  or (_05419_, _05371_, _04551_);
  and (_05420_, _05419_, _05379_);
  nand (_05421_, _05420_, _05418_);
  nand (_05422_, _05421_, _05417_);
  nand (_05423_, _05422_, _05391_);
  nand (_05424_, _05423_, _05413_);
  nand (_05425_, _05424_, _05355_);
  and (_05426_, _05425_, _05403_);
  and (_05427_, _05426_, _03806_);
  or (_05428_, _05427_, _05339_);
  and (_05429_, _05428_, _03992_);
  and (_05430_, _05189_, _04889_);
  not (_05431_, _05036_);
  and (_05432_, _05431_, _04987_);
  and (_05433_, _05085_, _04938_);
  and (_05434_, _05433_, _05432_);
  and (_05435_, _05434_, _05430_);
  and (_05436_, _05435_, _04783_);
  nor (_05437_, _05436_, _04690_);
  and (_05438_, _05436_, _04690_);
  nor (_05439_, _05438_, _05437_);
  and (_05440_, _05439_, _03811_);
  or (_05441_, _05440_, _05429_);
  and (_05442_, _05441_, _05310_);
  not (_05443_, _04639_);
  nand (_05444_, _05307_, _05443_);
  and (_05445_, _05444_, _03810_);
  or (_05446_, _05445_, _04239_);
  or (_05447_, _05446_, _05442_);
  nor (_05448_, _05318_, _02540_);
  nor (_05449_, _05448_, _03818_);
  and (_05450_, _05449_, _05447_);
  and (_05451_, _05198_, _03818_);
  or (_05452_, _05451_, _03827_);
  or (_05453_, _05452_, _05450_);
  and (_05454_, _05453_, _05309_);
  or (_05455_, _05454_, _02795_);
  and (_05456_, _04679_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05457_, _04681_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05458_, _05457_, _05456_);
  and (_05459_, _04673_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05460_, _04676_, \oc8051_golden_model_1.P1INREG [7]);
  nor (_05461_, _05460_, _05459_);
  and (_05462_, _05461_, _05458_);
  and (_05463_, _05462_, _04672_);
  and (_05464_, _05463_, _04666_);
  and (_05465_, _05464_, _04638_);
  and (_05466_, _05465_, _04586_);
  nand (_05467_, _05466_, _02795_);
  and (_05468_, _05467_, _02793_);
  and (_05469_, _05468_, _05455_);
  nor (_05470_, _05307_, _05443_);
  not (_05471_, _05470_);
  and (_05472_, _05471_, _05444_);
  and (_05473_, _05472_, _02792_);
  or (_05474_, _05473_, _05469_);
  and (_05475_, _05474_, _02533_);
  not (_05476_, _05318_);
  or (_05477_, _05476_, _02533_);
  nand (_05478_, _05477_, _02922_);
  or (_05479_, _05478_, _05475_);
  nand (_05480_, _05466_, _02923_);
  and (_05481_, _05480_, _05479_);
  or (_05482_, _05481_, _03842_);
  and (_05483_, _05426_, _02743_);
  nand (_05484_, _05465_, _03842_);
  or (_05485_, _05484_, _05483_);
  and (_05486_, _05485_, _04289_);
  and (_05487_, _05486_, _05482_);
  and (_05488_, _05280_, \oc8051_golden_model_1.P3INREG [7]);
  nor (_05489_, _05488_, _05276_);
  and (_05490_, _05489_, _05299_);
  and (_05491_, _05300_, \oc8051_golden_model_1.P1INREG [7]);
  not (_05492_, _05491_);
  and (_05493_, _04613_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05494_, _05278_, \oc8051_golden_model_1.P2INREG [7]);
  nor (_05495_, _05494_, _05493_);
  and (_05496_, _05495_, _05492_);
  and (_05497_, _05496_, _05490_);
  and (_05498_, _05497_, _05294_);
  and (_05499_, _05498_, _04586_);
  nor (_05500_, _05499_, _04639_);
  and (_05501_, _04639_, \oc8051_golden_model_1.PSW [7]);
  nor (_05502_, _05501_, _05500_);
  nor (_05503_, _05502_, _04289_);
  or (_05504_, _05503_, _02518_);
  or (_05505_, _05504_, _05487_);
  and (_05506_, _05476_, _02518_);
  nor (_05507_, _05506_, _03862_);
  and (_05508_, _05507_, _05505_);
  and (_05509_, _05198_, _03862_);
  or (_05510_, _05509_, _03851_);
  or (_05511_, _05510_, _05508_);
  not (_05512_, _03853_);
  or (_05513_, _05426_, _03852_);
  and (_05514_, _05513_, _05512_);
  and (_05515_, _05514_, _05511_);
  not (_05516_, _05267_);
  not (_05517_, _05256_);
  nor (_05518_, _05517_, _04585_);
  and (_05519_, _03043_, _01525_);
  and (_05520_, _03046_, _01531_);
  nor (_05521_, _05520_, _05519_);
  and (_05522_, _03034_, _01521_);
  and (_05523_, _03071_, _01517_);
  nor (_05524_, _05523_, _05522_);
  and (_05525_, _05524_, _05521_);
  and (_05526_, _03055_, _01556_);
  and (_05527_, _03057_, _01541_);
  nor (_05528_, _05527_, _05526_);
  and (_05529_, _03050_, _01533_);
  and (_05530_, _03075_, _01539_);
  nor (_05531_, _05530_, _05529_);
  and (_05532_, _05531_, _05528_);
  and (_05533_, _05532_, _05525_);
  and (_05534_, _03063_, _01548_);
  and (_05535_, _03066_, _01546_);
  nor (_05536_, _05535_, _05534_);
  and (_05537_, _03069_, _01559_);
  and (_05538_, _03037_, _01519_);
  nor (_05539_, _05538_, _05537_);
  and (_05540_, _05539_, _05536_);
  and (_05541_, _03052_, _01535_);
  and (_05542_, _03077_, _01554_);
  nor (_05543_, _05542_, _05541_);
  and (_05544_, _03080_, _01527_);
  and (_05545_, _03082_, _01550_);
  nor (_05546_, _05545_, _05544_);
  and (_05547_, _05546_, _05543_);
  and (_05548_, _05547_, _05540_);
  and (_05549_, _05548_, _05533_);
  and (_05550_, _05549_, _05517_);
  and (_05551_, _03080_, _01440_);
  and (_05552_, _03043_, _01437_);
  nor (_05553_, _05552_, _05551_);
  and (_05554_, _03050_, _01460_);
  and (_05555_, _03057_, _01429_);
  nor (_05556_, _05555_, _05554_);
  and (_05557_, _05556_, _05553_);
  and (_05558_, _03069_, _01435_);
  and (_05559_, _03046_, _01442_);
  nor (_05560_, _05559_, _05558_);
  and (_05561_, _03034_, _01447_);
  and (_05562_, _03066_, _01427_);
  nor (_05563_, _05562_, _05561_);
  and (_05564_, _05563_, _05560_);
  and (_05565_, _05564_, _05557_);
  and (_05566_, _03052_, _01462_);
  and (_05567_, _03075_, _01464_);
  nor (_05568_, _05567_, _05566_);
  and (_05569_, _03063_, _01425_);
  and (_05570_, _03077_, _01453_);
  nor (_05571_, _05570_, _05569_);
  and (_05572_, _05571_, _05568_);
  and (_05573_, _03071_, _01449_);
  and (_05574_, _03055_, _01455_);
  nor (_05575_, _05574_, _05573_);
  and (_05576_, _03037_, _01433_);
  and (_05577_, _03082_, _01458_);
  nor (_05578_, _05577_, _05576_);
  and (_05579_, _05578_, _05575_);
  and (_05580_, _05579_, _05572_);
  and (_05581_, _05580_, _05565_);
  and (_05582_, _03043_, _01483_);
  and (_05583_, _03046_, _01488_);
  nor (_05584_, _05583_, _05582_);
  and (_05585_, _03037_, _01479_);
  and (_05586_, _03071_, _01495_);
  nor (_05587_, _05586_, _05585_);
  and (_05588_, _05587_, _05584_);
  and (_05589_, _03055_, _01501_);
  and (_05590_, _03057_, _01475_);
  nor (_05591_, _05590_, _05589_);
  and (_05592_, _03050_, _01508_);
  and (_05593_, _03075_, _01511_);
  nor (_05594_, _05593_, _05592_);
  and (_05595_, _05594_, _05591_);
  and (_05596_, _05595_, _05588_);
  and (_05597_, _03080_, _01486_);
  and (_05598_, _03063_, _01471_);
  nor (_05599_, _05598_, _05597_);
  and (_05600_, _03069_, _01481_);
  and (_05601_, _03082_, _01504_);
  nor (_05602_, _05601_, _05600_);
  and (_05603_, _05602_, _05599_);
  and (_05604_, _03052_, _01506_);
  and (_05605_, _03077_, _01499_);
  nor (_05606_, _05605_, _05604_);
  and (_05607_, _03034_, _01493_);
  and (_05608_, _03066_, _01473_);
  nor (_05609_, _05608_, _05607_);
  and (_05610_, _05609_, _05606_);
  and (_05611_, _05610_, _05603_);
  and (_05612_, _05611_, _05596_);
  and (_05613_, _05612_, _05581_);
  and (_05614_, _05613_, _05550_);
  and (_05615_, _03660_, _03471_);
  not (_05616_, _03087_);
  and (_05617_, _03223_, _05616_);
  and (_05618_, _05617_, _05615_);
  and (_05619_, _05618_, _05614_);
  and (_05620_, _05619_, \oc8051_golden_model_1.TCON [7]);
  nor (_05621_, _05612_, _05581_);
  and (_05622_, _03223_, _03087_);
  and (_05623_, _05622_, _05615_);
  nor (_05624_, _05549_, _05256_);
  and (_05625_, _05624_, _05623_);
  and (_05626_, _05625_, _05621_);
  and (_05627_, _05626_, \oc8051_golden_model_1.B [7]);
  or (_05628_, _05627_, _05620_);
  not (_05629_, _05581_);
  and (_05630_, _05612_, _05629_);
  and (_05631_, _05630_, _05625_);
  and (_05632_, _05631_, \oc8051_golden_model_1.PSW [7]);
  not (_05633_, _05612_);
  and (_05634_, _05633_, _05581_);
  and (_05635_, _05634_, _05625_);
  and (_05636_, _05635_, \oc8051_golden_model_1.ACC [7]);
  or (_05637_, _05636_, _05632_);
  or (_05638_, _05637_, _05628_);
  and (_05639_, _05623_, _05614_);
  and (_05640_, _05639_, \oc8051_golden_model_1.P0INREG [7]);
  and (_05641_, _05630_, _05550_);
  and (_05642_, _05641_, _05618_);
  and (_05643_, _05642_, \oc8051_golden_model_1.SCON [7]);
  or (_05644_, _05643_, _05640_);
  and (_05645_, _05641_, _05623_);
  and (_05646_, _05645_, \oc8051_golden_model_1.P1INREG [7]);
  not (_05647_, _03471_);
  and (_05648_, _03660_, _05647_);
  and (_05649_, _05648_, _05617_);
  and (_05650_, _05649_, _05641_);
  and (_05651_, _05650_, \oc8051_golden_model_1.SBUF [7]);
  or (_05652_, _05651_, _05646_);
  or (_05653_, _05652_, _05644_);
  nor (_05654_, _03223_, _03087_);
  and (_05655_, _05654_, _05614_);
  and (_05656_, _05655_, _05648_);
  and (_05657_, _05656_, \oc8051_golden_model_1.TH1 [7]);
  and (_05658_, _05634_, _05550_);
  and (_05659_, _05658_, _05618_);
  and (_05660_, _05659_, \oc8051_golden_model_1.IE [7]);
  and (_05661_, _05621_, _05550_);
  and (_05662_, _05661_, _05623_);
  and (_05663_, _05662_, \oc8051_golden_model_1.P3INREG [7]);
  or (_05664_, _05663_, _05660_);
  and (_05665_, _05658_, _05623_);
  and (_05666_, _05665_, \oc8051_golden_model_1.P2INREG [7]);
  and (_05667_, _05661_, _05618_);
  and (_05668_, _05667_, \oc8051_golden_model_1.IP [7]);
  or (_05669_, _05668_, _05666_);
  or (_05670_, _05669_, _05664_);
  or (_05671_, _05670_, _05657_);
  or (_05672_, _05671_, _05653_);
  or (_05673_, _05672_, _05638_);
  and (_05674_, _05622_, _05614_);
  not (_05675_, _03660_);
  and (_05676_, _05675_, _03471_);
  and (_05677_, _05676_, _05674_);
  and (_05678_, _05677_, \oc8051_golden_model_1.DPL [7]);
  nor (_05679_, _03660_, _03471_);
  and (_05680_, _05679_, _05614_);
  and (_05681_, _05680_, _05622_);
  and (_05682_, _05681_, \oc8051_golden_model_1.DPH [7]);
  or (_05683_, _05682_, _05678_);
  and (_05684_, _05648_, _05674_);
  and (_05685_, _05684_, \oc8051_golden_model_1.SP [7]);
  and (_05686_, _05655_, _05615_);
  and (_05687_, _05686_, \oc8051_golden_model_1.TH0 [7]);
  or (_05688_, _05687_, _05685_);
  or (_05689_, _05688_, _05683_);
  not (_05690_, _03223_);
  and (_05691_, _05690_, _03087_);
  and (_05692_, _05691_, _05680_);
  and (_05693_, _05692_, \oc8051_golden_model_1.PCON [7]);
  and (_05694_, _05617_, _05614_);
  and (_05695_, _05648_, _05694_);
  and (_05696_, _05695_, \oc8051_golden_model_1.TMOD [7]);
  or (_05697_, _05696_, _05693_);
  and (_05698_, _05676_, _05694_);
  and (_05699_, _05698_, \oc8051_golden_model_1.TL0 [7]);
  and (_05700_, _05680_, _05617_);
  and (_05701_, _05700_, \oc8051_golden_model_1.TL1 [7]);
  or (_05702_, _05701_, _05699_);
  or (_05703_, _05702_, _05697_);
  or (_05704_, _05703_, _05689_);
  or (_05705_, _05704_, _05673_);
  or (_05706_, _05705_, _05518_);
  and (_05707_, _05706_, _03853_);
  or (_05708_, _05707_, _05516_);
  or (_05709_, _05708_, _05515_);
  and (_05710_, _05709_, _05269_);
  and (_05711_, _05517_, _03874_);
  or (_05712_, _05711_, _02585_);
  or (_05713_, _05712_, _05710_);
  and (_05714_, _05476_, _02585_);
  nor (_05715_, _05714_, _05225_);
  and (_05716_, _05715_, _05713_);
  or (_05717_, _05716_, _05260_);
  and (_05718_, _05717_, _05224_);
  not (_05719_, \oc8051_golden_model_1.ACC [7]);
  nor (_05720_, _04689_, _05719_);
  and (_05721_, _04689_, _05719_);
  nor (_05722_, _05721_, _05720_);
  and (_05723_, _05722_, _05223_);
  or (_05724_, _05723_, _05718_);
  and (_05725_, _05724_, _05222_);
  and (_05726_, _05258_, _05221_);
  or (_05727_, _05726_, _05725_);
  and (_05728_, _05727_, _05220_);
  and (_05729_, _05720_, _03880_);
  or (_05730_, _05729_, _02594_);
  or (_05731_, _05730_, _05728_);
  and (_05732_, _02994_, _02743_);
  and (_05733_, _05476_, _02594_);
  nor (_05734_, _05733_, _05732_);
  and (_05735_, _05734_, _05731_);
  and (_05736_, _03099_, _02743_);
  not (_05737_, _05732_);
  nor (_05738_, _05257_, _05737_);
  or (_05739_, _05738_, _05736_);
  or (_05740_, _05739_, _05735_);
  not (_05741_, _02592_);
  nand (_05742_, _05721_, _05736_);
  and (_05743_, _05742_, _05741_);
  and (_05744_, _05743_, _05740_);
  and (_05745_, _03011_, _02571_);
  nor (_05746_, _05745_, _03563_);
  nor (_05747_, _04060_, _03898_);
  and (_05748_, _05747_, _05746_);
  and (_05749_, _05318_, _02592_);
  nor (_05750_, _05749_, _04108_);
  nand (_05751_, _05750_, _05748_);
  or (_05752_, _05751_, _05744_);
  not (_05753_, _03898_);
  or (_05754_, _05371_, \oc8051_golden_model_1.IRAM[1] [6]);
  or (_05755_, _05380_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_05756_, _05755_, _05379_);
  and (_05757_, _05756_, _05754_);
  or (_05758_, _05380_, \oc8051_golden_model_1.IRAM[2] [6]);
  or (_05759_, _05371_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_05760_, _05759_, _05385_);
  and (_05761_, _05760_, _05758_);
  nor (_05762_, _05761_, _05757_);
  nand (_05763_, _05762_, _05365_);
  or (_05764_, _05371_, \oc8051_golden_model_1.IRAM[5] [6]);
  or (_05765_, _05380_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_05766_, _05765_, _05379_);
  and (_05767_, _05766_, _05764_);
  or (_05768_, _05380_, \oc8051_golden_model_1.IRAM[6] [6]);
  or (_05769_, _05371_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_05770_, _05769_, _05385_);
  and (_05771_, _05770_, _05768_);
  nor (_05772_, _05771_, _05767_);
  nand (_05773_, _05772_, _05391_);
  nand (_05774_, _05773_, _05763_);
  nand (_05775_, _05774_, _05355_);
  or (_05776_, _05380_, \oc8051_golden_model_1.IRAM[8] [6]);
  or (_05777_, _05371_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand (_05778_, _05777_, _05776_);
  nand (_05779_, _05778_, _05379_);
  or (_05780_, _05380_, \oc8051_golden_model_1.IRAM[10] [6]);
  or (_05781_, _05371_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand (_05782_, _05781_, _05780_);
  nand (_05783_, _05782_, _05385_);
  nand (_05784_, _05783_, _05779_);
  nand (_05785_, _05784_, _05365_);
  or (_05786_, _05380_, \oc8051_golden_model_1.IRAM[12] [6]);
  or (_05787_, _05371_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand (_05788_, _05787_, _05786_);
  nand (_05789_, _05788_, _05379_);
  or (_05790_, _05380_, \oc8051_golden_model_1.IRAM[14] [6]);
  or (_05791_, _05371_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand (_05792_, _05791_, _05790_);
  nand (_05793_, _05792_, _05385_);
  nand (_05794_, _05793_, _05789_);
  nand (_05795_, _05794_, _05391_);
  nand (_05796_, _05795_, _05785_);
  nand (_05797_, _05796_, _05356_);
  and (_05798_, _05797_, _05775_);
  not (_05799_, _05798_);
  or (_05800_, _05371_, \oc8051_golden_model_1.IRAM[1] [1]);
  or (_05801_, _05380_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_05802_, _05801_, _05379_);
  and (_05803_, _05802_, _05800_);
  or (_05804_, _05380_, \oc8051_golden_model_1.IRAM[2] [1]);
  or (_05805_, _05371_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_05806_, _05805_, _05385_);
  and (_05807_, _05806_, _05804_);
  nor (_05808_, _05807_, _05803_);
  nand (_05809_, _05808_, _05365_);
  or (_05810_, _05371_, _03945_);
  or (_05811_, _05380_, _03947_);
  nand (_05812_, _05811_, _05810_);
  nand (_05813_, _05812_, _05385_);
  or (_05814_, _05371_, _03953_);
  or (_05815_, _05380_, _03951_);
  nand (_05816_, _05815_, _05814_);
  nand (_05817_, _05816_, _05379_);
  and (_05818_, _05817_, _05813_);
  nand (_05819_, _05818_, _05391_);
  and (_05820_, _05819_, _05355_);
  nand (_05821_, _05820_, _05809_);
  or (_05822_, _05380_, \oc8051_golden_model_1.IRAM[12] [1]);
  or (_05823_, _05371_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand (_05824_, _05823_, _05822_);
  nand (_05825_, _05824_, _05379_);
  or (_05826_, _05380_, \oc8051_golden_model_1.IRAM[14] [1]);
  or (_05827_, _05371_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand (_05828_, _05827_, _05826_);
  nand (_05829_, _05828_, _05385_);
  nand (_05830_, _05829_, _05825_);
  nand (_05831_, _05830_, _05391_);
  or (_05832_, _05380_, \oc8051_golden_model_1.IRAM[8] [1]);
  or (_05833_, _05371_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand (_05834_, _05833_, _05832_);
  nand (_05835_, _05834_, _05379_);
  or (_05836_, _05380_, \oc8051_golden_model_1.IRAM[10] [1]);
  or (_05837_, _05371_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand (_05838_, _05837_, _05836_);
  nand (_05839_, _05838_, _05385_);
  nand (_05840_, _05839_, _05835_);
  nand (_05841_, _05840_, _05365_);
  and (_05842_, _05841_, _05356_);
  nand (_05843_, _05842_, _05831_);
  and (_05844_, _05843_, _05821_);
  or (_05845_, _05371_, \oc8051_golden_model_1.IRAM[1] [0]);
  or (_05846_, _05380_, \oc8051_golden_model_1.IRAM[0] [0]);
  and (_05847_, _05846_, _05379_);
  and (_05848_, _05847_, _05845_);
  or (_05849_, _05380_, \oc8051_golden_model_1.IRAM[2] [0]);
  or (_05850_, _05371_, \oc8051_golden_model_1.IRAM[3] [0]);
  and (_05851_, _05850_, _05385_);
  and (_05852_, _05851_, _05849_);
  nor (_05853_, _05852_, _05848_);
  nand (_05854_, _05853_, _05365_);
  or (_05855_, _05371_, _03762_);
  or (_05856_, _05380_, _03764_);
  nand (_05857_, _05856_, _05855_);
  nand (_05858_, _05857_, _05385_);
  or (_05859_, _05371_, _03770_);
  or (_05860_, _05380_, _03768_);
  nand (_05861_, _05860_, _05859_);
  nand (_05862_, _05861_, _05379_);
  and (_05863_, _05862_, _05858_);
  nand (_05864_, _05863_, _05391_);
  and (_05865_, _05864_, _05355_);
  nand (_05866_, _05865_, _05854_);
  or (_05867_, _05380_, \oc8051_golden_model_1.IRAM[12] [0]);
  or (_05868_, _05371_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand (_05869_, _05868_, _05867_);
  nand (_05870_, _05869_, _05379_);
  or (_05871_, _05380_, \oc8051_golden_model_1.IRAM[14] [0]);
  or (_05872_, _05371_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand (_05873_, _05872_, _05871_);
  nand (_05874_, _05873_, _05385_);
  nand (_05875_, _05874_, _05870_);
  nand (_05876_, _05875_, _05391_);
  or (_05877_, _05380_, \oc8051_golden_model_1.IRAM[8] [0]);
  or (_05878_, _05371_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand (_05879_, _05878_, _05877_);
  nand (_05880_, _05879_, _05379_);
  or (_05881_, _05380_, \oc8051_golden_model_1.IRAM[10] [0]);
  or (_05882_, _05371_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand (_05883_, _05882_, _05881_);
  nand (_05884_, _05883_, _05385_);
  nand (_05885_, _05884_, _05880_);
  nand (_05886_, _05885_, _05365_);
  and (_05887_, _05886_, _05356_);
  nand (_05888_, _05887_, _05876_);
  and (_05889_, _05888_, _05866_);
  and (_05890_, _05889_, _05844_);
  or (_05891_, _05371_, \oc8051_golden_model_1.IRAM[1] [3]);
  or (_05892_, _05380_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_05893_, _05892_, _05379_);
  and (_05894_, _05893_, _05891_);
  or (_05895_, _05380_, \oc8051_golden_model_1.IRAM[2] [3]);
  or (_05896_, _05371_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_05897_, _05896_, _05385_);
  and (_05898_, _05897_, _05895_);
  nor (_05899_, _05898_, _05894_);
  nand (_05900_, _05899_, _05365_);
  or (_05901_, _05371_, _04187_);
  or (_05902_, _05380_, _04189_);
  nand (_05903_, _05902_, _05901_);
  nand (_05904_, _05903_, _05385_);
  or (_05905_, _05371_, _04195_);
  or (_05906_, _05380_, _04193_);
  nand (_05907_, _05906_, _05905_);
  nand (_05908_, _05907_, _05379_);
  and (_05909_, _05908_, _05904_);
  nand (_05910_, _05909_, _05391_);
  and (_05911_, _05910_, _05355_);
  nand (_05912_, _05911_, _05900_);
  or (_05913_, _05380_, \oc8051_golden_model_1.IRAM[12] [3]);
  or (_05914_, _05371_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand (_05915_, _05914_, _05913_);
  nand (_05916_, _05915_, _05379_);
  or (_05917_, _05380_, \oc8051_golden_model_1.IRAM[14] [3]);
  or (_05918_, _05371_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand (_05919_, _05918_, _05917_);
  nand (_05920_, _05919_, _05385_);
  nand (_05921_, _05920_, _05916_);
  nand (_05922_, _05921_, _05391_);
  or (_05923_, _05380_, \oc8051_golden_model_1.IRAM[8] [3]);
  or (_05924_, _05371_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand (_05925_, _05924_, _05923_);
  nand (_05926_, _05925_, _05379_);
  or (_05927_, _05380_, \oc8051_golden_model_1.IRAM[10] [3]);
  or (_05928_, _05371_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand (_05929_, _05928_, _05927_);
  nand (_05930_, _05929_, _05385_);
  nand (_05931_, _05930_, _05926_);
  nand (_05932_, _05931_, _05365_);
  and (_05933_, _05932_, _05356_);
  nand (_05934_, _05933_, _05922_);
  and (_05935_, _05934_, _05912_);
  or (_05936_, _05371_, \oc8051_golden_model_1.IRAM[1] [2]);
  or (_05937_, _05380_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_05938_, _05937_, _05379_);
  and (_05939_, _05938_, _05936_);
  or (_05940_, _05380_, \oc8051_golden_model_1.IRAM[2] [2]);
  or (_05941_, _05371_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_05942_, _05941_, _05385_);
  and (_05943_, _05942_, _05940_);
  nor (_05944_, _05943_, _05939_);
  nand (_05945_, _05944_, _05365_);
  or (_05946_, _05371_, _04371_);
  or (_05947_, _05380_, _04373_);
  nand (_05948_, _05947_, _05946_);
  nand (_05949_, _05948_, _05385_);
  or (_05950_, _05371_, _04379_);
  or (_05951_, _05380_, _04377_);
  nand (_05952_, _05951_, _05950_);
  nand (_05953_, _05952_, _05379_);
  and (_05954_, _05953_, _05949_);
  nand (_05955_, _05954_, _05391_);
  and (_05956_, _05955_, _05355_);
  nand (_05957_, _05956_, _05945_);
  or (_05958_, _05380_, \oc8051_golden_model_1.IRAM[12] [2]);
  or (_05959_, _05371_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand (_05960_, _05959_, _05958_);
  nand (_05961_, _05960_, _05379_);
  or (_05962_, _05380_, \oc8051_golden_model_1.IRAM[14] [2]);
  or (_05963_, _05371_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand (_05964_, _05963_, _05962_);
  nand (_05965_, _05964_, _05385_);
  nand (_05966_, _05965_, _05961_);
  nand (_05967_, _05966_, _05391_);
  or (_05968_, _05380_, \oc8051_golden_model_1.IRAM[8] [2]);
  or (_05969_, _05371_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand (_05970_, _05969_, _05968_);
  nand (_05971_, _05970_, _05379_);
  or (_05972_, _05380_, \oc8051_golden_model_1.IRAM[10] [2]);
  or (_05973_, _05371_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand (_05974_, _05973_, _05972_);
  nand (_05975_, _05974_, _05385_);
  nand (_05976_, _05975_, _05971_);
  nand (_05977_, _05976_, _05365_);
  and (_05978_, _05977_, _05356_);
  nand (_05979_, _05978_, _05967_);
  and (_05980_, _05979_, _05957_);
  and (_05981_, _05980_, _05935_);
  and (_05982_, _05981_, _05890_);
  or (_05983_, _05371_, \oc8051_golden_model_1.IRAM[1] [5]);
  or (_05984_, _05380_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_05985_, _05984_, _05379_);
  and (_05986_, _05985_, _05983_);
  or (_05987_, _05380_, \oc8051_golden_model_1.IRAM[2] [5]);
  or (_05988_, _05371_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_05989_, _05988_, _05385_);
  and (_05990_, _05989_, _05987_);
  nor (_05991_, _05990_, _05986_);
  nand (_05992_, _05991_, _05365_);
  or (_05993_, _05371_, _04797_);
  or (_05994_, _05380_, _04799_);
  nand (_05995_, _05994_, _05993_);
  nand (_05996_, _05995_, _05385_);
  or (_05997_, _05371_, _04805_);
  or (_05998_, _05380_, _04803_);
  nand (_05999_, _05998_, _05997_);
  nand (_06000_, _05999_, _05379_);
  and (_06001_, _06000_, _05996_);
  nand (_06002_, _06001_, _05391_);
  and (_06003_, _06002_, _05355_);
  nand (_06004_, _06003_, _05992_);
  or (_06005_, _05380_, \oc8051_golden_model_1.IRAM[12] [5]);
  or (_06006_, _05371_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand (_06007_, _06006_, _06005_);
  nand (_06008_, _06007_, _05379_);
  or (_06009_, _05380_, \oc8051_golden_model_1.IRAM[14] [5]);
  or (_06010_, _05371_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand (_06011_, _06010_, _06009_);
  nand (_06012_, _06011_, _05385_);
  nand (_06013_, _06012_, _06008_);
  nand (_06014_, _06013_, _05391_);
  or (_06015_, _05380_, \oc8051_golden_model_1.IRAM[8] [5]);
  or (_06016_, _05371_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand (_06017_, _06016_, _06015_);
  nand (_06018_, _06017_, _05379_);
  or (_06019_, _05380_, \oc8051_golden_model_1.IRAM[10] [5]);
  or (_06020_, _05371_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand (_06021_, _06020_, _06019_);
  nand (_06022_, _06021_, _05385_);
  nand (_06023_, _06022_, _06018_);
  nand (_06024_, _06023_, _05365_);
  and (_06025_, _06024_, _05356_);
  nand (_06026_, _06025_, _06014_);
  and (_06027_, _06026_, _06004_);
  or (_06028_, _05371_, \oc8051_golden_model_1.IRAM[1] [4]);
  or (_06029_, _05380_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_06030_, _06029_, _05379_);
  and (_06031_, _06030_, _06028_);
  or (_06032_, _05380_, \oc8051_golden_model_1.IRAM[2] [4]);
  or (_06033_, _05371_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_06034_, _06033_, _05385_);
  and (_06035_, _06034_, _06032_);
  nor (_06036_, _06035_, _06031_);
  nand (_06037_, _06036_, _05365_);
  or (_06038_, _05371_, _05101_);
  or (_06039_, _05380_, _05103_);
  nand (_06040_, _06039_, _06038_);
  nand (_06041_, _06040_, _05385_);
  or (_06042_, _05371_, _05109_);
  or (_06043_, _05380_, _05107_);
  nand (_06044_, _06043_, _06042_);
  nand (_06045_, _06044_, _05379_);
  and (_06046_, _06045_, _06041_);
  nand (_06047_, _06046_, _05391_);
  and (_06048_, _06047_, _05355_);
  nand (_06049_, _06048_, _06037_);
  or (_06050_, _05380_, \oc8051_golden_model_1.IRAM[12] [4]);
  or (_06051_, _05371_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand (_06052_, _06051_, _06050_);
  nand (_06053_, _06052_, _05379_);
  or (_06054_, _05380_, \oc8051_golden_model_1.IRAM[14] [4]);
  or (_06055_, _05371_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand (_06056_, _06055_, _06054_);
  nand (_06057_, _06056_, _05385_);
  nand (_06058_, _06057_, _06053_);
  nand (_06059_, _06058_, _05391_);
  or (_06060_, _05380_, \oc8051_golden_model_1.IRAM[8] [4]);
  or (_06061_, _05371_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand (_06062_, _06061_, _06060_);
  nand (_06063_, _06062_, _05379_);
  or (_06064_, _05380_, \oc8051_golden_model_1.IRAM[10] [4]);
  or (_06065_, _05371_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand (_06066_, _06065_, _06064_);
  nand (_06067_, _06066_, _05385_);
  nand (_06068_, _06067_, _06063_);
  nand (_06069_, _06068_, _05365_);
  and (_06070_, _06069_, _05356_);
  nand (_06071_, _06070_, _06059_);
  and (_06072_, _06071_, _06049_);
  and (_06073_, _06072_, _06027_);
  and (_06074_, _06073_, _05982_);
  and (_06075_, _06074_, _05799_);
  or (_06076_, _06075_, _05426_);
  nand (_06077_, _06075_, _05426_);
  and (_06078_, _06077_, _06076_);
  or (_06079_, _06078_, _05753_);
  not (_06080_, _03900_);
  and (_06081_, _03009_, _02571_);
  nor (_06082_, _06081_, _04108_);
  nor (_06083_, _05745_, _03228_);
  nand (_06084_, _06083_, _06082_);
  nor (_06085_, _06084_, _03557_);
  or (_06086_, _06085_, _05336_);
  and (_06087_, _06086_, _06080_);
  and (_06088_, _06087_, _06079_);
  and (_06089_, _06088_, _05752_);
  and (_06090_, _05439_, _03900_);
  or (_06091_, _06090_, _06089_);
  and (_06092_, _06091_, _05219_);
  and (_06093_, _02229_, \oc8051_golden_model_1.PC [2]);
  and (_06094_, _06093_, \oc8051_golden_model_1.PC [3]);
  and (_06095_, _06094_, _05314_);
  and (_06096_, _06095_, \oc8051_golden_model_1.PC [7]);
  nor (_06097_, _06095_, \oc8051_golden_model_1.PC [7]);
  nor (_06098_, _06097_, _06096_);
  and (_06099_, _06098_, _02988_);
  or (_06100_, _06099_, _06092_);
  and (_06101_, _06100_, _05218_);
  and (_06102_, _05318_, _02572_);
  or (_06103_, _06102_, _06101_);
  and (_06104_, _06103_, _02781_);
  not (_06105_, _05216_);
  and (_06106_, _05500_, _02780_);
  nor (_06107_, _06106_, _06105_);
  not (_06108_, _06107_);
  nor (_06109_, _06108_, _06104_);
  nor (_06110_, _06109_, _05217_);
  nor (_06111_, _06110_, _03912_);
  not (_06112_, _03912_);
  nand (_06113_, _05843_, _05821_);
  nand (_06114_, _05888_, _05866_);
  and (_06115_, _06114_, _06113_);
  nand (_06116_, _05934_, _05912_);
  nand (_06117_, _05979_, _05957_);
  and (_06118_, _06117_, _06116_);
  and (_06119_, _06118_, _06115_);
  nand (_06120_, _06026_, _06004_);
  nand (_06121_, _06071_, _06049_);
  and (_06122_, _06121_, _06120_);
  and (_06123_, _06122_, _06119_);
  and (_06124_, _06123_, _05798_);
  and (_06125_, _06124_, _05426_);
  nor (_06126_, _06124_, _05426_);
  nor (_06127_, _06126_, _06125_);
  nor (_06128_, _06127_, _06112_);
  nor (_06129_, _06128_, _03914_);
  not (_06130_, _06129_);
  nor (_06131_, _06130_, _06111_);
  nor (_06132_, _06131_, _05197_);
  nor (_06133_, _06132_, _04520_);
  or (_06134_, _06133_, _04528_);
  and (_06135_, _06134_, _04518_);
  and (_06136_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and (_06137_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and (_06138_, _06137_, _06136_);
  and (_06139_, _06138_, _06096_);
  and (_06140_, _06139_, \oc8051_golden_model_1.PC [12]);
  and (_06141_, _06140_, \oc8051_golden_model_1.PC [13]);
  and (_06142_, _06141_, \oc8051_golden_model_1.PC [14]);
  nor (_06143_, _06142_, \oc8051_golden_model_1.PC [15]);
  and (_06144_, _06142_, \oc8051_golden_model_1.PC [15]);
  nor (_06145_, _06144_, _06143_);
  not (_06146_, _06145_);
  nand (_06147_, _06146_, _02988_);
  and (_06148_, _06138_, _05316_);
  and (_06149_, _06148_, \oc8051_golden_model_1.PC [12]);
  and (_06150_, _06149_, \oc8051_golden_model_1.PC [13]);
  and (_06151_, _06150_, \oc8051_golden_model_1.PC [14]);
  nor (_06152_, _06151_, \oc8051_golden_model_1.PC [15]);
  and (_06153_, _06151_, \oc8051_golden_model_1.PC [15]);
  nor (_06154_, _06153_, _06152_);
  or (_06155_, _06154_, _02988_);
  and (_06156_, _06155_, _06147_);
  and (_06157_, _06156_, _04513_);
  and (_06158_, _06157_, _04516_);
  or (_35698_, _06158_, _06135_);
  not (_06159_, \oc8051_golden_model_1.B [7]);
  nor (_06160_, _34446_, _06159_);
  not (_06161_, _03094_);
  not (_06162_, _02932_);
  nor (_06163_, _04661_, _06159_);
  and (_06164_, _05439_, _04661_);
  or (_06165_, _06164_, _06163_);
  or (_06166_, _06165_, _06162_);
  and (_06167_, _04661_, \oc8051_golden_model_1.ACC [7]);
  or (_06168_, _06167_, _06163_);
  and (_06169_, _06168_, _02837_);
  nor (_06170_, _02837_, _06159_);
  or (_06171_, _06170_, _02932_);
  or (_06172_, _06171_, _06169_);
  and (_06173_, _06172_, _02939_);
  and (_06174_, _06173_, _06166_);
  not (_06175_, _04661_);
  nor (_06176_, _06175_, _04585_);
  or (_06177_, _06176_, _06163_);
  and (_06178_, _06177_, _02930_);
  nor (_06179_, _05286_, _06159_);
  and (_06180_, _05444_, _05286_);
  or (_06181_, _06180_, _06179_);
  and (_06182_, _06181_, _02799_);
  or (_06183_, _06182_, _06178_);
  or (_06184_, _06183_, _02928_);
  or (_06185_, _06184_, _06174_);
  or (_06186_, _06168_, _02943_);
  and (_06187_, _06186_, _06185_);
  or (_06188_, _06187_, _02796_);
  not (_06189_, _02790_);
  and (_06190_, _05308_, _05286_);
  or (_06191_, _06190_, _06179_);
  or (_06192_, _06191_, _02927_);
  and (_06193_, _06192_, _06189_);
  and (_06194_, _06193_, _06188_);
  and (_06195_, _02978_, _02900_);
  or (_06196_, _06179_, _05471_);
  and (_06197_, _06196_, _02790_);
  and (_06198_, _06197_, _06181_);
  or (_06199_, _06198_, _06195_);
  or (_06200_, _06199_, _06194_);
  not (_06201_, _06195_);
  and (_06202_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and (_06203_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and (_06204_, _06203_, _06202_);
  and (_06205_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [5]);
  and (_06206_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  and (_06207_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor (_06208_, _06207_, _06206_);
  nor (_06209_, _06208_, _06204_);
  and (_06210_, _06209_, _06205_);
  nor (_06211_, _06210_, _06204_);
  and (_06212_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and (_06213_, _06212_, _06207_);
  and (_06214_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor (_06215_, _06214_, _06202_);
  nor (_06216_, _06215_, _06213_);
  not (_06217_, _06216_);
  nor (_06218_, _06217_, _06211_);
  and (_06219_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and (_06220_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [5]);
  and (_06221_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [4]);
  and (_06222_, _06221_, _06220_);
  nor (_06223_, _06221_, _06220_);
  nor (_06224_, _06223_, _06222_);
  and (_06225_, _06224_, _06219_);
  nor (_06226_, _06224_, _06219_);
  nor (_06227_, _06226_, _06225_);
  and (_06228_, _06217_, _06211_);
  nor (_06229_, _06228_, _06218_);
  and (_06230_, _06229_, _06227_);
  nor (_06231_, _06230_, _06218_);
  not (_06232_, _06207_);
  and (_06233_, _06212_, _06232_);
  and (_06234_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [4]);
  and (_06235_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and (_06236_, _06235_, _06220_);
  and (_06237_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [5]);
  and (_06238_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor (_06239_, _06238_, _06237_);
  nor (_06240_, _06239_, _06236_);
  and (_06241_, _06240_, _06234_);
  nor (_06242_, _06240_, _06234_);
  nor (_06243_, _06242_, _06241_);
  and (_06244_, _06243_, _06233_);
  nor (_06245_, _06243_, _06233_);
  nor (_06246_, _06245_, _06244_);
  not (_06247_, _06246_);
  nor (_06248_, _06247_, _06231_);
  and (_06249_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and (_06250_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [1]);
  and (_06251_, _06250_, _06249_);
  nor (_06252_, _06225_, _06222_);
  and (_06253_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [2]);
  and (_06254_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and (_06255_, _06254_, _06253_);
  nor (_06256_, _06254_, _06253_);
  nor (_06257_, _06256_, _06255_);
  not (_06258_, _06257_);
  nor (_06259_, _06258_, _06252_);
  and (_06260_, _06258_, _06252_);
  nor (_06261_, _06260_, _06259_);
  and (_06262_, _06261_, _06251_);
  nor (_06263_, _06261_, _06251_);
  nor (_06264_, _06263_, _06262_);
  and (_06265_, _06247_, _06231_);
  nor (_06266_, _06265_, _06248_);
  and (_06267_, _06266_, _06264_);
  nor (_06268_, _06267_, _06248_);
  nor (_06269_, _06241_, _06236_);
  and (_06270_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [3]);
  and (_06271_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [4]);
  and (_06272_, _06271_, _06270_);
  nor (_06273_, _06271_, _06270_);
  nor (_06274_, _06273_, _06272_);
  not (_06275_, _06274_);
  nor (_06276_, _06275_, _06269_);
  and (_06277_, _06275_, _06269_);
  nor (_06278_, _06277_, _06276_);
  and (_06279_, _06278_, _06255_);
  nor (_06280_, _06278_, _06255_);
  nor (_06281_, _06280_, _06279_);
  nor (_06282_, _06244_, _06213_);
  and (_06283_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [5]);
  and (_06284_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and (_06285_, _06284_, _06235_);
  nor (_06286_, _06284_, _06235_);
  nor (_06287_, _06286_, _06285_);
  and (_06288_, _06287_, _06283_);
  nor (_06289_, _06287_, _06283_);
  nor (_06290_, _06289_, _06288_);
  not (_06291_, _06290_);
  nor (_06292_, _06291_, _06282_);
  and (_06293_, _06291_, _06282_);
  nor (_06294_, _06293_, _06292_);
  and (_06295_, _06294_, _06281_);
  nor (_06296_, _06294_, _06281_);
  nor (_06297_, _06296_, _06295_);
  not (_06298_, _06297_);
  nor (_06299_, _06298_, _06268_);
  nor (_06300_, _06262_, _06259_);
  not (_06301_, _06300_);
  and (_06302_, _06298_, _06268_);
  nor (_06303_, _06302_, _06299_);
  and (_06304_, _06303_, _06301_);
  nor (_06305_, _06304_, _06299_);
  nor (_06306_, _06279_, _06276_);
  not (_06307_, _06306_);
  nor (_06308_, _06295_, _06292_);
  not (_06309_, _06308_);
  and (_06310_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and (_06311_, _06310_, _06235_);
  and (_06312_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and (_06313_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor (_06314_, _06313_, _06312_);
  nor (_06315_, _06314_, _06311_);
  nor (_06316_, _06288_, _06285_);
  and (_06317_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [4]);
  and (_06318_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [5]);
  and (_06319_, _06318_, _06317_);
  nor (_06320_, _06318_, _06317_);
  nor (_06321_, _06320_, _06319_);
  not (_06322_, _06321_);
  nor (_06323_, _06322_, _06316_);
  and (_06324_, _06322_, _06316_);
  nor (_06325_, _06324_, _06323_);
  and (_06326_, _06325_, _06272_);
  nor (_06327_, _06325_, _06272_);
  nor (_06328_, _06327_, _06326_);
  and (_06329_, _06328_, _06315_);
  nor (_06330_, _06328_, _06315_);
  nor (_06331_, _06330_, _06329_);
  and (_06332_, _06331_, _06309_);
  nor (_06333_, _06331_, _06309_);
  nor (_06334_, _06333_, _06332_);
  and (_06335_, _06334_, _06307_);
  nor (_06336_, _06334_, _06307_);
  nor (_06337_, _06336_, _06335_);
  not (_06338_, _06337_);
  nor (_06339_, _06338_, _06305_);
  nor (_06340_, _06335_, _06332_);
  nor (_06341_, _06326_, _06323_);
  not (_06342_, _06341_);
  and (_06343_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [5]);
  and (_06344_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and (_06345_, _06344_, _06343_);
  nor (_06346_, _06344_, _06343_);
  nor (_06347_, _06346_, _06345_);
  and (_06348_, _06347_, _06311_);
  nor (_06349_, _06347_, _06311_);
  nor (_06350_, _06349_, _06348_);
  and (_06351_, _06350_, _06319_);
  nor (_06352_, _06350_, _06319_);
  nor (_06353_, _06352_, _06351_);
  and (_06354_, _06353_, _06310_);
  nor (_06355_, _06353_, _06310_);
  nor (_06356_, _06355_, _06354_);
  and (_06357_, _06356_, _06329_);
  nor (_06358_, _06356_, _06329_);
  nor (_06359_, _06358_, _06357_);
  and (_06360_, _06359_, _06342_);
  nor (_06361_, _06359_, _06342_);
  nor (_06362_, _06361_, _06360_);
  not (_06363_, _06362_);
  nor (_06364_, _06363_, _06340_);
  and (_06365_, _06363_, _06340_);
  nor (_06366_, _06365_, _06364_);
  and (_06367_, _06366_, _06339_);
  nor (_06368_, _06360_, _06357_);
  nor (_06369_, _06351_, _06348_);
  not (_06370_, _06369_);
  and (_06371_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [6]);
  and (_06372_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and (_06373_, _06372_, _06371_);
  nor (_06374_, _06372_, _06371_);
  nor (_06375_, _06374_, _06373_);
  and (_06376_, _06375_, _06345_);
  nor (_06377_, _06375_, _06345_);
  nor (_06378_, _06377_, _06376_);
  and (_06379_, _06378_, _06354_);
  nor (_06380_, _06378_, _06354_);
  nor (_06381_, _06380_, _06379_);
  and (_06382_, _06381_, _06370_);
  nor (_06383_, _06381_, _06370_);
  nor (_06384_, _06383_, _06382_);
  not (_06385_, _06384_);
  nor (_06386_, _06385_, _06368_);
  and (_06387_, _06385_, _06368_);
  nor (_06388_, _06387_, _06386_);
  and (_06389_, _06388_, _06364_);
  nor (_06390_, _06388_, _06364_);
  nor (_06391_, _06390_, _06389_);
  and (_06392_, _06391_, _06367_);
  nor (_06393_, _06391_, _06367_);
  nor (_06394_, _06393_, _06392_);
  and (_06395_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  and (_06396_, _06395_, _06207_);
  and (_06397_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [4]);
  and (_06398_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [5]);
  nor (_06399_, _06398_, _06203_);
  nor (_06400_, _06399_, _06396_);
  and (_06401_, _06400_, _06397_);
  nor (_06402_, _06401_, _06396_);
  not (_06403_, _06402_);
  nor (_06404_, _06209_, _06205_);
  nor (_06405_, _06404_, _06210_);
  and (_06406_, _06405_, _06403_);
  and (_06407_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and (_06408_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [4]);
  and (_06409_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and (_06410_, _06409_, _06408_);
  nor (_06411_, _06409_, _06408_);
  nor (_06412_, _06411_, _06410_);
  and (_06413_, _06412_, _06407_);
  nor (_06414_, _06412_, _06407_);
  nor (_06415_, _06414_, _06413_);
  nor (_06416_, _06405_, _06403_);
  nor (_06417_, _06416_, _06406_);
  and (_06418_, _06417_, _06415_);
  nor (_06419_, _06418_, _06406_);
  nor (_06420_, _06229_, _06227_);
  nor (_06421_, _06420_, _06230_);
  not (_06422_, _06421_);
  nor (_06423_, _06422_, _06419_);
  and (_06424_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and (_06425_, _06424_, _06250_);
  nor (_06426_, _06413_, _06410_);
  nor (_06427_, _06250_, _06249_);
  nor (_06428_, _06427_, _06251_);
  not (_06429_, _06428_);
  nor (_06430_, _06429_, _06426_);
  and (_06431_, _06429_, _06426_);
  nor (_06432_, _06431_, _06430_);
  and (_06433_, _06432_, _06425_);
  nor (_06434_, _06432_, _06425_);
  nor (_06435_, _06434_, _06433_);
  and (_06436_, _06422_, _06419_);
  nor (_06437_, _06436_, _06423_);
  and (_06438_, _06437_, _06435_);
  nor (_06439_, _06438_, _06423_);
  nor (_06440_, _06266_, _06264_);
  nor (_06441_, _06440_, _06267_);
  not (_06442_, _06441_);
  nor (_06443_, _06442_, _06439_);
  nor (_06444_, _06433_, _06430_);
  not (_06445_, _06444_);
  and (_06446_, _06442_, _06439_);
  nor (_06447_, _06446_, _06443_);
  and (_06448_, _06447_, _06445_);
  nor (_06449_, _06448_, _06443_);
  nor (_06450_, _06303_, _06301_);
  nor (_06451_, _06450_, _06304_);
  not (_06452_, _06451_);
  nor (_06453_, _06452_, _06449_);
  and (_06454_, _06338_, _06305_);
  nor (_06455_, _06454_, _06339_);
  and (_06456_, _06455_, _06453_);
  nor (_06457_, _06366_, _06339_);
  nor (_06458_, _06457_, _06367_);
  and (_06459_, _06458_, _06456_);
  and (_06460_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [4]);
  and (_06461_, _06460_, _06395_);
  and (_06462_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor (_06463_, _06460_, _06395_);
  nor (_06464_, _06463_, _06461_);
  and (_06465_, _06464_, _06462_);
  nor (_06466_, _06465_, _06461_);
  not (_06467_, _06466_);
  nor (_06468_, _06400_, _06397_);
  nor (_06469_, _06468_, _06401_);
  and (_06470_, _06469_, _06467_);
  and (_06471_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [1]);
  and (_06472_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and (_06473_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and (_06474_, _06473_, _06472_);
  nor (_06475_, _06473_, _06472_);
  nor (_06476_, _06475_, _06474_);
  and (_06477_, _06476_, _06471_);
  nor (_06478_, _06476_, _06471_);
  nor (_06479_, _06478_, _06477_);
  nor (_06480_, _06469_, _06467_);
  nor (_06481_, _06480_, _06470_);
  and (_06482_, _06481_, _06479_);
  nor (_06483_, _06482_, _06470_);
  not (_06484_, _06483_);
  nor (_06485_, _06417_, _06415_);
  nor (_06486_, _06485_, _06418_);
  and (_06487_, _06486_, _06484_);
  nor (_06488_, _06477_, _06474_);
  and (_06489_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [1]);
  and (_06490_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [0]);
  nor (_06491_, _06490_, _06489_);
  nor (_06492_, _06491_, _06425_);
  not (_06493_, _06492_);
  nor (_06494_, _06493_, _06488_);
  and (_06495_, _06493_, _06488_);
  nor (_06496_, _06495_, _06494_);
  nor (_06497_, _06486_, _06484_);
  nor (_06498_, _06497_, _06487_);
  and (_06499_, _06498_, _06496_);
  nor (_06500_, _06499_, _06487_);
  nor (_06501_, _06437_, _06435_);
  nor (_06502_, _06501_, _06438_);
  not (_06503_, _06502_);
  nor (_06504_, _06503_, _06500_);
  and (_06505_, _06503_, _06500_);
  nor (_06506_, _06505_, _06504_);
  and (_06507_, _06506_, _06494_);
  nor (_06508_, _06507_, _06504_);
  nor (_06509_, _06447_, _06445_);
  nor (_06510_, _06509_, _06448_);
  not (_06511_, _06510_);
  nor (_06512_, _06511_, _06508_);
  and (_06513_, _06452_, _06449_);
  nor (_06514_, _06513_, _06453_);
  and (_06515_, _06514_, _06512_);
  nor (_06516_, _06455_, _06453_);
  nor (_06517_, _06516_, _06456_);
  and (_06518_, _06517_, _06515_);
  nor (_06519_, _06517_, _06515_);
  nor (_06520_, _06519_, _06518_);
  and (_06521_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  and (_06522_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and (_06523_, _06522_, _06521_);
  and (_06524_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor (_06525_, _06522_, _06521_);
  nor (_06526_, _06525_, _06523_);
  and (_06527_, _06526_, _06524_);
  nor (_06528_, _06527_, _06523_);
  not (_06529_, _06528_);
  nor (_06530_, _06464_, _06462_);
  nor (_06531_, _06530_, _06465_);
  and (_06532_, _06531_, _06529_);
  and (_06533_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and (_06534_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and (_06535_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [1]);
  and (_06536_, _06535_, _06534_);
  nor (_06537_, _06535_, _06534_);
  nor (_06538_, _06537_, _06536_);
  and (_06539_, _06538_, _06533_);
  nor (_06540_, _06538_, _06533_);
  nor (_06541_, _06540_, _06539_);
  nor (_06542_, _06531_, _06529_);
  nor (_06543_, _06542_, _06532_);
  and (_06544_, _06543_, _06541_);
  nor (_06545_, _06544_, _06532_);
  not (_06546_, _06545_);
  nor (_06547_, _06481_, _06479_);
  nor (_06548_, _06547_, _06482_);
  and (_06549_, _06548_, _06546_);
  not (_06550_, _06424_);
  nor (_06551_, _06539_, _06536_);
  nor (_06552_, _06551_, _06550_);
  and (_06553_, _06551_, _06550_);
  nor (_06554_, _06553_, _06552_);
  nor (_06555_, _06548_, _06546_);
  nor (_06556_, _06555_, _06549_);
  and (_06557_, _06556_, _06554_);
  nor (_06558_, _06557_, _06549_);
  not (_06559_, _06558_);
  nor (_06560_, _06498_, _06496_);
  nor (_06561_, _06560_, _06499_);
  and (_06562_, _06561_, _06559_);
  nor (_06563_, _06561_, _06559_);
  nor (_06564_, _06563_, _06562_);
  and (_06565_, _06564_, _06552_);
  nor (_06566_, _06565_, _06562_);
  nor (_06567_, _06506_, _06494_);
  nor (_06568_, _06567_, _06507_);
  not (_06569_, _06568_);
  nor (_06570_, _06569_, _06566_);
  and (_06571_, _06511_, _06508_);
  nor (_06572_, _06571_, _06512_);
  and (_06573_, _06572_, _06570_);
  nor (_06574_, _06514_, _06512_);
  nor (_06575_, _06574_, _06515_);
  and (_06576_, _06575_, _06573_);
  nor (_06577_, _06575_, _06573_);
  nor (_06578_, _06577_, _06576_);
  and (_06579_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and (_06580_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and (_06581_, _06580_, _06579_);
  and (_06582_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [1]);
  nor (_06583_, _06580_, _06579_);
  nor (_06584_, _06583_, _06581_);
  and (_06585_, _06584_, _06582_);
  nor (_06586_, _06585_, _06581_);
  not (_06587_, _06586_);
  nor (_06588_, _06526_, _06524_);
  nor (_06589_, _06588_, _06527_);
  and (_06590_, _06589_, _06587_);
  and (_06591_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and (_06592_, _06591_, _06535_);
  and (_06593_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [1]);
  and (_06594_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor (_06595_, _06594_, _06593_);
  nor (_06596_, _06595_, _06592_);
  nor (_06597_, _06589_, _06587_);
  nor (_06598_, _06597_, _06590_);
  and (_06599_, _06598_, _06596_);
  nor (_06600_, _06599_, _06590_);
  not (_06601_, _06600_);
  nor (_06602_, _06543_, _06541_);
  nor (_06603_, _06602_, _06544_);
  and (_06604_, _06603_, _06601_);
  nor (_06605_, _06603_, _06601_);
  nor (_06606_, _06605_, _06604_);
  and (_06607_, _06606_, _06592_);
  nor (_06608_, _06607_, _06604_);
  not (_06609_, _06608_);
  nor (_06610_, _06556_, _06554_);
  nor (_06611_, _06610_, _06557_);
  and (_06612_, _06611_, _06609_);
  nor (_06613_, _06564_, _06552_);
  nor (_06614_, _06613_, _06565_);
  and (_06615_, _06614_, _06612_);
  and (_06616_, _06569_, _06566_);
  nor (_06617_, _06616_, _06570_);
  and (_06618_, _06617_, _06615_);
  nor (_06619_, _06572_, _06570_);
  nor (_06620_, _06619_, _06573_);
  nor (_06621_, _06620_, _06618_);
  and (_06622_, _06620_, _06618_);
  not (_06623_, _06622_);
  and (_06624_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and (_06625_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [1]);
  and (_06626_, _06625_, _06624_);
  and (_06627_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor (_06628_, _06625_, _06624_);
  nor (_06629_, _06628_, _06626_);
  and (_06630_, _06629_, _06627_);
  nor (_06631_, _06630_, _06626_);
  not (_06632_, _06631_);
  nor (_06633_, _06584_, _06582_);
  nor (_06634_, _06633_, _06585_);
  and (_06635_, _06634_, _06632_);
  nor (_06636_, _06634_, _06632_);
  nor (_06637_, _06636_, _06635_);
  and (_06638_, _06637_, _06591_);
  nor (_06639_, _06638_, _06635_);
  not (_06640_, _06639_);
  nor (_06641_, _06598_, _06596_);
  nor (_06642_, _06641_, _06599_);
  and (_06643_, _06642_, _06640_);
  nor (_06644_, _06606_, _06592_);
  nor (_06645_, _06644_, _06607_);
  and (_06646_, _06645_, _06643_);
  nor (_06647_, _06611_, _06609_);
  nor (_06648_, _06647_, _06612_);
  and (_06649_, _06648_, _06646_);
  nor (_06650_, _06614_, _06612_);
  nor (_06651_, _06650_, _06615_);
  and (_06652_, _06651_, _06649_);
  nor (_06653_, _06617_, _06615_);
  nor (_06654_, _06653_, _06618_);
  and (_06655_, _06654_, _06652_);
  and (_06656_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  and (_06657_, _06656_, _06625_);
  nor (_06658_, _06629_, _06627_);
  nor (_06659_, _06658_, _06630_);
  and (_06660_, _06659_, _06657_);
  nor (_06661_, _06637_, _06591_);
  nor (_06662_, _06661_, _06638_);
  and (_06663_, _06662_, _06660_);
  nor (_06664_, _06642_, _06640_);
  nor (_06665_, _06664_, _06643_);
  and (_06666_, _06665_, _06663_);
  nor (_06667_, _06645_, _06643_);
  nor (_06668_, _06667_, _06646_);
  and (_06669_, _06668_, _06666_);
  nor (_06670_, _06648_, _06646_);
  nor (_06671_, _06670_, _06649_);
  and (_06672_, _06671_, _06669_);
  nor (_06673_, _06651_, _06649_);
  nor (_06674_, _06673_, _06652_);
  and (_06675_, _06674_, _06672_);
  nor (_06676_, _06654_, _06652_);
  nor (_06677_, _06676_, _06655_);
  and (_06678_, _06677_, _06675_);
  nor (_06679_, _06678_, _06655_);
  and (_06680_, _06679_, _06623_);
  nor (_06681_, _06680_, _06621_);
  and (_06682_, _06681_, _06578_);
  nor (_06683_, _06682_, _06576_);
  not (_06684_, _06683_);
  and (_06685_, _06684_, _06520_);
  nor (_06686_, _06685_, _06518_);
  not (_06687_, _06686_);
  nor (_06688_, _06458_, _06456_);
  nor (_06689_, _06688_, _06459_);
  and (_06690_, _06689_, _06687_);
  nor (_06691_, _06690_, _06459_);
  not (_06692_, _06691_);
  and (_06693_, _06692_, _06394_);
  nor (_06694_, _06693_, _06392_);
  not (_06695_, _06694_);
  and (_06696_, \oc8051_golden_model_1.B [7], \oc8051_golden_model_1.ACC [7]);
  not (_06697_, _06696_);
  nor (_06698_, _06697_, _06344_);
  nor (_06699_, _06698_, _06376_);
  nor (_06700_, _06382_, _06379_);
  nor (_06701_, _06700_, _06699_);
  and (_06702_, _06700_, _06699_);
  nor (_06703_, _06702_, _06701_);
  not (_06704_, _06703_);
  nor (_06705_, _06389_, _06386_);
  and (_06706_, _06705_, _06704_);
  nor (_06707_, _06705_, _06704_);
  nor (_06708_, _06707_, _06706_);
  and (_06709_, _06708_, _06695_);
  or (_06710_, _06701_, _06373_);
  or (_06711_, _06710_, _06707_);
  or (_06712_, _06711_, _06709_);
  or (_06713_, _06712_, _06201_);
  and (_06714_, _06713_, _02966_);
  and (_06715_, _06714_, _06200_);
  not (_06716_, _05286_);
  nor (_06717_, _05502_, _06716_);
  or (_06718_, _06717_, _06179_);
  and (_06719_, _06718_, _02785_);
  or (_06720_, _06719_, _03861_);
  or (_06721_, _06720_, _06715_);
  or (_06722_, _06177_, _03860_);
  and (_06723_, _06722_, _06721_);
  or (_06724_, _06723_, _03850_);
  and (_06725_, _05426_, _04661_);
  not (_06726_, _03850_);
  or (_06727_, _06163_, _06726_);
  or (_06728_, _06727_, _06725_);
  and (_06729_, _06728_, _02970_);
  and (_06730_, _06729_, _06724_);
  and (_06731_, _02978_, _02347_);
  and (_06732_, _05706_, _04661_);
  or (_06733_, _06732_, _06163_);
  and (_06734_, _06733_, _02524_);
  or (_06735_, _06734_, _06731_);
  or (_06736_, _06735_, _06730_);
  not (_06737_, _06731_);
  not (_06738_, \oc8051_golden_model_1.B [1]);
  nor (_06739_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [5]);
  nor (_06740_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.B [3]);
  and (_06741_, _06740_, _06739_);
  and (_06742_, _06741_, _06738_);
  not (_06743_, \oc8051_golden_model_1.B [0]);
  and (_06744_, _06743_, \oc8051_golden_model_1.ACC [7]);
  nor (_06745_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  and (_06746_, _06745_, _06744_);
  and (_06747_, _06746_, _06742_);
  not (_06748_, _06745_);
  and (_06749_, \oc8051_golden_model_1.B [0], _05719_);
  nor (_06750_, _06749_, _06748_);
  and (_06751_, _06750_, _06742_);
  or (_06752_, _06751_, _05719_);
  not (_06753_, \oc8051_golden_model_1.B [2]);
  not (_06754_, \oc8051_golden_model_1.B [3]);
  not (_06755_, \oc8051_golden_model_1.B [4]);
  not (_06756_, \oc8051_golden_model_1.B [5]);
  nor (_06757_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and (_06758_, _06757_, _06756_);
  and (_06759_, _06758_, _06755_);
  and (_06760_, _06759_, _06754_);
  and (_06761_, _06760_, _06753_);
  not (_06762_, \oc8051_golden_model_1.ACC [6]);
  and (_06763_, \oc8051_golden_model_1.B [0], _06762_);
  nor (_06764_, _06763_, _05719_);
  nor (_06765_, _06764_, _06738_);
  not (_06766_, _06765_);
  and (_06767_, _06766_, _06761_);
  nor (_06768_, _06767_, _06752_);
  nor (_06769_, _06768_, _06747_);
  and (_06770_, _06767_, \oc8051_golden_model_1.B [0]);
  nor (_06771_, _06770_, _06762_);
  and (_06772_, _06771_, _06738_);
  nor (_06773_, _06771_, _06738_);
  nor (_06774_, _06773_, _06772_);
  nor (_06775_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [5]);
  nor (_06776_, _06775_, _06395_);
  nor (_06777_, _06776_, \oc8051_golden_model_1.ACC [4]);
  nor (_06778_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  and (_06779_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.ACC [4]);
  nor (_06780_, _06779_, _06743_);
  nor (_06781_, _06780_, _06778_);
  nor (_06782_, _06781_, _06777_);
  not (_06783_, _06782_);
  and (_06784_, _06783_, _06774_);
  nor (_06785_, _06769_, \oc8051_golden_model_1.B [2]);
  nor (_06786_, _06785_, _06772_);
  not (_06787_, _06786_);
  nor (_06788_, _06787_, _06784_);
  and (_06789_, \oc8051_golden_model_1.B [2], _05719_);
  nor (_06790_, _06789_, \oc8051_golden_model_1.B [7]);
  and (_06791_, _06790_, _06741_);
  not (_06792_, _06791_);
  nor (_06793_, _06792_, _06788_);
  nor (_06794_, _06793_, _06769_);
  nor (_06795_, _06794_, _06747_);
  and (_06796_, _06759_, \oc8051_golden_model_1.ACC [7]);
  nor (_06797_, _06796_, _06760_);
  nor (_06798_, _06783_, _06774_);
  nor (_06799_, _06798_, _06784_);
  not (_06800_, _06799_);
  and (_06801_, _06800_, _06793_);
  nor (_06802_, _06793_, _06771_);
  nor (_06803_, _06802_, _06801_);
  and (_06804_, _06803_, _06753_);
  nor (_06805_, _06803_, _06753_);
  nor (_06806_, _06805_, _06804_);
  not (_06807_, _06806_);
  not (_06808_, \oc8051_golden_model_1.ACC [5]);
  nor (_06809_, _06793_, _06808_);
  and (_06810_, _06793_, _06776_);
  or (_06811_, _06810_, _06809_);
  and (_06812_, _06811_, _06738_);
  nor (_06813_, _06811_, _06738_);
  not (_06814_, \oc8051_golden_model_1.ACC [4]);
  and (_06815_, \oc8051_golden_model_1.B [0], _06814_);
  nor (_06816_, _06815_, _06813_);
  nor (_06817_, _06816_, _06812_);
  nor (_06818_, _06817_, _06807_);
  nor (_06819_, _06795_, \oc8051_golden_model_1.B [3]);
  nor (_06820_, _06819_, _06804_);
  not (_06821_, _06820_);
  nor (_06822_, _06821_, _06818_);
  nor (_06823_, _06822_, _06797_);
  nor (_06824_, _06823_, _06795_);
  nor (_06825_, _06824_, _06747_);
  nor (_06826_, _06825_, \oc8051_golden_model_1.B [4]);
  not (_06827_, _06823_);
  and (_06828_, _06817_, _06807_);
  nor (_06829_, _06828_, _06818_);
  nor (_06830_, _06829_, _06827_);
  nor (_06831_, _06823_, _06803_);
  nor (_06832_, _06831_, _06830_);
  and (_06833_, _06832_, _06754_);
  nor (_06834_, _06832_, _06754_);
  nor (_06835_, _06834_, _06833_);
  not (_06836_, _06835_);
  nor (_06837_, _06823_, _06811_);
  nor (_06838_, _06813_, _06812_);
  and (_06839_, _06838_, _06815_);
  nor (_06840_, _06838_, _06815_);
  nor (_06841_, _06840_, _06839_);
  and (_06842_, _06841_, _06823_);
  or (_06843_, _06842_, _06837_);
  nor (_06844_, _06843_, \oc8051_golden_model_1.B [2]);
  and (_06845_, _06843_, \oc8051_golden_model_1.B [2]);
  nor (_06846_, _06823_, _06814_);
  nor (_06847_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [4]);
  nor (_06848_, _06847_, _06521_);
  and (_06849_, _06823_, _06848_);
  or (_06850_, _06849_, _06846_);
  and (_06851_, _06850_, _06738_);
  nor (_06852_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor (_06853_, _06852_, _06579_);
  nor (_06854_, _06853_, \oc8051_golden_model_1.ACC [2]);
  nor (_06855_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  and (_06856_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.ACC [2]);
  nor (_06857_, _06856_, _06743_);
  nor (_06858_, _06857_, _06855_);
  nor (_06859_, _06858_, _06854_);
  not (_06860_, _06859_);
  nor (_06861_, _06850_, _06738_);
  nor (_06862_, _06861_, _06851_);
  and (_06863_, _06862_, _06860_);
  nor (_06864_, _06863_, _06851_);
  nor (_06865_, _06864_, _06845_);
  nor (_06866_, _06865_, _06844_);
  nor (_06867_, _06866_, _06836_);
  or (_06868_, _06867_, _06833_);
  nor (_06869_, _06868_, _06826_);
  and (_06870_, _06758_, \oc8051_golden_model_1.ACC [7]);
  or (_06871_, _06870_, _06759_);
  not (_06872_, _06871_);
  nor (_06873_, _06872_, _06869_);
  nor (_06874_, _06873_, _06825_);
  nor (_06875_, _06874_, _06747_);
  and (_06876_, _06866_, _06836_);
  nor (_06877_, _06876_, _06867_);
  not (_06878_, _06877_);
  and (_06879_, _06878_, _06873_);
  nor (_06880_, _06873_, _06832_);
  nor (_06881_, _06880_, _06879_);
  and (_06882_, _06881_, _06755_);
  nor (_06883_, _06881_, _06755_);
  nor (_06884_, _06883_, _06882_);
  not (_06885_, _06884_);
  nor (_06886_, _06873_, _06843_);
  nor (_06887_, _06845_, _06844_);
  and (_06888_, _06887_, _06864_);
  nor (_06889_, _06887_, _06864_);
  nor (_06890_, _06889_, _06888_);
  not (_06891_, _06890_);
  and (_06892_, _06891_, _06873_);
  nor (_06893_, _06892_, _06886_);
  nor (_06894_, _06893_, \oc8051_golden_model_1.B [3]);
  and (_06895_, _06893_, \oc8051_golden_model_1.B [3]);
  nor (_06896_, _06862_, _06860_);
  nor (_06897_, _06896_, _06863_);
  not (_06898_, _06897_);
  and (_06899_, _06898_, _06873_);
  nor (_06900_, _06873_, _06850_);
  nor (_06901_, _06900_, _06899_);
  and (_06902_, _06901_, _06753_);
  nor (_06903_, _06873_, _02605_);
  and (_06904_, _06873_, _06853_);
  or (_06905_, _06904_, _06903_);
  and (_06906_, _06905_, _06738_);
  nor (_06907_, _06905_, _06738_);
  not (_06908_, \oc8051_golden_model_1.ACC [2]);
  and (_06909_, \oc8051_golden_model_1.B [0], _06908_);
  nor (_06910_, _06909_, _06907_);
  nor (_06911_, _06910_, _06906_);
  nor (_06912_, _06901_, _06753_);
  nor (_06913_, _06912_, _06902_);
  not (_06914_, _06913_);
  nor (_06915_, _06914_, _06911_);
  nor (_06916_, _06915_, _06902_);
  nor (_06917_, _06916_, _06895_);
  nor (_06918_, _06917_, _06894_);
  nor (_06919_, _06918_, _06885_);
  nor (_06920_, _06875_, \oc8051_golden_model_1.B [5]);
  nor (_06921_, _06920_, _06882_);
  not (_06922_, _06921_);
  nor (_06923_, _06922_, _06919_);
  not (_06924_, _06923_);
  not (_06925_, _06757_);
  and (_06926_, \oc8051_golden_model_1.B [5], _05719_);
  nor (_06927_, _06926_, _06925_);
  and (_06928_, _06927_, _06924_);
  nor (_06929_, _06928_, _06875_);
  nor (_06930_, _06929_, _06747_);
  nor (_06931_, _06930_, \oc8051_golden_model_1.B [6]);
  and (_06932_, \oc8051_golden_model_1.B [6], _05719_);
  not (_06933_, _06928_);
  and (_06934_, _06918_, _06885_);
  nor (_06935_, _06934_, _06919_);
  nor (_06936_, _06935_, _06933_);
  nor (_06937_, _06928_, _06881_);
  nor (_06938_, _06937_, _06936_);
  and (_06939_, _06938_, _06756_);
  nor (_06940_, _06938_, _06756_);
  nor (_06941_, _06940_, _06939_);
  not (_06942_, _06941_);
  nor (_06943_, _06895_, _06894_);
  nor (_06944_, _06943_, _06916_);
  and (_06945_, _06943_, _06916_);
  or (_06946_, _06945_, _06944_);
  nor (_06947_, _06946_, _06933_);
  and (_06948_, _06933_, _06893_);
  nor (_06949_, _06948_, _06947_);
  and (_06950_, _06949_, _06755_);
  nor (_06951_, _06949_, _06755_);
  and (_06952_, _06914_, _06911_);
  nor (_06953_, _06952_, _06915_);
  nor (_06954_, _06953_, _06933_);
  nor (_06955_, _06928_, _06901_);
  nor (_06956_, _06955_, _06954_);
  and (_06957_, _06956_, _06754_);
  nor (_06958_, _06907_, _06906_);
  nor (_06959_, _06958_, _06909_);
  and (_06960_, _06958_, _06909_);
  or (_06961_, _06960_, _06959_);
  nor (_06962_, _06961_, _06933_);
  nor (_06963_, _06928_, _06905_);
  nor (_06964_, _06963_, _06962_);
  and (_06965_, _06964_, _06753_);
  nor (_06966_, _06964_, _06753_);
  nor (_06967_, _06928_, \oc8051_golden_model_1.ACC [2]);
  nor (_06968_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  nor (_06969_, _06968_, _06624_);
  nor (_06970_, _06933_, _06969_);
  nor (_06971_, _06970_, _06967_);
  and (_06972_, _06971_, _06738_);
  and (_06973_, \oc8051_golden_model_1.B [0], _02477_);
  not (_06974_, _06973_);
  nor (_06975_, _06971_, _06738_);
  nor (_06976_, _06975_, _06972_);
  and (_06977_, _06976_, _06974_);
  nor (_06978_, _06977_, _06972_);
  nor (_06979_, _06978_, _06966_);
  nor (_06980_, _06979_, _06965_);
  nor (_06981_, _06956_, _06754_);
  nor (_06982_, _06981_, _06957_);
  not (_06983_, _06982_);
  nor (_06984_, _06983_, _06980_);
  nor (_06985_, _06984_, _06957_);
  nor (_06986_, _06985_, _06951_);
  nor (_06987_, _06986_, _06950_);
  nor (_06988_, _06987_, _06942_);
  nor (_06989_, _06988_, _06939_);
  nor (_06990_, _06989_, _06932_);
  nor (_06991_, _06990_, _06931_);
  nor (_06992_, _06991_, \oc8051_golden_model_1.B [7]);
  nor (_06993_, _06992_, _06930_);
  or (_06994_, _06993_, _06747_);
  nor (_06995_, _06994_, \oc8051_golden_model_1.B [7]);
  nor (_06996_, _06995_, _06696_);
  not (_06997_, \oc8051_golden_model_1.B [6]);
  and (_06998_, _06987_, _06942_);
  nor (_06999_, _06998_, _06988_);
  not (_07000_, _06999_);
  and (_07001_, _07000_, _06992_);
  nor (_07002_, _06992_, _06938_);
  nor (_07003_, _07002_, _07001_);
  nor (_07004_, _07003_, _06997_);
  not (_07005_, _07004_);
  nor (_07006_, _07005_, _06996_);
  nor (_07007_, _06966_, _06965_);
  and (_07008_, _07007_, _06978_);
  nor (_07009_, _07007_, _06978_);
  or (_07010_, _07009_, _07008_);
  and (_07011_, _07010_, _06992_);
  not (_07012_, _06964_);
  nor (_07013_, _06992_, _07012_);
  nor (_07014_, _07013_, _07011_);
  nor (_07015_, _07014_, \oc8051_golden_model_1.B [3]);
  and (_07016_, _07014_, \oc8051_golden_model_1.B [3]);
  nor (_07017_, _07016_, _07015_);
  nor (_07018_, _06976_, _06974_);
  nor (_07019_, _07018_, _06977_);
  and (_07020_, _07019_, _06992_);
  not (_07021_, _06971_);
  nor (_07022_, _06992_, _07021_);
  nor (_07023_, _07022_, _07020_);
  and (_07024_, _07023_, \oc8051_golden_model_1.B [2]);
  nor (_07025_, _07023_, \oc8051_golden_model_1.B [2]);
  nor (_07026_, _07025_, _07024_);
  and (_07027_, _07026_, _07017_);
  nor (_07028_, _06992_, \oc8051_golden_model_1.ACC [1]);
  and (_07029_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  nor (_07030_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [1]);
  or (_07031_, _07030_, _07029_);
  and (_07032_, _06992_, _07031_);
  nor (_07033_, _07032_, _07028_);
  and (_07034_, _07033_, _06738_);
  nor (_07035_, _07033_, _06738_);
  and (_07036_, _06743_, \oc8051_golden_model_1.ACC [0]);
  not (_07037_, _07036_);
  nor (_07038_, _07037_, _07035_);
  nor (_07039_, _07038_, _07034_);
  and (_07040_, _07039_, _07027_);
  not (_07041_, _07040_);
  and (_07042_, _07024_, _07017_);
  nor (_07043_, _07042_, _07016_);
  and (_07044_, _07043_, _07041_);
  and (_07045_, _06983_, _06980_);
  or (_07046_, _07045_, _06984_);
  and (_07047_, _07046_, _06992_);
  nor (_07048_, _06992_, _06956_);
  nor (_07049_, _07048_, _07047_);
  nor (_07050_, _07049_, _06755_);
  and (_07051_, _07049_, _06755_);
  nor (_07052_, _07051_, _07050_);
  nor (_07053_, _06951_, _06950_);
  nor (_07054_, _07053_, _06985_);
  and (_07055_, _07053_, _06985_);
  nor (_07056_, _07055_, _07054_);
  and (_07057_, _07056_, _06992_);
  nor (_07058_, _06992_, _06949_);
  or (_07059_, _07058_, _07057_);
  and (_07060_, _07059_, \oc8051_golden_model_1.B [5]);
  nor (_07061_, _07059_, \oc8051_golden_model_1.B [5]);
  nor (_07062_, _07061_, _07060_);
  and (_07063_, _07062_, _07052_);
  and (_07064_, _07003_, _06997_);
  nor (_07065_, _07064_, _07004_);
  not (_07066_, _07065_);
  nor (_07067_, _07066_, _06996_);
  and (_07068_, _07067_, _07063_);
  not (_07069_, _07068_);
  nor (_07070_, _07069_, _07044_);
  and (_07071_, _06930_, \oc8051_golden_model_1.B [7]);
  and (_07072_, _07062_, _07050_);
  nor (_07073_, _07072_, _07060_);
  not (_07074_, _07073_);
  and (_07075_, _07074_, _07067_);
  or (_07076_, _07075_, _07071_);
  or (_07077_, _07076_, _07070_);
  nor (_07078_, _07077_, _07006_);
  and (_07079_, \oc8051_golden_model_1.B [0], _02658_);
  not (_07080_, _07079_);
  nor (_07081_, _07035_, _07034_);
  and (_07082_, _07081_, _07080_);
  and (_07083_, _07082_, _07037_);
  and (_07084_, _07083_, _07027_);
  and (_07085_, _07084_, _07068_);
  nor (_07086_, _07085_, _07078_);
  or (_07087_, _07086_, _06747_);
  and (_07088_, _07087_, _06994_);
  or (_07089_, _07088_, _06737_);
  and (_07090_, _07089_, _06736_);
  or (_07091_, _07090_, _02974_);
  not (_07092_, _02977_);
  and (_07093_, _05517_, _04661_);
  or (_07094_, _07093_, _06163_);
  or (_07095_, _07094_, _05261_);
  and (_07096_, _07095_, _07092_);
  and (_07097_, _07096_, _07091_);
  and (_07098_, _05259_, _04661_);
  or (_07099_, _06163_, _03107_);
  nor (_07100_, _07099_, _07098_);
  nor (_07101_, _07100_, _03108_);
  or (_07102_, _07101_, _07097_);
  and (_07103_, _05722_, _04661_);
  not (_07104_, _03107_);
  or (_07105_, _06163_, _07104_);
  or (_07106_, _07105_, _07103_);
  and (_07107_, _07106_, _03881_);
  and (_07108_, _07107_, _07102_);
  or (_07109_, _06163_, _04690_);
  and (_07110_, _07094_, _02991_);
  and (_07111_, _07110_, _07109_);
  or (_07112_, _07111_, _07108_);
  and (_07113_, _07112_, _06161_);
  and (_07114_, _06168_, _03094_);
  and (_07115_, _07114_, _07109_);
  or (_07116_, _07115_, _02994_);
  or (_07117_, _07116_, _07113_);
  not (_07118_, _03099_);
  nor (_07119_, _05257_, _06175_);
  not (_07120_, _02994_);
  or (_07121_, _06163_, _07120_);
  or (_07122_, _07121_, _07119_);
  and (_07123_, _07122_, _07118_);
  and (_07124_, _07123_, _07117_);
  nor (_07125_, _05721_, _06175_);
  or (_07126_, _07125_, _06163_);
  and (_07127_, _07126_, _03099_);
  or (_07128_, _07127_, _03133_);
  or (_07129_, _07128_, _07124_);
  or (_07130_, _06165_, _03138_);
  and (_07131_, _07130_, _03142_);
  and (_07132_, _07131_, _07129_);
  and (_07133_, _06191_, _02778_);
  or (_07134_, _07133_, _02852_);
  or (_07135_, _07134_, _07132_);
  and (_07136_, _05196_, _04661_);
  or (_07137_, _06163_, _02853_);
  or (_07138_, _07137_, _07136_);
  and (_07139_, _07138_, _34446_);
  and (_07140_, _07139_, _07135_);
  or (_07141_, _07140_, _06160_);
  and (_35615_[7], _07141_, _35583_);
  nor (_07142_, _34446_, _05719_);
  and (_07143_, _02574_, _02475_);
  nand (_07144_, _07143_, _06762_);
  nor (_07145_, _05426_, \oc8051_golden_model_1.ACC [7]);
  and (_07146_, _05426_, \oc8051_golden_model_1.ACC [7]);
  nor (_07147_, _07146_, _07145_);
  and (_07148_, _05798_, \oc8051_golden_model_1.ACC [6]);
  nor (_07149_, _05798_, \oc8051_golden_model_1.ACC [6]);
  nor (_07150_, _07149_, _07148_);
  and (_07151_, _06120_, \oc8051_golden_model_1.ACC [5]);
  and (_07152_, _06027_, _06808_);
  nor (_07153_, _07152_, _07151_);
  not (_07154_, _07153_);
  and (_07155_, _06121_, \oc8051_golden_model_1.ACC [4]);
  and (_07156_, _06072_, _06814_);
  nor (_07157_, _07156_, _07155_);
  and (_07158_, _06116_, \oc8051_golden_model_1.ACC [3]);
  and (_07159_, _05935_, _02605_);
  and (_07160_, _06117_, \oc8051_golden_model_1.ACC [2]);
  and (_07161_, _05980_, _06908_);
  nor (_07162_, _07161_, _07160_);
  not (_07163_, _07162_);
  and (_07164_, _06113_, \oc8051_golden_model_1.ACC [1]);
  and (_07165_, _05844_, _02477_);
  nor (_07166_, _07165_, _07164_);
  and (_07167_, _06114_, \oc8051_golden_model_1.ACC [0]);
  and (_07168_, _07167_, _07166_);
  nor (_07169_, _07168_, _07164_);
  nor (_07170_, _07169_, _07163_);
  nor (_07171_, _07170_, _07160_);
  nor (_07172_, _07171_, _07159_);
  or (_07173_, _07172_, _07158_);
  and (_07174_, _07173_, _07157_);
  nor (_07175_, _07174_, _07155_);
  nor (_07176_, _07175_, _07154_);
  or (_07177_, _07176_, _07151_);
  and (_07178_, _07177_, _07150_);
  nor (_07179_, _07178_, _07148_);
  nor (_07180_, _07179_, _07147_);
  and (_07181_, _07179_, _07147_);
  nor (_07182_, _07181_, _07180_);
  and (_07183_, _02971_, _02574_);
  nand (_07184_, _07183_, _07182_);
  and (_07185_, _02999_, _02574_);
  or (_07186_, _07185_, _03260_);
  not (_07187_, _07186_);
  and (_07188_, _02907_, _02574_);
  nor (_07189_, _03702_, _07188_);
  and (_07190_, _07189_, _07187_);
  and (_07191_, _03857_, _02574_);
  not (_07192_, _07191_);
  and (_07193_, _07192_, _07190_);
  and (_07194_, _04585_, _05719_);
  nor (_07195_, _04585_, _05719_);
  nor (_07196_, _07195_, _07194_);
  nor (_07197_, _04735_, _06762_);
  and (_07198_, _04735_, _06762_);
  nor (_07199_, _07198_, _07197_);
  nor (_07200_, _04839_, _06808_);
  and (_07201_, _04839_, _06808_);
  nor (_07202_, _07201_, _07200_);
  not (_07203_, _07202_);
  nor (_07204_, _05143_, _06814_);
  and (_07205_, _05143_, _06814_);
  nor (_07206_, _07205_, _07204_);
  not (_07207_, _07206_);
  nor (_07208_, _04226_, _02605_);
  not (_07209_, _07208_);
  and (_07210_, _04226_, _02605_);
  nor (_07211_, _04413_, _06908_);
  and (_07212_, _04413_, _06908_);
  nor (_07213_, _07212_, _07211_);
  not (_07214_, _07213_);
  nor (_07215_, _03989_, _02477_);
  and (_07216_, _03989_, _02477_);
  nor (_07217_, _07216_, _07215_);
  and (_07218_, _03805_, \oc8051_golden_model_1.ACC [0]);
  and (_07219_, _07218_, _07217_);
  nor (_07220_, _07219_, _07215_);
  nor (_07221_, _07220_, _07214_);
  nor (_07222_, _07221_, _07211_);
  or (_07223_, _07222_, _07210_);
  and (_07224_, _07223_, _07209_);
  nor (_07225_, _07224_, _07207_);
  nor (_07226_, _07225_, _07204_);
  nor (_07227_, _07226_, _07203_);
  or (_07228_, _07227_, _07200_);
  and (_07229_, _07228_, _07199_);
  nor (_07230_, _07229_, _07197_);
  nor (_07231_, _07230_, _07196_);
  and (_07232_, _07230_, _07196_);
  nor (_07233_, _07232_, _07231_);
  nor (_07234_, _07233_, _03542_);
  or (_07235_, _07234_, _07193_);
  and (_07236_, _02971_, _02591_);
  not (_07237_, _02591_);
  nor (_07238_, _03011_, _02906_);
  nor (_07239_, _07238_, _07237_);
  and (_07240_, _03857_, _02591_);
  nor (_07241_, _07240_, _07239_);
  not (_07242_, _04735_);
  and (_07243_, _05205_, \oc8051_golden_model_1.PSW [7]);
  and (_07244_, _07243_, _07242_);
  nor (_07245_, _07244_, _04585_);
  and (_07246_, _07244_, _04585_);
  nor (_07247_, _07246_, _07245_);
  and (_07248_, _07247_, \oc8051_golden_model_1.ACC [7]);
  nor (_07249_, _07247_, \oc8051_golden_model_1.ACC [7]);
  nor (_07250_, _07249_, _07248_);
  nor (_07251_, _07243_, _07242_);
  nor (_07252_, _07251_, _07244_);
  and (_07253_, _07252_, \oc8051_golden_model_1.ACC [6]);
  and (_07254_, _07252_, _06762_);
  nor (_07255_, _07252_, _06762_);
  nor (_07256_, _07255_, _07254_);
  and (_07257_, _05204_, \oc8051_golden_model_1.PSW [7]);
  nor (_07258_, _07257_, _05199_);
  nor (_07259_, _07258_, _07243_);
  and (_07260_, _07259_, \oc8051_golden_model_1.ACC [5]);
  and (_07261_, _07259_, _06808_);
  nor (_07262_, _07259_, _06808_);
  nor (_07263_, _07262_, _07261_);
  and (_07264_, _05201_, \oc8051_golden_model_1.PSW [7]);
  and (_07265_, _07264_, _05202_);
  nor (_07266_, _07265_, _05200_);
  nor (_07267_, _07266_, _07257_);
  and (_07268_, _07267_, \oc8051_golden_model_1.ACC [4]);
  nor (_07269_, _07267_, _06814_);
  and (_07270_, _07267_, _06814_);
  nor (_07271_, _07270_, _07269_);
  not (_07272_, _04226_);
  and (_07273_, _05201_, _04414_);
  and (_07274_, _07273_, \oc8051_golden_model_1.PSW [7]);
  nor (_07275_, _07274_, _07272_);
  nor (_07276_, _07275_, _07265_);
  and (_07277_, _07276_, \oc8051_golden_model_1.ACC [3]);
  nor (_07278_, _07276_, _02605_);
  and (_07279_, _07276_, _02605_);
  nor (_07280_, _07279_, _07278_);
  nor (_07281_, _07264_, _04414_);
  nor (_07282_, _07281_, _07274_);
  and (_07283_, _07282_, \oc8051_golden_model_1.ACC [2]);
  nor (_07284_, _07282_, _06908_);
  and (_07285_, _07282_, _06908_);
  nor (_07286_, _07285_, _07284_);
  and (_07287_, _03805_, \oc8051_golden_model_1.PSW [7]);
  nor (_07288_, _07287_, _03990_);
  nor (_07289_, _07288_, _07264_);
  and (_07290_, _07289_, \oc8051_golden_model_1.ACC [1]);
  and (_07291_, _07289_, _02477_);
  nor (_07292_, _07289_, _02477_);
  nor (_07293_, _07292_, _07291_);
  not (_07294_, \oc8051_golden_model_1.PSW [7]);
  and (_07295_, _03823_, _07294_);
  nor (_07296_, _07295_, _07287_);
  and (_07297_, _07296_, \oc8051_golden_model_1.ACC [0]);
  not (_07298_, _07297_);
  nor (_07299_, _07298_, _07293_);
  nor (_07300_, _07299_, _07290_);
  nor (_07301_, _07300_, _07286_);
  nor (_07302_, _07301_, _07283_);
  nor (_07303_, _07302_, _07280_);
  nor (_07304_, _07303_, _07277_);
  nor (_07305_, _07304_, _07271_);
  nor (_07306_, _07305_, _07268_);
  nor (_07307_, _07306_, _07263_);
  nor (_07308_, _07307_, _07260_);
  nor (_07309_, _07308_, _07256_);
  nor (_07310_, _07309_, _07253_);
  nor (_07311_, _07310_, _07250_);
  and (_07312_, _07310_, _07250_);
  nor (_07313_, _07312_, _07311_);
  or (_07314_, _07313_, _07241_);
  and (_07315_, _02971_, _02588_);
  nand (_07316_, _02588_, _02409_);
  not (_07317_, _07316_);
  nand (_07318_, _07317_, _07194_);
  and (_07319_, _02978_, _02581_);
  nor (_07320_, _04654_, _05719_);
  and (_07321_, _05426_, _04654_);
  nor (_07322_, _07321_, _07320_);
  nand (_07323_, _07322_, _03850_);
  and (_07324_, _07323_, _02970_);
  not (_07325_, _04654_);
  nor (_07326_, _07325_, _04585_);
  nor (_07327_, _07326_, _07320_);
  nand (_07328_, _07327_, _03861_);
  and (_07329_, _02971_, _02782_);
  not (_07330_, _07329_);
  not (_07331_, _05426_);
  and (_07332_, _06124_, \oc8051_golden_model_1.PSW [7]);
  and (_07333_, _07332_, _07331_);
  nor (_07334_, _07332_, _07331_);
  or (_07335_, _07334_, _07333_);
  nor (_07336_, _07335_, _05719_);
  and (_07337_, _07335_, _05719_);
  nor (_07338_, _07337_, _07336_);
  not (_07339_, _07338_);
  and (_07340_, _06123_, \oc8051_golden_model_1.PSW [7]);
  nor (_07341_, _07340_, _05798_);
  nor (_07342_, _07341_, _07332_);
  nor (_07343_, _07342_, _06762_);
  and (_07344_, _07342_, _06762_);
  and (_07345_, _06119_, _06121_);
  and (_07346_, _07345_, \oc8051_golden_model_1.PSW [7]);
  nor (_07347_, _07346_, _06120_);
  nor (_07348_, _07347_, _07340_);
  and (_07349_, _07348_, _06808_);
  nor (_07350_, _07348_, _06808_);
  and (_07351_, _06115_, \oc8051_golden_model_1.PSW [7]);
  and (_07352_, _07351_, _06118_);
  nor (_07353_, _07352_, _06121_);
  nor (_07354_, _07353_, _07346_);
  nor (_07355_, _07354_, _06814_);
  nor (_07356_, _07355_, _07350_);
  nor (_07357_, _07356_, _07349_);
  nor (_07358_, _07350_, _07349_);
  and (_07359_, _07354_, _06814_);
  nor (_07360_, _07359_, _07355_);
  and (_07361_, _07360_, _07358_);
  and (_07362_, _06115_, _06117_);
  and (_07363_, _07362_, \oc8051_golden_model_1.PSW [7]);
  nor (_07364_, _07363_, _06116_);
  nor (_07365_, _07364_, _07352_);
  nor (_07366_, _07365_, _02605_);
  and (_07367_, _07365_, _02605_);
  nor (_07368_, _07367_, _07366_);
  nor (_07369_, _07351_, _06117_);
  nor (_07370_, _07369_, _07363_);
  nor (_07371_, _07370_, _06908_);
  and (_07372_, _07370_, _06908_);
  nor (_07373_, _07372_, _07371_);
  and (_07374_, _07373_, _07368_);
  and (_07375_, _06114_, \oc8051_golden_model_1.PSW [7]);
  nor (_07376_, _07375_, _06113_);
  nor (_07377_, _07376_, _07351_);
  nor (_07378_, _07377_, _02477_);
  and (_07379_, _07377_, _02477_);
  and (_07380_, _05889_, _07294_);
  nor (_07381_, _07380_, _07375_);
  and (_07382_, _07381_, _02658_);
  nor (_07383_, _07382_, _07379_);
  or (_07384_, _07383_, _07378_);
  and (_07385_, _07384_, _07374_);
  and (_07386_, _07371_, _07368_);
  or (_07387_, _07386_, _07366_);
  nor (_07388_, _07387_, _07385_);
  not (_07389_, _07388_);
  and (_07390_, _07389_, _07361_);
  nor (_07391_, _07390_, _07357_);
  nor (_07392_, _07391_, _07344_);
  or (_07393_, _07392_, _07343_);
  and (_07394_, _07393_, _07339_);
  nor (_07395_, _07393_, _07339_);
  nor (_07396_, _07395_, _07394_);
  nor (_07397_, _07396_, _07330_);
  and (_07398_, _03857_, _02782_);
  nor (_07399_, _07238_, _02498_);
  nor (_07400_, _07399_, _07398_);
  not (_07401_, _07400_);
  and (_07402_, _02978_, _02798_);
  and (_07403_, _05439_, _04654_);
  nor (_07404_, _07403_, _07320_);
  nand (_07405_, _07404_, _02932_);
  not (_07406_, _02934_);
  nor (_07407_, _05466_, _07406_);
  not (_07408_, _03343_);
  or (_07409_, _05426_, _07408_);
  and (_07410_, _03857_, _02933_);
  not (_07411_, _07410_);
  nor (_07412_, _03703_, _03344_);
  and (_07413_, _07412_, _07411_);
  nor (_07414_, _07413_, _04585_);
  and (_07415_, _02978_, _02803_);
  or (_07416_, _07415_, \oc8051_golden_model_1.ACC [7]);
  nand (_07417_, _07415_, \oc8051_golden_model_1.ACC [7]);
  and (_07418_, _07417_, _07416_);
  and (_07419_, _07418_, _07413_);
  or (_07420_, _07419_, _03343_);
  or (_07421_, _07420_, _07414_);
  and (_07422_, _07421_, _07406_);
  and (_07423_, _07422_, _07409_);
  or (_07424_, _07423_, _07407_);
  and (_07425_, _02777_, _02933_);
  nor (_07426_, _02978_, _02475_);
  nor (_07427_, _07426_, _02543_);
  or (_07428_, _07427_, _03363_);
  nor (_07429_, _07428_, _07425_);
  and (_07430_, _07429_, _07424_);
  and (_07431_, _02515_, _02563_);
  and (_07432_, _07431_, _02933_);
  nor (_07433_, _07432_, _07425_);
  not (_07434_, _07433_);
  and (_07435_, _07434_, \oc8051_golden_model_1.XRAM_DATA_IN [7]);
  or (_07436_, _07435_, _02932_);
  or (_07437_, _07436_, _07430_);
  and (_07438_, _07437_, _07405_);
  or (_07439_, _07438_, _07402_);
  nor (_07440_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_07441_, _07440_, _02605_);
  and (_07442_, _07441_, _06779_);
  and (_07443_, _07442_, \oc8051_golden_model_1.ACC [6]);
  and (_07444_, _07443_, \oc8051_golden_model_1.ACC [7]);
  nor (_07445_, _07443_, \oc8051_golden_model_1.ACC [7]);
  nor (_07446_, _07445_, _07444_);
  and (_07447_, _07441_, \oc8051_golden_model_1.ACC [4]);
  nor (_07448_, _07447_, \oc8051_golden_model_1.ACC [5]);
  nor (_07449_, _07448_, _07442_);
  nor (_07450_, _07442_, \oc8051_golden_model_1.ACC [6]);
  nor (_07451_, _07450_, _07443_);
  nor (_07452_, _07451_, _07449_);
  not (_07453_, _07452_);
  and (_07454_, _07453_, _07446_);
  nor (_07455_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_07456_, _07455_, _07452_);
  nor (_07457_, _07456_, _07446_);
  nor (_07458_, _07457_, _07454_);
  not (_07459_, _07458_);
  nand (_07460_, _07459_, _07402_);
  and (_07461_, _07460_, _02939_);
  and (_07462_, _07461_, _07439_);
  nor (_07463_, _05291_, _05719_);
  and (_07464_, _05444_, _05291_);
  nor (_07465_, _07464_, _07463_);
  nor (_07466_, _07465_, _03186_);
  nor (_07467_, _07327_, _03693_);
  and (_07468_, _02919_, _02794_);
  nor (_07469_, _07468_, _03274_);
  not (_07470_, _03241_);
  and (_07471_, _03680_, _02794_);
  and (_07472_, _03008_, _02794_);
  nor (_07473_, _07472_, _07471_);
  and (_07474_, _07473_, _07470_);
  and (_07475_, _07474_, _07469_);
  not (_07476_, _07475_);
  or (_07477_, _07476_, _07467_);
  or (_07478_, _07477_, _07466_);
  or (_07479_, _07478_, _07462_);
  nand (_07480_, _07476_, _04585_);
  and (_07481_, _07480_, _07479_);
  or (_07482_, _07481_, _03374_);
  or (_07483_, _05426_, _03375_);
  and (_07484_, _07483_, _02943_);
  and (_07485_, _07484_, _07482_);
  and (_07486_, _02978_, _02794_);
  nor (_07487_, _05466_, _02943_);
  or (_07488_, _07487_, _07486_);
  or (_07489_, _07488_, _07485_);
  nand (_07490_, _07486_, _02605_);
  and (_07491_, _07490_, _07489_);
  or (_07492_, _07491_, _02796_);
  and (_07493_, _05308_, _05291_);
  nor (_07494_, _07493_, _07463_);
  nand (_07495_, _07494_, _02796_);
  and (_07496_, _07495_, _06189_);
  and (_07497_, _07496_, _07492_);
  and (_07498_, _07464_, _05471_);
  nor (_07499_, _07498_, _07463_);
  nor (_07500_, _07499_, _06189_);
  or (_07501_, _07500_, _06195_);
  or (_07502_, _07501_, _07497_);
  nor (_07503_, _06674_, _06672_);
  nor (_07504_, _07503_, _06675_);
  or (_07505_, _07504_, _06201_);
  and (_07506_, _07505_, _07502_);
  or (_07507_, _07506_, _07401_);
  not (_07508_, _07250_);
  nor (_07509_, _07269_, _07262_);
  nor (_07510_, _07509_, _07261_);
  and (_07511_, _07271_, _07263_);
  not (_07512_, _07511_);
  and (_07513_, _07286_, _07280_);
  nor (_07514_, _07296_, _02658_);
  nor (_07515_, _07514_, _07292_);
  nor (_07516_, _07515_, _07291_);
  not (_07517_, _07516_);
  and (_07518_, _07517_, _07513_);
  not (_07519_, _07518_);
  and (_07520_, _07285_, _07280_);
  nor (_07521_, _07520_, _07279_);
  and (_07522_, _07521_, _07519_);
  and (_07523_, _07296_, _02658_);
  nor (_07524_, _07514_, _07523_);
  and (_07525_, _07524_, _07293_);
  and (_07526_, _07525_, _07513_);
  nor (_07527_, _07526_, _07522_);
  nor (_07528_, _07527_, _07512_);
  nor (_07529_, _07528_, _07510_);
  nor (_07530_, _07529_, _07254_);
  or (_07531_, _07530_, _07255_);
  and (_07532_, _07531_, _07508_);
  nor (_07533_, _07531_, _07508_);
  or (_07534_, _07533_, _07532_);
  or (_07535_, _07534_, _07400_);
  and (_07536_, _07535_, _07330_);
  and (_07537_, _07536_, _07507_);
  or (_07538_, _07537_, _02898_);
  or (_07539_, _07538_, _07397_);
  and (_07540_, _02978_, _02782_);
  not (_07541_, _07540_);
  and (_07542_, _05466_, _05719_);
  nor (_07543_, _05466_, _05719_);
  nor (_07544_, _07543_, _07542_);
  not (_07545_, _07544_);
  and (_07546_, _04679_, \oc8051_golden_model_1.P2INREG [6]);
  and (_07547_, _04681_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_07548_, _07547_, _07546_);
  and (_07549_, _04673_, \oc8051_golden_model_1.P0INREG [6]);
  and (_07550_, _04676_, \oc8051_golden_model_1.P1INREG [6]);
  nor (_07551_, _07550_, _07549_);
  and (_07552_, _07551_, _07548_);
  and (_07553_, _07552_, _04770_);
  and (_07554_, _07553_, _04767_);
  and (_07555_, _07554_, _04754_);
  and (_07556_, _07555_, _04736_);
  and (_07557_, _07556_, \oc8051_golden_model_1.ACC [6]);
  nor (_07558_, _07556_, \oc8051_golden_model_1.ACC [6]);
  nor (_07559_, _07558_, _07557_);
  and (_07560_, _04673_, \oc8051_golden_model_1.P0INREG [5]);
  not (_07561_, _07560_);
  and (_07562_, _04676_, \oc8051_golden_model_1.P1INREG [5]);
  not (_07563_, _07562_);
  and (_07564_, _04679_, \oc8051_golden_model_1.P2INREG [5]);
  and (_07565_, _04681_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_07566_, _07565_, _07564_);
  and (_07567_, _07566_, _07563_);
  and (_07568_, _07567_, _07561_);
  and (_07569_, _07568_, _04876_);
  and (_07570_, _07569_, _04870_);
  and (_07571_, _07570_, _04854_);
  and (_07572_, _07571_, _04840_);
  and (_07573_, _07572_, \oc8051_golden_model_1.ACC [5]);
  nor (_07574_, _07572_, \oc8051_golden_model_1.ACC [5]);
  not (_07575_, _05149_);
  and (_07576_, _05160_, _07575_);
  nor (_07577_, _05152_, _05148_);
  and (_07578_, _07577_, _07576_);
  and (_07579_, _04679_, \oc8051_golden_model_1.P2INREG [4]);
  and (_07580_, _04681_, \oc8051_golden_model_1.P3INREG [4]);
  nor (_07581_, _07580_, _07579_);
  and (_07582_, _04673_, \oc8051_golden_model_1.P0INREG [4]);
  and (_07583_, _04676_, \oc8051_golden_model_1.P1INREG [4]);
  nor (_07584_, _07583_, _07582_);
  and (_07585_, _07584_, _07581_);
  and (_07586_, _07585_, _07578_);
  and (_07587_, _05157_, _05172_);
  not (_07588_, _05184_);
  and (_07589_, _07588_, _05147_);
  and (_07590_, _07589_, _05180_);
  and (_07591_, _07590_, _07587_);
  and (_07592_, _07591_, _07586_);
  and (_07593_, _07592_, _05144_);
  and (_07594_, _07593_, \oc8051_golden_model_1.ACC [4]);
  not (_07595_, _04910_);
  and (_07596_, _04924_, _07595_);
  nor (_07597_, _04916_, _04909_);
  and (_07598_, _07597_, _07596_);
  and (_07599_, _04679_, \oc8051_golden_model_1.P2INREG [3]);
  and (_07600_, _04681_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_07601_, _07600_, _07599_);
  and (_07602_, _04676_, \oc8051_golden_model_1.P1INREG [3]);
  and (_07603_, _04673_, \oc8051_golden_model_1.P0INREG [3]);
  nor (_07604_, _07603_, _07602_);
  and (_07605_, _07604_, _07601_);
  and (_07606_, _07605_, _07598_);
  and (_07607_, _04921_, _04897_);
  and (_07608_, _04935_, _04908_);
  and (_07609_, _07608_, _07607_);
  and (_07610_, _07609_, _07606_);
  and (_07611_, _07610_, _04891_);
  and (_07612_, _07611_, \oc8051_golden_model_1.ACC [3]);
  nor (_07613_, _07611_, \oc8051_golden_model_1.ACC [3]);
  not (_07614_, _05038_);
  and (_07615_, _04679_, \oc8051_golden_model_1.P2INREG [2]);
  and (_07616_, _04681_, \oc8051_golden_model_1.P3INREG [2]);
  or (_07617_, _07616_, _07615_);
  and (_07618_, _04673_, \oc8051_golden_model_1.P0INREG [2]);
  and (_07619_, _04676_, \oc8051_golden_model_1.P1INREG [2]);
  or (_07620_, _07619_, _07618_);
  nor (_07621_, _07620_, _07617_);
  and (_07622_, _07621_, _05072_);
  and (_07623_, _07622_, _05069_);
  nand (_07624_, _07623_, _05056_);
  nor (_07625_, _07624_, _07614_);
  and (_07626_, _07625_, \oc8051_golden_model_1.ACC [2]);
  not (_07627_, _04940_);
  and (_07628_, _04679_, \oc8051_golden_model_1.P2INREG [1]);
  and (_07629_, _04681_, \oc8051_golden_model_1.P3INREG [1]);
  or (_07630_, _07629_, _07628_);
  and (_07631_, _04673_, \oc8051_golden_model_1.P0INREG [1]);
  and (_07632_, _04676_, \oc8051_golden_model_1.P1INREG [1]);
  or (_07633_, _07632_, _07631_);
  nor (_07634_, _07633_, _07630_);
  and (_07635_, _07634_, _04974_);
  and (_07636_, _07635_, _04971_);
  nand (_07637_, _07636_, _04958_);
  nor (_07638_, _07637_, _07627_);
  and (_07639_, _07638_, \oc8051_golden_model_1.ACC [1]);
  nor (_07640_, _07638_, \oc8051_golden_model_1.ACC [1]);
  and (_07641_, _04679_, \oc8051_golden_model_1.P2INREG [0]);
  and (_07642_, _04681_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_07643_, _07642_, _07641_);
  and (_07644_, _04673_, \oc8051_golden_model_1.P0INREG [0]);
  and (_07645_, _04676_, \oc8051_golden_model_1.P1INREG [0]);
  nor (_07646_, _07645_, _07644_);
  and (_07647_, _07646_, _07643_);
  and (_07648_, _07647_, _04998_);
  and (_07649_, _07648_, _05016_);
  and (_07650_, _07649_, _05034_);
  and (_07651_, _07650_, _04989_);
  nor (_07652_, _07651_, \oc8051_golden_model_1.ACC [0]);
  nor (_07653_, _07652_, _07640_);
  or (_07654_, _07653_, _07639_);
  nor (_07655_, _07625_, \oc8051_golden_model_1.ACC [2]);
  nor (_07656_, _07655_, _07626_);
  and (_07657_, _07656_, _07654_);
  nor (_07658_, _07657_, _07626_);
  nor (_07659_, _07658_, _07613_);
  or (_07660_, _07659_, _07612_);
  nor (_07661_, _07593_, \oc8051_golden_model_1.ACC [4]);
  nor (_07662_, _07661_, _07594_);
  and (_07663_, _07662_, _07660_);
  nor (_07664_, _07663_, _07594_);
  nor (_07665_, _07664_, _07574_);
  or (_07666_, _07665_, _07573_);
  and (_07667_, _07666_, _07559_);
  nor (_07668_, _07667_, _07557_);
  and (_07669_, _07668_, _07545_);
  nor (_07670_, _07668_, _07545_);
  nor (_07671_, _07670_, _07669_);
  nor (_07672_, _07666_, _07559_);
  nor (_07673_, _07672_, _07667_);
  nor (_07674_, _07573_, _07574_);
  nor (_07675_, _07674_, _07664_);
  and (_07676_, _07674_, _07664_);
  or (_07677_, _07676_, _07675_);
  nor (_07678_, _07662_, _07660_);
  nor (_07679_, _07678_, _07663_);
  nor (_07680_, _07612_, _07613_);
  and (_07681_, _07680_, _07656_);
  nor (_07682_, _07639_, _07640_);
  and (_07683_, _07651_, \oc8051_golden_model_1.ACC [0]);
  nor (_07684_, _07683_, _07652_);
  and (_07685_, _07684_, _07682_);
  and (_07686_, _07685_, _07681_);
  and (_07687_, _07686_, \oc8051_golden_model_1.PSW [7]);
  not (_07688_, _07687_);
  nor (_07689_, _07688_, _07679_);
  not (_07690_, _07689_);
  nor (_07691_, _07690_, _07677_);
  not (_07692_, _07691_);
  nor (_07693_, _07692_, _07673_);
  and (_07694_, _07693_, _07671_);
  nor (_07695_, _07693_, _07671_);
  nor (_07696_, _07695_, _07694_);
  nand (_07697_, _07696_, _02898_);
  and (_07698_, _07697_, _07541_);
  and (_07699_, _07698_, _07539_);
  not (_07700_, _02499_);
  and (_07701_, _04614_, \oc8051_golden_model_1.PSW [7]);
  and (_07702_, _07701_, _04591_);
  and (_07703_, _07702_, _04646_);
  and (_07704_, _07703_, _02890_);
  and (_07705_, _07703_, _04340_);
  nor (_07706_, _07705_, _02743_);
  or (_07707_, _07706_, _07704_);
  nor (_07708_, _07707_, _05719_);
  and (_07709_, _07707_, _05719_);
  nor (_07710_, _07709_, _07708_);
  not (_07711_, _07710_);
  nor (_07712_, _07703_, _04340_);
  nor (_07713_, _07712_, _07705_);
  nor (_07714_, _07713_, _06762_);
  and (_07715_, _07713_, _06762_);
  and (_07716_, _07702_, _04597_);
  nor (_07717_, _07716_, _04621_);
  nor (_07718_, _07717_, _07703_);
  and (_07719_, _07718_, _06808_);
  nor (_07720_, _07718_, _06808_);
  nor (_07721_, _07702_, _04597_);
  nor (_07722_, _07721_, _07716_);
  nor (_07723_, _07722_, _06814_);
  nor (_07724_, _07723_, _07720_);
  nor (_07725_, _07724_, _07719_);
  nor (_07726_, _07720_, _07719_);
  and (_07727_, _07722_, _06814_);
  nor (_07728_, _07727_, _07723_);
  and (_07729_, _07728_, _07726_);
  not (_07730_, _07729_);
  nor (_07731_, _05501_, _02774_);
  nor (_07732_, _07731_, _07702_);
  and (_07733_, _07732_, _02605_);
  nor (_07734_, _07732_, _02605_);
  nor (_07735_, _07734_, _07733_);
  nor (_07736_, _07701_, _03321_);
  nor (_07737_, _07736_, _05501_);
  nor (_07738_, _07737_, _06908_);
  and (_07739_, _07737_, _06908_);
  nor (_07740_, _07739_, _07738_);
  and (_07741_, _07740_, _07735_);
  not (_07742_, _07741_);
  nor (_07743_, _02835_, _07294_);
  nor (_07744_, _07743_, _03743_);
  nor (_07745_, _07744_, _07701_);
  and (_07746_, _07745_, _02477_);
  nor (_07747_, _07745_, _02477_);
  and (_07748_, _02835_, _07294_);
  nor (_07749_, _07748_, _07743_);
  nor (_07750_, _07749_, _02658_);
  nor (_07751_, _07750_, _07747_);
  nor (_07752_, _07751_, _07746_);
  nor (_07753_, _07752_, _07742_);
  and (_07754_, _07739_, _07735_);
  nor (_07755_, _07754_, _07733_);
  not (_07756_, _07755_);
  nor (_07757_, _07756_, _07753_);
  and (_07758_, _07749_, _02658_);
  nor (_07759_, _07750_, _07758_);
  and (_07760_, _03742_, _02477_);
  nor (_07761_, _03742_, _02477_);
  nor (_07762_, _07761_, _07760_);
  and (_07763_, \oc8051_golden_model_1.PSW [7], _02658_);
  and (_07764_, _07294_, \oc8051_golden_model_1.ACC [0]);
  nor (_07765_, _07764_, _02835_);
  nor (_07766_, _07765_, _07763_);
  and (_07767_, _07766_, _07762_);
  nor (_07768_, _07766_, _07762_);
  nor (_07769_, _07768_, _07767_);
  nand (_07770_, _07769_, _07759_);
  nor (_07771_, _07770_, _07742_);
  nor (_07772_, _07771_, _07757_);
  nor (_07773_, _07772_, _07730_);
  nor (_07774_, _07773_, _07725_);
  nor (_07775_, _07774_, _07715_);
  or (_07776_, _07775_, _07714_);
  and (_07777_, _07776_, _07711_);
  nor (_07778_, _07776_, _07711_);
  or (_07779_, _07778_, _07777_);
  and (_07780_, _07779_, _07540_);
  or (_07781_, _07780_, _07700_);
  or (_07782_, _07781_, _07699_);
  nand (_07783_, _02743_, _07700_);
  and (_07784_, _07783_, _02966_);
  and (_07785_, _07784_, _07782_);
  not (_07786_, _05291_);
  nor (_07787_, _05502_, _07786_);
  nor (_07788_, _07787_, _07463_);
  nor (_07789_, _07788_, _02966_);
  or (_07790_, _07789_, _03861_);
  or (_07791_, _07790_, _07785_);
  and (_07792_, _07791_, _07328_);
  or (_07793_, _07792_, _03850_);
  and (_07794_, _07793_, _07324_);
  and (_07795_, _05706_, _04654_);
  nor (_07796_, _07795_, _07320_);
  nor (_07797_, _07796_, _02970_);
  or (_07798_, _07797_, _06731_);
  or (_07799_, _07798_, _07794_);
  not (_07800_, _06751_);
  nand (_07801_, _07800_, _06731_);
  and (_07802_, _07801_, _07799_);
  and (_07803_, _07802_, _02552_);
  nor (_07804_, _02743_, _02552_);
  or (_07805_, _07804_, _02974_);
  or (_07806_, _07805_, _07803_);
  and (_07807_, _02978_, _02584_);
  not (_07808_, _07807_);
  and (_07809_, _05517_, _04654_);
  nor (_07810_, _07809_, _07320_);
  nand (_07811_, _07810_, _02974_);
  and (_07812_, _07811_, _07808_);
  and (_07813_, _07812_, _07806_);
  nor (_07814_, _07808_, _02743_);
  and (_07815_, _02999_, _02581_);
  nor (_07816_, _07815_, _03259_);
  not (_07817_, _07816_);
  or (_07818_, _07817_, _07814_);
  or (_07819_, _07818_, _07813_);
  nor (_07820_, _07816_, _07196_);
  and (_07821_, _03680_, _02581_);
  nor (_07822_, _07821_, _03488_);
  not (_07823_, _07822_);
  nor (_07824_, _07823_, _07820_);
  and (_07825_, _07824_, _07819_);
  and (_07826_, _07823_, _07196_);
  and (_07827_, _03008_, _02581_);
  nor (_07828_, _07827_, _03484_);
  not (_07829_, _07828_);
  or (_07830_, _07829_, _07826_);
  or (_07831_, _07830_, _07825_);
  and (_07832_, _02971_, _02581_);
  not (_07833_, _07832_);
  or (_07834_, _07828_, _07196_);
  and (_07835_, _07834_, _07833_);
  and (_07836_, _07835_, _07831_);
  and (_07837_, _07147_, _07832_);
  or (_07838_, _07837_, _03105_);
  or (_07839_, _07838_, _07836_);
  or (_07840_, _05722_, _03106_);
  and (_07841_, _07840_, _07839_);
  or (_07842_, _07841_, _07319_);
  and (_07843_, _02743_, _05719_);
  nor (_07844_, _02743_, _05719_);
  nor (_07845_, _07844_, _07843_);
  not (_07846_, _07319_);
  or (_07847_, _07846_, _07845_);
  and (_07848_, _07847_, _07842_);
  or (_07849_, _07848_, _02977_);
  and (_07850_, _05259_, _04654_);
  nor (_07851_, _07850_, _07320_);
  nand (_07852_, _07851_, _02977_);
  and (_07853_, _07852_, _07104_);
  and (_07854_, _07853_, _07849_);
  and (_07855_, _07320_, _03107_);
  or (_07856_, _07855_, _07854_);
  not (_07857_, _02593_);
  nor (_07858_, _03012_, _07857_);
  and (_07859_, _03009_, _02593_);
  and (_07860_, _02912_, _02593_);
  or (_07861_, _07860_, _07859_);
  nor (_07862_, _07861_, _07858_);
  and (_07863_, _07862_, _07856_);
  not (_07864_, _03278_);
  and (_07865_, _07864_, _03227_);
  and (_07866_, _02904_, _02593_);
  not (_07867_, _07866_);
  and (_07868_, _07867_, _07865_);
  not (_07869_, _07868_);
  or (_07870_, _07195_, _03497_);
  and (_07871_, _07870_, _07869_);
  or (_07872_, _07871_, _07863_);
  or (_07873_, _07195_, _03498_);
  and (_07874_, _07873_, _07872_);
  or (_07875_, _07874_, _03499_);
  not (_07876_, _03499_);
  or (_07877_, _07146_, _07876_);
  and (_07878_, _07877_, _03093_);
  and (_07879_, _07878_, _07875_);
  and (_07880_, _02978_, _02593_);
  nor (_07881_, _07880_, _03092_);
  not (_07882_, _07881_);
  or (_07883_, _07880_, _05720_);
  and (_07884_, _07883_, _07882_);
  or (_07885_, _07884_, _07879_);
  not (_07886_, _07880_);
  or (_07887_, _07886_, _07844_);
  and (_07888_, _07887_, _03881_);
  and (_07889_, _07888_, _07885_);
  or (_07890_, _07810_, _05721_);
  nor (_07891_, _07890_, _03881_);
  or (_07892_, _07891_, _07317_);
  or (_07893_, _07892_, _07889_);
  and (_07894_, _07893_, _07318_);
  or (_07895_, _07894_, _07315_);
  nand (_07896_, _07145_, _07315_);
  and (_07897_, _07896_, _03098_);
  and (_07898_, _07897_, _07895_);
  and (_07899_, _02978_, _02588_);
  nor (_07900_, _07899_, _03097_);
  not (_07901_, _07900_);
  not (_07902_, _07899_);
  nand (_07903_, _07902_, _05721_);
  and (_07904_, _07903_, _07901_);
  or (_07905_, _07904_, _07898_);
  nand (_07906_, _07899_, _07843_);
  and (_07907_, _07906_, _07120_);
  and (_07908_, _07907_, _07905_);
  nor (_07909_, _05257_, _07325_);
  nor (_07910_, _07909_, _07320_);
  nor (_07911_, _07910_, _07120_);
  not (_07912_, _07241_);
  or (_07913_, _07912_, _07911_);
  or (_07914_, _07913_, _07908_);
  and (_07915_, _07914_, _07314_);
  or (_07916_, _07915_, _07236_);
  not (_07917_, _07236_);
  and (_07918_, _07342_, \oc8051_golden_model_1.ACC [6]);
  nor (_07919_, _07343_, _07344_);
  and (_07920_, _07348_, \oc8051_golden_model_1.ACC [5]);
  and (_07921_, _07354_, \oc8051_golden_model_1.ACC [4]);
  and (_07922_, _07365_, \oc8051_golden_model_1.ACC [3]);
  and (_07923_, _07370_, \oc8051_golden_model_1.ACC [2]);
  and (_07924_, _07377_, \oc8051_golden_model_1.ACC [1]);
  nor (_07925_, _07378_, _07379_);
  and (_07926_, _07381_, \oc8051_golden_model_1.ACC [0]);
  not (_07927_, _07926_);
  nor (_07928_, _07927_, _07925_);
  nor (_07929_, _07928_, _07924_);
  nor (_07930_, _07929_, _07373_);
  nor (_07931_, _07930_, _07923_);
  nor (_07932_, _07931_, _07368_);
  nor (_07933_, _07932_, _07922_);
  nor (_07934_, _07933_, _07360_);
  nor (_07935_, _07934_, _07921_);
  nor (_07936_, _07935_, _07358_);
  nor (_07937_, _07936_, _07920_);
  nor (_07938_, _07937_, _07919_);
  nor (_07939_, _07938_, _07918_);
  nor (_07940_, _07939_, _07338_);
  and (_07941_, _07939_, _07338_);
  nor (_07942_, _07941_, _07940_);
  or (_07943_, _07942_, _07917_);
  and (_07944_, _07943_, _03104_);
  and (_07945_, _07944_, _07916_);
  and (_07946_, _02978_, _02591_);
  nor (_07947_, _07946_, _03103_);
  not (_07948_, _07947_);
  not (_07949_, _07556_);
  not (_07950_, _07611_);
  not (_07951_, _07625_);
  not (_07952_, _07638_);
  nor (_07953_, _07651_, _07294_);
  and (_07954_, _07953_, _07952_);
  and (_07955_, _07954_, _07951_);
  and (_07956_, _07955_, _07950_);
  nor (_07957_, _07593_, _07572_);
  and (_07958_, _07957_, _07956_);
  and (_07959_, _07958_, _07949_);
  nor (_07960_, _07959_, _05466_);
  and (_07961_, _07959_, _05466_);
  nor (_07962_, _07961_, _07960_);
  and (_07963_, _07962_, \oc8051_golden_model_1.ACC [7]);
  nor (_07964_, _07962_, \oc8051_golden_model_1.ACC [7]);
  nor (_07965_, _07964_, _07963_);
  nor (_07966_, _07958_, _07949_);
  nor (_07967_, _07966_, _07959_);
  and (_07968_, _07967_, \oc8051_golden_model_1.ACC [6]);
  and (_07969_, _07967_, _06762_);
  nor (_07970_, _07967_, _06762_);
  nor (_07971_, _07970_, _07969_);
  not (_07972_, _07572_);
  not (_07973_, _07593_);
  and (_07974_, _07956_, _07973_);
  nor (_07975_, _07974_, _07972_);
  nor (_07976_, _07975_, _07958_);
  and (_07977_, _07976_, \oc8051_golden_model_1.ACC [5]);
  and (_07978_, _07976_, _06808_);
  nor (_07979_, _07976_, _06808_);
  nor (_07980_, _07979_, _07978_);
  nor (_07981_, _07956_, _07973_);
  nor (_07982_, _07981_, _07974_);
  and (_07983_, _07982_, \oc8051_golden_model_1.ACC [4]);
  nor (_07984_, _07982_, _06814_);
  and (_07985_, _07982_, _06814_);
  nor (_07986_, _07985_, _07984_);
  nor (_07987_, _07955_, _07950_);
  nor (_07988_, _07987_, _07956_);
  and (_07989_, _07988_, \oc8051_golden_model_1.ACC [3]);
  nor (_07990_, _07988_, _02605_);
  and (_07991_, _07988_, _02605_);
  nor (_07992_, _07991_, _07990_);
  nor (_07993_, _07954_, _07951_);
  nor (_07994_, _07993_, _07955_);
  and (_07995_, _07994_, \oc8051_golden_model_1.ACC [2]);
  nor (_07996_, _07994_, _06908_);
  and (_07997_, _07994_, _06908_);
  nor (_07998_, _07997_, _07996_);
  nor (_07999_, _07953_, _07952_);
  nor (_08000_, _07999_, _07954_);
  and (_08001_, _08000_, \oc8051_golden_model_1.ACC [1]);
  nor (_08002_, _08000_, _02477_);
  and (_08003_, _08000_, _02477_);
  nor (_08004_, _08003_, _08002_);
  and (_08005_, _07651_, _07294_);
  nor (_08006_, _08005_, _07953_);
  and (_08007_, _08006_, \oc8051_golden_model_1.ACC [0]);
  not (_08008_, _08007_);
  nor (_08009_, _08008_, _08004_);
  nor (_08010_, _08009_, _08001_);
  nor (_08011_, _08010_, _07998_);
  nor (_08012_, _08011_, _07995_);
  nor (_08013_, _08012_, _07992_);
  nor (_08014_, _08013_, _07989_);
  nor (_08015_, _08014_, _07986_);
  nor (_08016_, _08015_, _07983_);
  nor (_08017_, _08016_, _07980_);
  nor (_08018_, _08017_, _07977_);
  nor (_08019_, _08018_, _07971_);
  nor (_08020_, _08019_, _07968_);
  nor (_08021_, _08020_, _07965_);
  and (_08022_, _08020_, _07965_);
  nor (_08023_, _08022_, _08021_);
  or (_08024_, _08023_, _07946_);
  and (_08025_, _08024_, _07948_);
  or (_08026_, _08025_, _07945_);
  and (_08027_, _02591_, _02475_);
  not (_08028_, _08027_);
  not (_08029_, _07946_);
  and (_08030_, _07713_, \oc8051_golden_model_1.ACC [6]);
  nor (_08031_, _07714_, _07715_);
  and (_08032_, _07718_, \oc8051_golden_model_1.ACC [5]);
  and (_08033_, _07722_, \oc8051_golden_model_1.ACC [4]);
  and (_08034_, _07732_, \oc8051_golden_model_1.ACC [3]);
  and (_08035_, _07737_, \oc8051_golden_model_1.ACC [2]);
  and (_08036_, _07745_, \oc8051_golden_model_1.ACC [1]);
  nor (_08037_, _07747_, _07746_);
  and (_08038_, _07749_, \oc8051_golden_model_1.ACC [0]);
  not (_08039_, _08038_);
  nor (_08040_, _08039_, _08037_);
  nor (_08041_, _08040_, _08036_);
  nor (_08042_, _08041_, _07740_);
  nor (_08043_, _08042_, _08035_);
  nor (_08044_, _08043_, _07735_);
  nor (_08045_, _08044_, _08034_);
  nor (_08046_, _08045_, _07728_);
  nor (_08047_, _08046_, _08033_);
  nor (_08048_, _08047_, _07726_);
  nor (_08049_, _08048_, _08032_);
  nor (_08050_, _08049_, _08031_);
  nor (_08051_, _08050_, _08030_);
  nor (_08052_, _08051_, _07710_);
  and (_08053_, _08051_, _07710_);
  nor (_08054_, _08053_, _08052_);
  or (_08055_, _08054_, _08029_);
  and (_08056_, _08055_, _08028_);
  and (_08057_, _08056_, _08026_);
  not (_08058_, _03539_);
  and (_08059_, _07190_, _08058_);
  and (_08060_, _03008_, _02574_);
  not (_08061_, _08060_);
  and (_08062_, _08061_, _08059_);
  nand (_08063_, _08027_, \oc8051_golden_model_1.ACC [6]);
  nand (_08064_, _08063_, _08062_);
  or (_08065_, _08064_, _08057_);
  and (_08066_, _08065_, _07235_);
  not (_08067_, _03542_);
  nor (_08068_, _07233_, _08067_);
  or (_08069_, _08068_, _07183_);
  or (_08070_, _08069_, _08066_);
  and (_08071_, _08070_, _07184_);
  or (_08072_, _08071_, _02856_);
  and (_08073_, _02978_, _02574_);
  not (_08074_, _08073_);
  nor (_08075_, _07556_, _06762_);
  nor (_08076_, _07572_, _06808_);
  nor (_08077_, _07593_, _06814_);
  not (_08078_, _07662_);
  nor (_08079_, _07625_, _06908_);
  nor (_08080_, _07638_, _02477_);
  nor (_08081_, _07651_, _02658_);
  not (_08082_, _08081_);
  nor (_08083_, _08082_, _07682_);
  nor (_08084_, _08083_, _08080_);
  nor (_08085_, _08084_, _07656_);
  nor (_08086_, _08085_, _08079_);
  nor (_08087_, _08086_, _07611_);
  or (_08088_, _08087_, \oc8051_golden_model_1.ACC [3]);
  nand (_08089_, _08086_, _07611_);
  and (_08090_, _08089_, _08088_);
  and (_08091_, _08090_, _08078_);
  nor (_08092_, _08091_, _08077_);
  nor (_08093_, _08092_, _07674_);
  nor (_08094_, _08093_, _08076_);
  nor (_08095_, _08094_, _07559_);
  nor (_08096_, _08095_, _08075_);
  nor (_08097_, _08096_, _07544_);
  and (_08098_, _08096_, _07544_);
  nor (_08099_, _08098_, _08097_);
  nand (_08100_, _08099_, _02856_);
  and (_08101_, _08100_, _08074_);
  and (_08102_, _08101_, _08072_);
  nor (_08103_, _02889_, _06762_);
  and (_08104_, _02889_, _06762_);
  nor (_08105_, _08103_, _08104_);
  nor (_08106_, _03179_, _06808_);
  and (_08107_, _03179_, _06808_);
  nor (_08108_, _03620_, _06814_);
  and (_08109_, _03620_, _06814_);
  nor (_08110_, _08108_, _08109_);
  and (_08111_, _02774_, \oc8051_golden_model_1.ACC [3]);
  nor (_08112_, _02774_, \oc8051_golden_model_1.ACC [3]);
  nor (_08113_, _03320_, _06908_);
  and (_08114_, _03320_, _06908_);
  nor (_08115_, _08113_, _08114_);
  not (_08116_, _08115_);
  nor (_08117_, _02835_, _02658_);
  and (_08118_, _08117_, _07762_);
  nor (_08119_, _08118_, _07761_);
  nor (_08120_, _08119_, _08116_);
  nor (_08121_, _08120_, _08113_);
  nor (_08122_, _08121_, _08112_);
  or (_08123_, _08122_, _08111_);
  and (_08124_, _08123_, _08110_);
  nor (_08125_, _08124_, _08108_);
  nor (_08126_, _08125_, _08107_);
  or (_08127_, _08126_, _08106_);
  and (_08128_, _08127_, _08105_);
  nor (_08129_, _08128_, _08103_);
  nor (_08130_, _08129_, _07845_);
  and (_08131_, _08129_, _07845_);
  or (_08132_, _08131_, _08130_);
  and (_08133_, _08132_, _08073_);
  or (_08134_, _08133_, _07143_);
  or (_08135_, _08134_, _08102_);
  and (_08136_, _08135_, _07144_);
  or (_08137_, _08136_, _03133_);
  and (_08138_, _02978_, _02571_);
  not (_08139_, _08138_);
  nand (_08140_, _07404_, _03133_);
  and (_08141_, _08140_, _08139_);
  and (_08142_, _08141_, _08137_);
  and (_08143_, _02571_, _02475_);
  nor (_08144_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  and (_08145_, _08144_, _06855_);
  and (_08146_, _08145_, _06778_);
  and (_08147_, _08146_, _06762_);
  nor (_08148_, _08147_, _05719_);
  and (_08149_, _08147_, _05719_);
  nor (_08150_, _08149_, _08148_);
  nor (_08151_, _08150_, _08139_);
  or (_08152_, _08151_, _08143_);
  or (_08153_, _08152_, _08142_);
  nand (_08154_, _08143_, _07294_);
  and (_08155_, _08154_, _03142_);
  and (_08156_, _08155_, _08153_);
  nor (_08157_, _07494_, _03142_);
  or (_08158_, _08157_, _02852_);
  or (_08159_, _08158_, _08156_);
  and (_08160_, _02978_, _02567_);
  not (_08161_, _08160_);
  and (_08162_, _05196_, _04654_);
  nor (_08163_, _08162_, _07320_);
  nand (_08164_, _08163_, _02852_);
  and (_08165_, _08164_, _08161_);
  and (_08166_, _08165_, _08159_);
  and (_08167_, _02567_, _02475_);
  and (_08168_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.ACC [1]);
  nand (_08169_, _08168_, _06856_);
  nor (_08170_, _08169_, _06814_);
  and (_08171_, _08170_, \oc8051_golden_model_1.ACC [5]);
  and (_08172_, _08171_, \oc8051_golden_model_1.ACC [6]);
  nor (_08173_, _08172_, \oc8051_golden_model_1.ACC [7]);
  and (_08174_, _08172_, \oc8051_golden_model_1.ACC [7]);
  nor (_08175_, _08174_, _08173_);
  and (_08176_, _08175_, _08160_);
  or (_08177_, _08176_, _08167_);
  or (_08178_, _08177_, _08166_);
  nand (_08179_, _08167_, _02658_);
  and (_08180_, _08179_, _34446_);
  and (_08181_, _08180_, _08178_);
  or (_08182_, _08181_, _07142_);
  and (_35614_[7], _08182_, _35583_);
  or (_08183_, _34446_, \oc8051_golden_model_1.DPL [7]);
  and (_08184_, _08183_, _35583_);
  not (_08185_, \oc8051_golden_model_1.DPL [7]);
  nor (_08186_, _04670_, _08185_);
  and (_08187_, _05722_, _04670_);
  or (_08188_, _08187_, _08186_);
  and (_08189_, _08188_, _03107_);
  not (_08190_, _04670_);
  nor (_08191_, _08190_, _04585_);
  or (_08192_, _08191_, _08186_);
  or (_08193_, _08192_, _03860_);
  not (_08194_, _02975_);
  and (_08195_, _05439_, _04670_);
  or (_08196_, _08195_, _08186_);
  or (_08197_, _08196_, _06162_);
  and (_08198_, _04670_, \oc8051_golden_model_1.ACC [7]);
  or (_08199_, _08198_, _08186_);
  and (_08200_, _08199_, _02837_);
  nor (_08201_, _02837_, _08185_);
  or (_08202_, _08201_, _02932_);
  or (_08203_, _08202_, _08200_);
  and (_08204_, _08203_, _03693_);
  and (_08205_, _08204_, _08197_);
  and (_08206_, _08192_, _02930_);
  or (_08207_, _08206_, _02928_);
  or (_08208_, _08207_, _08205_);
  nor (_08209_, _02529_, _02474_);
  not (_08210_, _08209_);
  or (_08211_, _08199_, _02943_);
  and (_08212_, _08211_, _08210_);
  and (_08213_, _08212_, _08208_);
  and (_08214_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and (_08215_, _08214_, \oc8051_golden_model_1.DPL [2]);
  and (_08216_, _08215_, \oc8051_golden_model_1.DPL [3]);
  and (_08217_, _08216_, \oc8051_golden_model_1.DPL [4]);
  and (_08218_, _08217_, \oc8051_golden_model_1.DPL [5]);
  and (_08219_, _08218_, \oc8051_golden_model_1.DPL [6]);
  nor (_08220_, _08219_, \oc8051_golden_model_1.DPL [7]);
  and (_08221_, _08219_, \oc8051_golden_model_1.DPL [7]);
  nor (_08222_, _08221_, _08220_);
  and (_08223_, _08222_, _08209_);
  or (_08224_, _08223_, _08213_);
  and (_08225_, _08224_, _08194_);
  nor (_08226_, _05256_, _08194_);
  or (_08227_, _08226_, _03861_);
  or (_08228_, _08227_, _08225_);
  and (_08229_, _08228_, _08193_);
  or (_08230_, _08229_, _03850_);
  and (_08231_, _05426_, _04670_);
  or (_08232_, _08186_, _06726_);
  or (_08233_, _08232_, _08231_);
  and (_08234_, _08233_, _02970_);
  and (_08235_, _08234_, _08230_);
  and (_08236_, _05706_, _04670_);
  or (_08237_, _08236_, _08186_);
  and (_08238_, _08237_, _02524_);
  or (_08239_, _08238_, _02974_);
  or (_08240_, _08239_, _08235_);
  and (_08241_, _05517_, _04670_);
  or (_08242_, _08241_, _08186_);
  or (_08243_, _08242_, _05261_);
  and (_08244_, _08243_, _08240_);
  or (_08245_, _08244_, _02977_);
  and (_08246_, _05259_, _04670_);
  or (_08247_, _08186_, _07092_);
  or (_08248_, _08247_, _08246_);
  and (_08249_, _08248_, _07104_);
  and (_08250_, _08249_, _08245_);
  or (_08251_, _08250_, _08189_);
  and (_08252_, _08251_, _03095_);
  or (_08253_, _08186_, _04690_);
  and (_08254_, _08199_, _03094_);
  and (_08255_, _08242_, _02991_);
  or (_08256_, _08255_, _08254_);
  and (_08257_, _08256_, _08253_);
  or (_08258_, _08257_, _02994_);
  or (_08259_, _08258_, _08252_);
  nor (_08260_, _05257_, _08190_);
  or (_08261_, _08186_, _07120_);
  or (_08262_, _08261_, _08260_);
  and (_08263_, _08262_, _07118_);
  and (_08264_, _08263_, _08259_);
  nor (_08265_, _05721_, _08190_);
  or (_08266_, _08265_, _08186_);
  and (_08267_, _08266_, _03099_);
  or (_08268_, _08267_, _03133_);
  or (_08269_, _08268_, _08264_);
  or (_08270_, _08196_, _03138_);
  and (_08271_, _08270_, _02853_);
  and (_08272_, _08271_, _08269_);
  and (_08273_, _05196_, _04670_);
  or (_08274_, _08273_, _08186_);
  and (_08275_, _08274_, _02852_);
  or (_08276_, _08275_, _34450_);
  or (_08277_, _08276_, _08272_);
  and (_35617_[7], _08277_, _08184_);
  or (_08278_, _34446_, \oc8051_golden_model_1.DPH [7]);
  and (_08279_, _08278_, _35583_);
  not (_08280_, \oc8051_golden_model_1.DPH [7]);
  nor (_08281_, _05183_, _08280_);
  and (_08282_, _05722_, _04616_);
  or (_08283_, _08282_, _08281_);
  and (_08284_, _08283_, _03107_);
  not (_08285_, _04616_);
  nor (_08286_, _08285_, _04585_);
  or (_08287_, _08286_, _08281_);
  or (_08288_, _08287_, _03860_);
  and (_08289_, _05439_, _04616_);
  or (_08290_, _08289_, _08281_);
  or (_08291_, _08290_, _06162_);
  and (_08292_, _05183_, \oc8051_golden_model_1.ACC [7]);
  or (_08293_, _08292_, _08281_);
  and (_08294_, _08293_, _02837_);
  nor (_08295_, _02837_, _08280_);
  or (_08296_, _08295_, _02932_);
  or (_08297_, _08296_, _08294_);
  and (_08298_, _08297_, _03693_);
  and (_08299_, _08298_, _08291_);
  and (_08300_, _08287_, _02930_);
  or (_08301_, _08300_, _02928_);
  or (_08302_, _08301_, _08299_);
  or (_08303_, _08293_, _02943_);
  and (_08304_, _08303_, _08210_);
  and (_08305_, _08304_, _08302_);
  and (_08306_, _08221_, \oc8051_golden_model_1.DPH [0]);
  and (_08307_, _08306_, \oc8051_golden_model_1.DPH [1]);
  and (_08308_, _08307_, \oc8051_golden_model_1.DPH [2]);
  and (_08309_, _08308_, \oc8051_golden_model_1.DPH [3]);
  and (_08310_, _08309_, \oc8051_golden_model_1.DPH [4]);
  and (_08311_, _08310_, \oc8051_golden_model_1.DPH [5]);
  and (_08312_, _08311_, \oc8051_golden_model_1.DPH [6]);
  nand (_08313_, _08312_, \oc8051_golden_model_1.DPH [7]);
  or (_08314_, _08312_, \oc8051_golden_model_1.DPH [7]);
  and (_08315_, _08314_, _08313_);
  and (_08316_, _08315_, _08209_);
  or (_08317_, _08316_, _08305_);
  and (_08318_, _08317_, _08194_);
  nor (_08319_, _08194_, _02743_);
  or (_08320_, _08319_, _03861_);
  or (_08321_, _08320_, _08318_);
  and (_08322_, _08321_, _08288_);
  or (_08323_, _08322_, _03850_);
  or (_08324_, _08281_, _06726_);
  and (_08325_, _05426_, _05183_);
  or (_08326_, _08325_, _08324_);
  and (_08327_, _08326_, _02970_);
  and (_08328_, _08327_, _08323_);
  and (_08329_, _05706_, _05183_);
  or (_08330_, _08329_, _08281_);
  and (_08331_, _08330_, _02524_);
  or (_08332_, _08331_, _02974_);
  or (_08333_, _08332_, _08328_);
  and (_08334_, _05517_, _05183_);
  or (_08335_, _08334_, _08281_);
  or (_08336_, _08335_, _05261_);
  and (_08337_, _08336_, _08333_);
  or (_08338_, _08337_, _02977_);
  and (_08339_, _05259_, _04616_);
  or (_08340_, _08281_, _07092_);
  or (_08341_, _08340_, _08339_);
  and (_08342_, _08341_, _07104_);
  and (_08343_, _08342_, _08338_);
  or (_08344_, _08343_, _08284_);
  and (_08345_, _08344_, _03095_);
  or (_08346_, _08281_, _04690_);
  and (_08347_, _08293_, _03094_);
  and (_08348_, _08335_, _02991_);
  or (_08349_, _08348_, _08347_);
  and (_08350_, _08349_, _08346_);
  or (_08351_, _08350_, _02994_);
  or (_08352_, _08351_, _08345_);
  nor (_08353_, _05257_, _08285_);
  or (_08354_, _08281_, _07120_);
  or (_08355_, _08354_, _08353_);
  and (_08356_, _08355_, _07118_);
  and (_08357_, _08356_, _08352_);
  nor (_08358_, _05721_, _08285_);
  or (_08359_, _08358_, _08281_);
  and (_08360_, _08359_, _03099_);
  or (_08361_, _08360_, _03133_);
  or (_08362_, _08361_, _08357_);
  or (_08363_, _08290_, _03138_);
  and (_08364_, _08363_, _02853_);
  and (_08365_, _08364_, _08362_);
  and (_08366_, _05196_, _04616_);
  or (_08367_, _08366_, _08281_);
  and (_08368_, _08367_, _02852_);
  or (_08369_, _08368_, _34450_);
  or (_08370_, _08369_, _08365_);
  and (_35616_[7], _08370_, _08279_);
  and (_35618_[7], \oc8051_golden_model_1.IE [7], _35583_);
  and (_35619_[7], \oc8051_golden_model_1.IP [7], _35583_);
  not (_08371_, \oc8051_golden_model_1.P0 [7]);
  nor (_08372_, _34446_, _08371_);
  or (_08373_, _08372_, rst);
  nor (_08374_, _04673_, _08371_);
  and (_08375_, _05722_, _04673_);
  or (_08376_, _08375_, _08374_);
  and (_08377_, _08376_, _03107_);
  nor (_08378_, _04613_, _08371_);
  and (_08379_, _05444_, _04613_);
  or (_08380_, _08379_, _08378_);
  or (_08381_, _08378_, _05471_);
  and (_08382_, _08381_, _02790_);
  and (_08383_, _08382_, _08380_);
  and (_08384_, _05439_, _04673_);
  or (_08385_, _08384_, _08374_);
  or (_08386_, _08385_, _06162_);
  and (_08387_, _04673_, \oc8051_golden_model_1.ACC [7]);
  or (_08388_, _08387_, _08374_);
  and (_08389_, _08388_, _02837_);
  nor (_08390_, _02837_, _08371_);
  or (_08391_, _08390_, _02932_);
  or (_08392_, _08391_, _08389_);
  and (_08393_, _08392_, _02939_);
  and (_08394_, _08393_, _08386_);
  not (_08395_, _04673_);
  nor (_08396_, _08395_, _04585_);
  or (_08397_, _08396_, _08374_);
  and (_08398_, _08397_, _02930_);
  and (_08399_, _08380_, _02799_);
  or (_08400_, _08399_, _08398_);
  or (_08401_, _08400_, _02928_);
  or (_08402_, _08401_, _08394_);
  or (_08403_, _08388_, _02943_);
  and (_08404_, _08403_, _08402_);
  or (_08405_, _08404_, _02796_);
  and (_08406_, _05308_, _04613_);
  or (_08407_, _08406_, _08378_);
  or (_08408_, _08407_, _02927_);
  and (_08409_, _08408_, _06189_);
  and (_08410_, _08409_, _08405_);
  or (_08411_, _08410_, _08383_);
  and (_08412_, _08411_, _02966_);
  or (_08413_, _05501_, _05308_);
  and (_08414_, _08413_, _04613_);
  or (_08415_, _08414_, _08378_);
  and (_08416_, _08415_, _02785_);
  or (_08417_, _08416_, _03861_);
  or (_08418_, _08417_, _08412_);
  or (_08419_, _08397_, _03860_);
  and (_08420_, _08419_, _08418_);
  or (_08421_, _08420_, _03850_);
  and (_08422_, _05426_, _04673_);
  or (_08423_, _08374_, _06726_);
  or (_08424_, _08423_, _08422_);
  and (_08425_, _08424_, _02970_);
  and (_08426_, _08425_, _08421_);
  and (_08427_, _05706_, _04673_);
  or (_08428_, _08427_, _08374_);
  and (_08429_, _08428_, _02524_);
  or (_08430_, _08429_, _02974_);
  or (_08431_, _08430_, _08426_);
  and (_08432_, _05517_, _04673_);
  or (_08433_, _08432_, _08374_);
  or (_08434_, _08433_, _05261_);
  and (_08435_, _08434_, _08431_);
  or (_08436_, _08435_, _02977_);
  and (_08437_, _05259_, _04673_);
  or (_08438_, _08374_, _07092_);
  or (_08439_, _08438_, _08437_);
  and (_08440_, _08439_, _07104_);
  and (_08441_, _08440_, _08436_);
  or (_08442_, _08441_, _08377_);
  and (_08443_, _08442_, _03095_);
  or (_08444_, _08374_, _04690_);
  and (_08445_, _08388_, _03094_);
  and (_08446_, _08433_, _02991_);
  or (_08447_, _08446_, _08445_);
  and (_08448_, _08447_, _08444_);
  or (_08449_, _08448_, _02994_);
  or (_08450_, _08449_, _08443_);
  nor (_08451_, _05257_, _08395_);
  or (_08452_, _08374_, _07120_);
  or (_08453_, _08452_, _08451_);
  and (_08454_, _08453_, _07118_);
  and (_08455_, _08454_, _08450_);
  nor (_08456_, _05721_, _08395_);
  or (_08457_, _08456_, _08374_);
  and (_08458_, _08457_, _03099_);
  or (_08459_, _08458_, _03133_);
  or (_08460_, _08459_, _08455_);
  or (_08461_, _08385_, _03138_);
  and (_08462_, _08461_, _03142_);
  and (_08463_, _08462_, _08460_);
  and (_08464_, _08407_, _02778_);
  or (_08465_, _08464_, _02852_);
  or (_08466_, _08465_, _08463_);
  and (_08467_, _05196_, _04673_);
  or (_08468_, _08374_, _02853_);
  or (_08469_, _08468_, _08467_);
  and (_08470_, _08469_, _34446_);
  and (_08471_, _08470_, _08466_);
  or (_35621_[7], _08471_, _08373_);
  not (_08472_, \oc8051_golden_model_1.P1 [7]);
  nor (_08473_, _34446_, _08472_);
  or (_08474_, _08473_, rst);
  nor (_08475_, _04676_, _08472_);
  and (_08476_, _05722_, _04676_);
  or (_08477_, _08476_, _08475_);
  and (_08478_, _08477_, _03107_);
  and (_08479_, _05439_, _04676_);
  or (_08480_, _08479_, _08475_);
  or (_08481_, _08480_, _06162_);
  and (_08482_, _04676_, \oc8051_golden_model_1.ACC [7]);
  or (_08483_, _08482_, _08475_);
  and (_08484_, _08483_, _02837_);
  nor (_08485_, _02837_, _08472_);
  or (_08486_, _08485_, _02932_);
  or (_08487_, _08486_, _08484_);
  and (_08488_, _08487_, _02939_);
  and (_08489_, _08488_, _08481_);
  not (_08490_, _04676_);
  nor (_08491_, _08490_, _04585_);
  or (_08492_, _08491_, _08475_);
  and (_08493_, _08492_, _02930_);
  nor (_08494_, _05300_, _08472_);
  and (_08495_, _05444_, _05300_);
  or (_08496_, _08495_, _08494_);
  and (_08497_, _08496_, _02799_);
  or (_08498_, _08497_, _08493_);
  or (_08499_, _08498_, _02928_);
  or (_08500_, _08499_, _08489_);
  or (_08501_, _08483_, _02943_);
  and (_08502_, _08501_, _08500_);
  or (_08503_, _08502_, _02796_);
  and (_08504_, _05308_, _05300_);
  or (_08505_, _08504_, _08494_);
  or (_08506_, _08505_, _02927_);
  and (_08507_, _08506_, _06189_);
  and (_08508_, _08507_, _08503_);
  and (_08509_, _05472_, _05300_);
  or (_08510_, _08509_, _08494_);
  and (_08511_, _08510_, _02790_);
  or (_08512_, _08511_, _08508_);
  and (_08513_, _08512_, _02966_);
  and (_08514_, _08413_, _05300_);
  or (_08515_, _08514_, _08494_);
  and (_08516_, _08515_, _02785_);
  or (_08517_, _08516_, _03861_);
  or (_08518_, _08517_, _08513_);
  or (_08519_, _08492_, _03860_);
  and (_08520_, _08519_, _08518_);
  or (_08521_, _08520_, _03850_);
  and (_08522_, _05426_, _04676_);
  or (_08523_, _08475_, _06726_);
  or (_08524_, _08523_, _08522_);
  and (_08525_, _08524_, _02970_);
  and (_08526_, _08525_, _08521_);
  and (_08527_, _05706_, _04676_);
  or (_08528_, _08527_, _08475_);
  and (_08529_, _08528_, _02524_);
  or (_08530_, _08529_, _02974_);
  or (_08531_, _08530_, _08526_);
  and (_08532_, _05517_, _04676_);
  or (_08533_, _08532_, _08475_);
  or (_08534_, _08533_, _05261_);
  and (_08535_, _08534_, _08531_);
  or (_08536_, _08535_, _02977_);
  and (_08537_, _05259_, _04676_);
  or (_08538_, _08475_, _07092_);
  or (_08539_, _08538_, _08537_);
  and (_08540_, _08539_, _07104_);
  and (_08541_, _08540_, _08536_);
  or (_08542_, _08541_, _08478_);
  and (_08543_, _08542_, _03095_);
  or (_08544_, _08475_, _04690_);
  and (_08545_, _08483_, _03094_);
  and (_08546_, _08533_, _02991_);
  or (_08547_, _08546_, _08545_);
  and (_08548_, _08547_, _08544_);
  or (_08549_, _08548_, _02994_);
  or (_08550_, _08549_, _08543_);
  nor (_08551_, _05257_, _08490_);
  or (_08552_, _08475_, _07120_);
  or (_08553_, _08552_, _08551_);
  and (_08554_, _08553_, _07118_);
  and (_08555_, _08554_, _08550_);
  nor (_08556_, _05721_, _08490_);
  or (_08557_, _08556_, _08475_);
  and (_08558_, _08557_, _03099_);
  or (_08559_, _08558_, _03133_);
  or (_08560_, _08559_, _08555_);
  or (_08561_, _08480_, _03138_);
  and (_08562_, _08561_, _03142_);
  and (_08563_, _08562_, _08560_);
  and (_08564_, _08505_, _02778_);
  or (_08565_, _08564_, _02852_);
  or (_08566_, _08565_, _08563_);
  and (_08567_, _05196_, _04676_);
  or (_08568_, _08475_, _02853_);
  or (_08569_, _08568_, _08567_);
  and (_08570_, _08569_, _34446_);
  and (_08571_, _08570_, _08566_);
  or (_35623_[7], _08571_, _08474_);
  not (_08572_, \oc8051_golden_model_1.P2 [7]);
  nor (_08573_, _34446_, _08572_);
  or (_08574_, _08573_, rst);
  nor (_08575_, _04679_, _08572_);
  and (_08576_, _05722_, _04679_);
  or (_08577_, _08576_, _08575_);
  and (_08578_, _08577_, _03107_);
  nor (_08579_, _05278_, _08572_);
  and (_08580_, _05444_, _05278_);
  or (_08581_, _08580_, _08579_);
  or (_08582_, _08579_, _05471_);
  and (_08583_, _08582_, _02790_);
  and (_08584_, _08583_, _08581_);
  and (_08585_, _05439_, _04679_);
  or (_08586_, _08585_, _08575_);
  or (_08587_, _08586_, _06162_);
  and (_08588_, _04679_, \oc8051_golden_model_1.ACC [7]);
  or (_08589_, _08588_, _08575_);
  and (_08590_, _08589_, _02837_);
  nor (_08591_, _02837_, _08572_);
  or (_08592_, _08591_, _02932_);
  or (_08593_, _08592_, _08590_);
  and (_08594_, _08593_, _02939_);
  and (_08595_, _08594_, _08587_);
  not (_08596_, _04679_);
  nor (_08597_, _08596_, _04585_);
  or (_08598_, _08597_, _08575_);
  and (_08599_, _08598_, _02930_);
  and (_08600_, _08581_, _02799_);
  or (_08601_, _08600_, _08599_);
  or (_08602_, _08601_, _02928_);
  or (_08603_, _08602_, _08595_);
  or (_08604_, _08589_, _02943_);
  and (_08605_, _08604_, _08603_);
  or (_08606_, _08605_, _02796_);
  and (_08607_, _05308_, _05278_);
  or (_08608_, _08607_, _08579_);
  or (_08609_, _08608_, _02927_);
  and (_08610_, _08609_, _06189_);
  and (_08611_, _08610_, _08606_);
  or (_08612_, _08611_, _08584_);
  and (_08613_, _08612_, _02966_);
  and (_08614_, _08413_, _05278_);
  or (_08615_, _08614_, _08579_);
  and (_08616_, _08615_, _02785_);
  or (_08617_, _08616_, _03861_);
  or (_08618_, _08617_, _08613_);
  or (_08619_, _08598_, _03860_);
  and (_08620_, _08619_, _08618_);
  or (_08621_, _08620_, _03850_);
  and (_08622_, _05426_, _04679_);
  or (_08623_, _08575_, _06726_);
  or (_08624_, _08623_, _08622_);
  and (_08625_, _08624_, _02970_);
  and (_08626_, _08625_, _08621_);
  and (_08627_, _05706_, _04679_);
  or (_08628_, _08627_, _08575_);
  and (_08629_, _08628_, _02524_);
  or (_08630_, _08629_, _02974_);
  or (_08631_, _08630_, _08626_);
  and (_08632_, _05517_, _04679_);
  or (_08633_, _08632_, _08575_);
  or (_08634_, _08633_, _05261_);
  and (_08635_, _08634_, _08631_);
  or (_08636_, _08635_, _02977_);
  and (_08637_, _05259_, _04679_);
  or (_08638_, _08575_, _07092_);
  or (_08639_, _08638_, _08637_);
  and (_08640_, _08639_, _07104_);
  and (_08641_, _08640_, _08636_);
  or (_08642_, _08641_, _08578_);
  and (_08643_, _08642_, _03095_);
  or (_08644_, _08575_, _04690_);
  and (_08645_, _08589_, _03094_);
  and (_08646_, _08633_, _02991_);
  or (_08647_, _08646_, _08645_);
  and (_08648_, _08647_, _08644_);
  or (_08649_, _08648_, _02994_);
  or (_08650_, _08649_, _08643_);
  nor (_08651_, _05257_, _08596_);
  or (_08652_, _08575_, _07120_);
  or (_08653_, _08652_, _08651_);
  and (_08654_, _08653_, _07118_);
  and (_08655_, _08654_, _08650_);
  nor (_08656_, _05721_, _08596_);
  or (_08657_, _08656_, _08575_);
  and (_08658_, _08657_, _03099_);
  or (_08659_, _08658_, _03133_);
  or (_08660_, _08659_, _08655_);
  or (_08661_, _08586_, _03138_);
  and (_08662_, _08661_, _03142_);
  and (_08663_, _08662_, _08660_);
  and (_08664_, _08608_, _02778_);
  or (_08665_, _08664_, _02852_);
  or (_08666_, _08665_, _08663_);
  and (_08667_, _05196_, _04679_);
  or (_08668_, _08575_, _02853_);
  or (_08669_, _08668_, _08667_);
  and (_08670_, _08669_, _34446_);
  and (_08671_, _08670_, _08666_);
  or (_35625_[7], _08671_, _08574_);
  not (_08672_, \oc8051_golden_model_1.P3 [7]);
  nor (_08673_, _34446_, _08672_);
  or (_08674_, _08673_, rst);
  nor (_08675_, _04681_, _08672_);
  and (_08676_, _05722_, _04681_);
  or (_08677_, _08676_, _08675_);
  and (_08678_, _08677_, _03107_);
  and (_08679_, _05439_, _04681_);
  or (_08680_, _08679_, _08675_);
  or (_08681_, _08680_, _06162_);
  and (_08682_, _04681_, \oc8051_golden_model_1.ACC [7]);
  or (_08683_, _08682_, _08675_);
  and (_08684_, _08683_, _02837_);
  nor (_08685_, _02837_, _08672_);
  or (_08686_, _08685_, _02932_);
  or (_08687_, _08686_, _08684_);
  and (_08688_, _08687_, _02939_);
  and (_08689_, _08688_, _08681_);
  not (_08690_, _04681_);
  nor (_08691_, _08690_, _04585_);
  or (_08692_, _08691_, _08675_);
  and (_08693_, _08692_, _02930_);
  nor (_08694_, _05280_, _08672_);
  and (_08695_, _05444_, _05280_);
  or (_08696_, _08695_, _08694_);
  and (_08697_, _08696_, _02799_);
  or (_08698_, _08697_, _08693_);
  or (_08699_, _08698_, _02928_);
  or (_08700_, _08699_, _08689_);
  or (_08701_, _08683_, _02943_);
  and (_08702_, _08701_, _08700_);
  or (_08703_, _08702_, _02796_);
  and (_08704_, _05308_, _05280_);
  or (_08705_, _08704_, _08694_);
  or (_08706_, _08705_, _02927_);
  and (_08707_, _08706_, _06189_);
  and (_08708_, _08707_, _08703_);
  and (_08709_, _05472_, _05280_);
  or (_08710_, _08709_, _08694_);
  and (_08711_, _08710_, _02790_);
  or (_08712_, _08711_, _08708_);
  and (_08713_, _08712_, _02966_);
  and (_08714_, _08413_, _05280_);
  or (_08715_, _08714_, _08694_);
  and (_08716_, _08715_, _02785_);
  or (_08717_, _08716_, _03861_);
  or (_08718_, _08717_, _08713_);
  or (_08719_, _08692_, _03860_);
  and (_08720_, _08719_, _08718_);
  or (_08721_, _08720_, _03850_);
  and (_08722_, _05426_, _04681_);
  or (_08723_, _08675_, _06726_);
  or (_08724_, _08723_, _08722_);
  and (_08725_, _08724_, _02970_);
  and (_08726_, _08725_, _08721_);
  and (_08727_, _05706_, _04681_);
  or (_08728_, _08727_, _08675_);
  and (_08729_, _08728_, _02524_);
  or (_08730_, _08729_, _02974_);
  or (_08731_, _08730_, _08726_);
  and (_08732_, _05517_, _04681_);
  or (_08733_, _08732_, _08675_);
  or (_08734_, _08733_, _05261_);
  and (_08735_, _08734_, _08731_);
  or (_08736_, _08735_, _02977_);
  and (_08737_, _05259_, _04681_);
  or (_08738_, _08675_, _07092_);
  or (_08739_, _08738_, _08737_);
  and (_08740_, _08739_, _07104_);
  and (_08741_, _08740_, _08736_);
  or (_08742_, _08741_, _08678_);
  and (_08743_, _08742_, _03095_);
  or (_08744_, _08675_, _04690_);
  and (_08745_, _08683_, _03094_);
  and (_08746_, _08733_, _02991_);
  or (_08747_, _08746_, _08745_);
  and (_08748_, _08747_, _08744_);
  or (_08749_, _08748_, _02994_);
  or (_08750_, _08749_, _08743_);
  nor (_08751_, _05257_, _08690_);
  or (_08752_, _08675_, _07120_);
  or (_08753_, _08752_, _08751_);
  and (_08754_, _08753_, _07118_);
  and (_08755_, _08754_, _08750_);
  nor (_08756_, _05721_, _08690_);
  or (_08757_, _08756_, _08675_);
  and (_08758_, _08757_, _03099_);
  or (_08759_, _08758_, _03133_);
  or (_08760_, _08759_, _08755_);
  or (_08761_, _08680_, _03138_);
  and (_08762_, _08761_, _03142_);
  and (_08763_, _08762_, _08760_);
  and (_08764_, _08705_, _02778_);
  or (_08765_, _08764_, _02852_);
  or (_08766_, _08765_, _08763_);
  and (_08767_, _05196_, _04681_);
  or (_08768_, _08675_, _02853_);
  or (_08769_, _08768_, _08767_);
  and (_08770_, _08769_, _34446_);
  and (_08771_, _08770_, _08766_);
  or (_35627_[7], _08771_, _08674_);
  or (_08772_, _08073_, _02856_);
  and (_08773_, _06136_, \oc8051_golden_model_1.PC [10]);
  not (_08774_, _02212_);
  and (_08775_, _05314_, _08774_);
  and (_08776_, _08775_, \oc8051_golden_model_1.PC [7]);
  and (_08777_, _08776_, _08773_);
  and (_08778_, _08777_, \oc8051_golden_model_1.PC [11]);
  and (_08779_, _08778_, \oc8051_golden_model_1.PC [12]);
  and (_08780_, _08779_, \oc8051_golden_model_1.PC [13]);
  and (_08781_, _08780_, \oc8051_golden_model_1.PC [14]);
  nor (_08782_, _08781_, \oc8051_golden_model_1.PC [15]);
  and (_08783_, _08776_, \oc8051_golden_model_1.PC [8]);
  and (_08784_, _08783_, \oc8051_golden_model_1.PC [9]);
  and (_08785_, _08784_, \oc8051_golden_model_1.PC [10]);
  and (_08786_, _08785_, \oc8051_golden_model_1.PC [11]);
  and (_08787_, _08786_, \oc8051_golden_model_1.PC [12]);
  and (_08788_, _08787_, \oc8051_golden_model_1.PC [13]);
  and (_08789_, _08788_, \oc8051_golden_model_1.PC [14]);
  and (_08790_, _08789_, \oc8051_golden_model_1.PC [15]);
  nor (_08791_, _08790_, _08782_);
  not (_08792_, _07183_);
  nor (_08793_, _07191_, _03702_);
  and (_08794_, _08793_, _08792_);
  and (_08795_, _08794_, _03544_);
  or (_08796_, _08795_, _08791_);
  and (_08797_, _07241_, _07917_);
  or (_08798_, _08797_, _08791_);
  and (_08799_, _02777_, _02588_);
  not (_08800_, _08799_);
  nor (_08801_, _03099_, _02589_);
  or (_08802_, _08801_, _06154_);
  and (_08803_, _08802_, _08800_);
  not (_08804_, _07315_);
  and (_08805_, _07316_, _08804_);
  or (_08806_, _08805_, _08791_);
  and (_08807_, _02777_, _02593_);
  not (_08808_, _08807_);
  nor (_08809_, _03094_, _02594_);
  or (_08810_, _08809_, _06154_);
  and (_08811_, _08810_, _08808_);
  and (_08812_, _07868_, _07876_);
  or (_08813_, _08812_, _08791_);
  nor (_08814_, _07319_, _03105_);
  not (_08815_, _08814_);
  and (_08816_, _03011_, _02581_);
  or (_08817_, _08816_, _03488_);
  nor (_08818_, _08817_, _07817_);
  and (_08819_, _03857_, _02581_);
  not (_08820_, _08819_);
  and (_08821_, _08820_, _08818_);
  and (_08822_, _08821_, _07833_);
  or (_08823_, _08822_, _08791_);
  or (_08824_, _06731_, _02476_);
  not (_08825_, _08824_);
  or (_08826_, _08825_, _08791_);
  nor (_08827_, _02532_, _02474_);
  not (_08828_, _08827_);
  and (_08829_, _02835_, _02658_);
  nor (_08830_, _08829_, _08117_);
  nor (_08831_, _08830_, _07762_);
  nor (_08832_, _08111_, _08112_);
  nor (_08833_, _08832_, _08115_);
  nor (_08834_, _08106_, _08107_);
  nor (_08835_, _08834_, _08110_);
  nor (_08836_, _08105_, _07845_);
  and (_08837_, _08836_, _08835_);
  and (_08838_, _08837_, _08833_);
  and (_08839_, _08838_, _08831_);
  nor (_08840_, _06141_, \oc8051_golden_model_1.PC [14]);
  nor (_08841_, _08840_, _06142_);
  not (_08842_, _08841_);
  nor (_08843_, _08842_, _05256_);
  and (_08844_, _08842_, _05256_);
  nor (_08845_, _08844_, _08843_);
  not (_08846_, _08845_);
  nor (_08847_, _06140_, \oc8051_golden_model_1.PC [13]);
  nor (_08848_, _08847_, _06141_);
  not (_08849_, _08848_);
  nor (_08850_, _08849_, _05256_);
  and (_08851_, _08849_, _05256_);
  nor (_08852_, _06139_, \oc8051_golden_model_1.PC [12]);
  nor (_08853_, _08852_, _06140_);
  not (_08854_, _08853_);
  nor (_08855_, _08854_, _05256_);
  and (_08856_, _08773_, _06096_);
  nor (_08857_, _08856_, \oc8051_golden_model_1.PC [11]);
  nor (_08858_, _08857_, _06139_);
  not (_08859_, _08858_);
  nor (_08860_, _08859_, _05256_);
  and (_08861_, _08859_, _05256_);
  nor (_08862_, _08861_, _08860_);
  and (_08863_, _06136_, _06096_);
  nor (_08864_, _08863_, \oc8051_golden_model_1.PC [10]);
  nor (_08865_, _08864_, _08856_);
  not (_08866_, _08865_);
  nor (_08867_, _08866_, _05256_);
  and (_08868_, _08866_, _05256_);
  nor (_08869_, _08868_, _08867_);
  and (_08870_, _08869_, _08862_);
  and (_08871_, _06096_, \oc8051_golden_model_1.PC [8]);
  nor (_08872_, _08871_, \oc8051_golden_model_1.PC [9]);
  nor (_08873_, _08872_, _08863_);
  not (_08874_, _08873_);
  nor (_08875_, _08874_, _05256_);
  and (_08876_, _08874_, _05256_);
  nor (_08877_, _08876_, _08875_);
  not (_08878_, _06098_);
  nor (_08879_, _05256_, _08878_);
  and (_08880_, _05256_, _08878_);
  nor (_08881_, _08880_, _08879_);
  not (_08882_, _08881_);
  and (_08883_, _06094_, _05313_);
  nor (_08884_, _08883_, \oc8051_golden_model_1.PC [6]);
  nor (_08885_, _08884_, _06095_);
  not (_08886_, _08885_);
  nor (_08887_, _08886_, _05549_);
  and (_08888_, _08886_, _05549_);
  nor (_08889_, _08888_, _08887_);
  and (_08890_, _06094_, \oc8051_golden_model_1.PC [4]);
  nor (_08891_, _08890_, \oc8051_golden_model_1.PC [5]);
  nor (_08892_, _08891_, _08883_);
  not (_08893_, _08892_);
  nor (_08894_, _08893_, _05612_);
  and (_08895_, _08893_, _05612_);
  nor (_08896_, _06094_, \oc8051_golden_model_1.PC [4]);
  nor (_08897_, _08896_, _08890_);
  not (_08898_, _08897_);
  nor (_08899_, _08898_, _05581_);
  nor (_08900_, _06093_, \oc8051_golden_model_1.PC [3]);
  nor (_08901_, _08900_, _06094_);
  not (_08902_, _08901_);
  nor (_08903_, _08902_, _03087_);
  and (_08904_, _08902_, _03087_);
  nor (_08905_, _02229_, \oc8051_golden_model_1.PC [2]);
  nor (_08906_, _08905_, _06093_);
  not (_08907_, _08906_);
  nor (_08908_, _08907_, _03223_);
  not (_08909_, _02478_);
  nor (_08910_, _03660_, _08909_);
  nor (_08911_, _03471_, \oc8051_golden_model_1.PC [0]);
  and (_08912_, _03660_, _08909_);
  nor (_08913_, _08912_, _08910_);
  and (_08914_, _08913_, _08911_);
  nor (_08915_, _08914_, _08910_);
  and (_08916_, _08907_, _03223_);
  nor (_08917_, _08916_, _08908_);
  not (_08918_, _08917_);
  nor (_08919_, _08918_, _08915_);
  nor (_08920_, _08919_, _08908_);
  nor (_08921_, _08920_, _08904_);
  nor (_08922_, _08921_, _08903_);
  and (_08923_, _08898_, _05581_);
  nor (_08924_, _08923_, _08899_);
  not (_08925_, _08924_);
  nor (_08926_, _08925_, _08922_);
  nor (_08927_, _08926_, _08899_);
  nor (_08928_, _08927_, _08895_);
  or (_08929_, _08928_, _08894_);
  and (_08930_, _08929_, _08889_);
  nor (_08931_, _08930_, _08887_);
  nor (_08932_, _08931_, _08882_);
  nor (_08933_, _08932_, _08879_);
  nor (_08934_, _06096_, \oc8051_golden_model_1.PC [8]);
  nor (_08935_, _08934_, _08871_);
  not (_08936_, _08935_);
  nor (_08937_, _08936_, _05256_);
  and (_08938_, _08936_, _05256_);
  nor (_08939_, _08938_, _08937_);
  not (_08940_, _08939_);
  nor (_08941_, _08940_, _08933_);
  and (_08942_, _08941_, _08877_);
  and (_08943_, _08942_, _08870_);
  nor (_08944_, _08937_, _08875_);
  not (_08945_, _08944_);
  and (_08946_, _08945_, _08870_);
  or (_08947_, _08946_, _08867_);
  or (_08948_, _08947_, _08943_);
  nor (_08949_, _08948_, _08860_);
  and (_08950_, _08854_, _05256_);
  nor (_08951_, _08950_, _08855_);
  not (_08952_, _08951_);
  nor (_08953_, _08952_, _08949_);
  nor (_08954_, _08953_, _08855_);
  nor (_08955_, _08954_, _08851_);
  nor (_08956_, _08955_, _08850_);
  nor (_08957_, _08956_, _08846_);
  nor (_08958_, _08957_, _08843_);
  and (_08959_, _06146_, _05256_);
  nor (_08960_, _06146_, _05256_);
  nor (_08961_, _08960_, _08959_);
  and (_08962_, _08961_, _08958_);
  nor (_08963_, _08961_, _08958_);
  or (_08964_, _08963_, _08962_);
  or (_08965_, _08964_, _08839_);
  nand (_08966_, _08839_, _06146_);
  and (_08967_, _08966_, _02979_);
  and (_08968_, _08967_, _08965_);
  not (_08969_, _02979_);
  not (_08970_, _05483_);
  or (_08971_, _06027_, _04621_);
  and (_08972_, _08971_, _08970_);
  nand (_08973_, _05798_, _02889_);
  or (_08974_, _05426_, _02743_);
  or (_08975_, _05798_, _02889_);
  and (_08976_, _08975_, _08974_);
  and (_08977_, _08976_, _08973_);
  and (_08978_, _08977_, _08972_);
  or (_08979_, _06072_, _04597_);
  or (_08980_, _06120_, _03179_);
  or (_08981_, _06121_, _03620_);
  and (_08982_, _08981_, _08980_);
  and (_08983_, _08982_, _08979_);
  and (_08984_, _08983_, _08978_);
  or (_08985_, _06116_, _04318_);
  or (_08986_, _05935_, _02774_);
  and (_08987_, _08986_, _08985_);
  and (_08988_, _05980_, _03321_);
  and (_08989_, _06117_, _03320_);
  nor (_08990_, _08989_, _08988_);
  and (_08991_, _08990_, _08987_);
  or (_08992_, _05889_, _02836_);
  and (_08993_, _05844_, _03743_);
  and (_08994_, _06113_, _03742_);
  nor (_08995_, _08994_, _08993_);
  and (_08996_, _08995_, _08992_);
  and (_08997_, _08996_, _08991_);
  or (_08998_, _06114_, _02835_);
  and (_08999_, _08998_, _08997_);
  and (_09000_, _08999_, _08984_);
  or (_09001_, _09000_, _08964_);
  nand (_09002_, _09000_, _06146_);
  and (_09003_, _09002_, _09001_);
  and (_09004_, _09003_, _02972_);
  and (_09005_, _07674_, _07662_);
  and (_09006_, _07559_, _07545_);
  and (_09007_, _09006_, _09005_);
  and (_09008_, _09007_, _07686_);
  not (_09009_, _09008_);
  and (_09010_, _09009_, _08964_);
  and (_09011_, _09008_, _06145_);
  or (_09012_, _09011_, _09010_);
  and (_09013_, _09012_, _02944_);
  nor (_09014_, _02799_, _04239_);
  and (_09015_, _09014_, _03693_);
  or (_09016_, _09015_, _06154_);
  nor (_09017_, _02539_, _02474_);
  nor (_09018_, _09017_, _07402_);
  and (_09019_, _05036_, _04987_);
  and (_09020_, _05433_, _09019_);
  and (_09021_, _04783_, _04689_);
  and (_09022_, _09021_, _05430_);
  nand (_09023_, _09022_, _09020_);
  or (_09024_, _09023_, _06145_);
  and (_09025_, _09022_, _09020_);
  or (_09026_, _09025_, _08964_);
  and (_09027_, _09026_, _02932_);
  and (_09028_, _09027_, _09024_);
  nor (_09029_, _06150_, \oc8051_golden_model_1.PC [14]);
  nor (_09030_, _09029_, _06151_);
  not (_09031_, _09030_);
  nor (_09032_, _09031_, _02743_);
  and (_09033_, _09031_, _02743_);
  nor (_09034_, _09033_, _09032_);
  not (_09035_, _09034_);
  nor (_09036_, _06149_, \oc8051_golden_model_1.PC [13]);
  nor (_09037_, _09036_, _06150_);
  not (_09038_, _09037_);
  and (_09039_, _09038_, _02743_);
  nor (_09040_, _09038_, _02743_);
  not (_09041_, _09040_);
  nor (_09042_, _06148_, \oc8051_golden_model_1.PC [12]);
  nor (_09043_, _09042_, _06149_);
  not (_09044_, _09043_);
  nor (_09045_, _09044_, _02743_);
  and (_09046_, _08773_, _05316_);
  nor (_09047_, _09046_, \oc8051_golden_model_1.PC [11]);
  nor (_09048_, _09047_, _06148_);
  not (_09049_, _09048_);
  nor (_09050_, _09049_, _02743_);
  and (_09051_, _09049_, _02743_);
  and (_09052_, _06136_, _05316_);
  nor (_09053_, _09052_, \oc8051_golden_model_1.PC [10]);
  nor (_09054_, _09053_, _09046_);
  not (_09055_, _09054_);
  nor (_09056_, _09055_, _02743_);
  and (_09057_, _09055_, _02743_);
  nor (_09058_, _09057_, _09056_);
  and (_09059_, _05316_, \oc8051_golden_model_1.PC [8]);
  nor (_09060_, _09059_, \oc8051_golden_model_1.PC [9]);
  nor (_09061_, _09060_, _09052_);
  not (_09062_, _09061_);
  and (_09063_, _09062_, _02743_);
  nor (_09064_, _09062_, _02743_);
  not (_09065_, _09064_);
  nor (_09066_, _05316_, \oc8051_golden_model_1.PC [8]);
  nor (_09067_, _09066_, _09059_);
  not (_09068_, _09067_);
  nor (_09069_, _09068_, _02743_);
  nor (_09070_, _05476_, _02743_);
  and (_09071_, _05476_, _02743_);
  nor (_09072_, _09071_, _09070_);
  not (_09073_, _09072_);
  and (_09074_, _05313_, _02618_);
  nor (_09075_, _09074_, \oc8051_golden_model_1.PC [6]);
  nor (_09076_, _09075_, _05315_);
  not (_09077_, _09076_);
  nor (_09078_, _09077_, _02889_);
  and (_09079_, _09077_, _02889_);
  nor (_09080_, _09079_, _09078_);
  and (_09081_, _02618_, \oc8051_golden_model_1.PC [4]);
  nor (_09082_, _09081_, \oc8051_golden_model_1.PC [5]);
  nor (_09083_, _09082_, _09074_);
  not (_09084_, _09083_);
  nor (_09085_, _09084_, _03179_);
  and (_09086_, _09084_, _03179_);
  nor (_09087_, _02618_, \oc8051_golden_model_1.PC [4]);
  nor (_09088_, _09087_, _09081_);
  not (_09089_, _09088_);
  nor (_09090_, _09089_, _03620_);
  and (_09091_, _02774_, _02620_);
  nor (_09092_, _02774_, _02620_);
  nor (_09093_, _03320_, _02600_);
  nor (_09094_, _03742_, \oc8051_golden_model_1.PC [1]);
  nor (_09095_, _02835_, _02225_);
  and (_09096_, _03742_, \oc8051_golden_model_1.PC [1]);
  nor (_09097_, _09096_, _09094_);
  and (_09098_, _09097_, _09095_);
  nor (_09099_, _09098_, _09094_);
  and (_09100_, _03320_, _02600_);
  nor (_09101_, _09100_, _09093_);
  not (_09102_, _09101_);
  nor (_09103_, _09102_, _09099_);
  nor (_09104_, _09103_, _09093_);
  nor (_09105_, _09104_, _09092_);
  nor (_09106_, _09105_, _09091_);
  and (_09107_, _09089_, _03620_);
  nor (_09108_, _09107_, _09090_);
  not (_09109_, _09108_);
  nor (_09110_, _09109_, _09106_);
  nor (_09111_, _09110_, _09090_);
  nor (_09112_, _09111_, _09086_);
  or (_09113_, _09112_, _09085_);
  and (_09114_, _09113_, _09080_);
  nor (_09115_, _09114_, _09078_);
  nor (_09116_, _09115_, _09073_);
  nor (_09117_, _09116_, _09070_);
  and (_09118_, _09068_, _02743_);
  nor (_09119_, _09118_, _09069_);
  not (_09120_, _09119_);
  nor (_09121_, _09120_, _09117_);
  nor (_09122_, _09121_, _09069_);
  and (_09123_, _09122_, _09065_);
  or (_09124_, _09123_, _09063_);
  not (_09125_, _09124_);
  and (_09126_, _09125_, _09058_);
  nor (_09127_, _09126_, _09056_);
  nor (_09128_, _09127_, _09051_);
  or (_09129_, _09128_, _09050_);
  and (_09130_, _09044_, _02743_);
  nor (_09131_, _09130_, _09045_);
  and (_09132_, _09131_, _09129_);
  nor (_09133_, _09132_, _09045_);
  and (_09134_, _09133_, _09041_);
  or (_09135_, _09134_, _09039_);
  nor (_09136_, _09135_, _09035_);
  nor (_09137_, _09136_, _09032_);
  not (_09138_, _06154_);
  and (_09139_, _09138_, _02743_);
  nor (_09140_, _09138_, _02743_);
  nor (_09141_, _09140_, _09139_);
  and (_09142_, _09141_, _09137_);
  nor (_09143_, _09141_, _09137_);
  or (_09144_, _09143_, _09142_);
  and (_09145_, _05330_, _05328_);
  and (_09146_, _03989_, _03805_);
  and (_09147_, _09146_, _05207_);
  nand (_09148_, _09147_, _09145_);
  and (_09149_, _09148_, _09144_);
  and (_09150_, _09147_, _09145_);
  and (_09151_, _09150_, _06154_);
  or (_09152_, _09151_, _09149_);
  or (_09153_, _09152_, _05325_);
  and (_09154_, _08791_, _07428_);
  not (_09155_, _08791_);
  and (_09156_, _02777_, _02803_);
  not (_09157_, _09156_);
  and (_09158_, _07413_, _07408_);
  and (_09159_, _09158_, _09157_);
  nor (_09160_, _02971_, _02409_);
  or (_09161_, _09160_, _02545_);
  and (_09162_, _07431_, _02803_);
  nor (_09163_, _09162_, _07415_);
  and (_09164_, _09163_, _09161_);
  and (_09165_, _09164_, _09159_);
  nor (_09166_, _09165_, _09155_);
  not (_09167_, _02837_);
  and (_09168_, _09161_, _09167_);
  and (_09169_, _02546_, \oc8051_golden_model_1.PC [15]);
  and (_09170_, _09169_, _09163_);
  and (_09171_, _09170_, _09168_);
  and (_09172_, _09171_, _07429_);
  and (_09173_, _09172_, _09159_);
  or (_09174_, _09173_, _09166_);
  and (_09175_, _09174_, _07406_);
  or (_09176_, _09175_, _09154_);
  and (_09177_, _09176_, _02544_);
  and (_09178_, _02933_, _02564_);
  or (_09179_, _02837_, _02804_);
  or (_09180_, _09179_, _02934_);
  or (_09181_, _09180_, _09178_);
  nor (_09182_, _07425_, _09138_);
  and (_09183_, _09182_, _09181_);
  nand (_09184_, _08791_, _07425_);
  nand (_09185_, _09184_, _05325_);
  or (_09186_, _09185_, _09183_);
  or (_09187_, _09186_, _09177_);
  nor (_09188_, _03806_, _02932_);
  and (_09189_, _09188_, _09187_);
  and (_09190_, _09189_, _09153_);
  or (_09191_, _09190_, _09028_);
  and (_09192_, _09191_, _09018_);
  not (_09193_, _09015_);
  nand (_09194_, _09018_, _05311_);
  and (_09195_, _09194_, _08791_);
  or (_09196_, _09195_, _09193_);
  or (_09197_, _09196_, _09192_);
  and (_09198_, _09197_, _09016_);
  and (_09199_, _07475_, _03375_);
  not (_09200_, _09199_);
  or (_09201_, _09200_, _09198_);
  or (_09202_, _09199_, _08791_);
  and (_09203_, _09202_, _02943_);
  and (_09204_, _09203_, _09201_);
  and (_09205_, _06154_, _02928_);
  nor (_09206_, _07426_, _02537_);
  or (_09207_, _09206_, _09205_);
  or (_09208_, _09207_, _09204_);
  not (_09209_, _02538_);
  nor (_09210_, _02796_, _09209_);
  and (_09211_, _09210_, _03932_);
  not (_09212_, _09206_);
  or (_09213_, _09212_, _08791_);
  and (_09214_, _09213_, _09211_);
  and (_09215_, _09214_, _09208_);
  nor (_09216_, _03232_, _03001_);
  and (_09217_, _09216_, _03015_);
  or (_09218_, _09211_, _09138_);
  nand (_09219_, _09218_, _09217_);
  or (_09220_, _09219_, _09215_);
  and (_09221_, _04585_, _02858_);
  not (_09222_, _09221_);
  and (_09223_, _09222_, _04586_);
  nor (_09224_, _04735_, _04340_);
  and (_09225_, _04735_, _04340_);
  nor (_09226_, _09225_, _09224_);
  and (_09227_, _09226_, _09223_);
  and (_09228_, _04839_, _04621_);
  nor (_09229_, _04839_, _04621_);
  nor (_09230_, _09229_, _09228_);
  and (_09231_, _05143_, _04597_);
  nor (_09232_, _05143_, _04597_);
  nor (_09233_, _09232_, _09231_);
  and (_09234_, _09233_, _09230_);
  and (_09235_, _09234_, _09227_);
  and (_09236_, _04226_, _02774_);
  nor (_09237_, _04226_, _02774_);
  nor (_09238_, _09237_, _09236_);
  and (_09239_, _04413_, _03321_);
  nor (_09240_, _04413_, _03321_);
  nor (_09241_, _09240_, _09239_);
  and (_09242_, _09241_, _09238_);
  nor (_09243_, _03989_, _03743_);
  and (_09244_, _03805_, _02835_);
  and (_09245_, _03989_, _03743_);
  or (_09246_, _09245_, _09244_);
  nor (_09247_, _09246_, _09243_);
  and (_09248_, _09247_, _09242_);
  and (_09249_, _03823_, _02836_);
  not (_09250_, _09249_);
  and (_09251_, _09250_, _09248_);
  and (_09252_, _09251_, _09235_);
  or (_09253_, _09252_, _08964_);
  nand (_09254_, _09252_, _06146_);
  and (_09255_, _09254_, _09253_);
  or (_09256_, _09255_, _09217_);
  and (_09257_, _09256_, _02973_);
  and (_09258_, _09257_, _09220_);
  or (_09259_, _09258_, _09013_);
  or (_09260_, _09259_, _09004_);
  and (_09261_, _09260_, _08969_);
  or (_09262_, _09261_, _08968_);
  and (_09263_, _09262_, _08828_);
  nand (_09264_, _08827_, _08791_);
  nor (_09265_, _03842_, _04230_);
  and (_09266_, _09265_, _02926_);
  and (_09267_, _09266_, _02922_);
  nand (_09268_, _09267_, _09264_);
  or (_09269_, _09268_, _09263_);
  or (_09270_, _09267_, _06154_);
  and (_09271_, _02900_, _02523_);
  nor (_09272_, _09271_, _06195_);
  and (_09273_, _09272_, _08210_);
  and (_09274_, _09273_, _09270_);
  and (_09275_, _09274_, _09269_);
  not (_09276_, _02902_);
  not (_09277_, _02530_);
  nor (_09278_, _02901_, _09277_);
  and (_09279_, _09278_, _09276_);
  not (_09280_, _09279_);
  not (_09281_, _09273_);
  and (_09282_, _09281_, _08791_);
  or (_09283_, _09282_, _09280_);
  or (_09284_, _09283_, _09275_);
  and (_09285_, _07400_, _07330_);
  or (_09286_, _09279_, _06154_);
  and (_09287_, _09286_, _09285_);
  and (_09288_, _09287_, _09284_);
  nor (_09289_, _07540_, _02898_);
  not (_09290_, _09289_);
  nor (_09291_, _09285_, _09155_);
  or (_09292_, _09291_, _09290_);
  or (_09293_, _09292_, _09288_);
  or (_09294_, _09289_, _06154_);
  and (_09295_, _09294_, _02499_);
  and (_09296_, _09295_, _09293_);
  nand (_09297_, _08791_, _07700_);
  nor (_09298_, _02785_, _02518_);
  nand (_09299_, _09298_, _09297_);
  or (_09300_, _09299_, _09296_);
  or (_09301_, _09298_, _06154_);
  and (_09302_, _09301_, _08194_);
  and (_09303_, _09302_, _09300_);
  nand (_09304_, _06145_, _02975_);
  and (_09305_, _03860_, _06726_);
  nand (_09306_, _09305_, _09304_);
  or (_09307_, _09306_, _09303_);
  or (_09308_, _09305_, _06154_);
  and (_09309_, _09308_, _02970_);
  and (_09310_, _09309_, _09307_);
  and (_09311_, _06145_, _02524_);
  or (_09312_, _09311_, _08824_);
  or (_09313_, _09312_, _09310_);
  and (_09314_, _09313_, _08826_);
  nor (_09315_, _02894_, _02578_);
  not (_09316_, _09315_);
  or (_09317_, _09316_, _09314_);
  and (_09318_, _02777_, _02347_);
  not (_09319_, _09318_);
  or (_09320_, _09315_, _06154_);
  and (_09321_, _09320_, _09319_);
  and (_09322_, _09321_, _09317_);
  and (_09323_, _09318_, _09144_);
  or (_09324_, _09323_, _05516_);
  or (_09325_, _09324_, _09322_);
  or (_09326_, _06154_, _05267_);
  and (_09327_, _09326_, _09325_);
  or (_09328_, _09327_, _02974_);
  nand (_09329_, _06146_, _02974_);
  and (_09330_, _09329_, _07808_);
  and (_09331_, _09330_, _09328_);
  and (_09332_, _07807_, _06154_);
  or (_09333_, _09332_, _09331_);
  and (_09334_, _02584_, _02475_);
  not (_09335_, _09334_);
  and (_09336_, _09335_, _09333_);
  not (_09337_, \oc8051_golden_model_1.DPH [0]);
  and (_09338_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_09339_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor (_09340_, _09339_, _09338_);
  not (_09341_, _09340_);
  and (_09342_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_09343_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor (_09344_, _09343_, _09342_);
  and (_09345_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor (_09346_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  and (_09347_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_09348_, _02629_, _02625_);
  nor (_09349_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor (_09350_, _09349_, _09347_);
  not (_09351_, _09350_);
  nor (_09352_, _09351_, _09348_);
  nor (_09353_, _09352_, _09347_);
  nor (_09354_, _09353_, _09346_);
  or (_09355_, _09354_, _09345_);
  and (_09356_, _09355_, _09344_);
  nor (_09357_, _09356_, _09342_);
  nor (_09358_, _09357_, _09341_);
  nor (_09359_, _09358_, _09338_);
  nor (_09360_, _09359_, _09337_);
  and (_09361_, _09360_, \oc8051_golden_model_1.DPH [1]);
  and (_09362_, _09361_, \oc8051_golden_model_1.DPH [2]);
  and (_09363_, _09362_, \oc8051_golden_model_1.DPH [3]);
  and (_09364_, _09363_, \oc8051_golden_model_1.DPH [4]);
  and (_09365_, _09364_, \oc8051_golden_model_1.DPH [5]);
  and (_09366_, _09365_, \oc8051_golden_model_1.DPH [6]);
  or (_09367_, _09366_, \oc8051_golden_model_1.DPH [7]);
  nand (_09368_, _09366_, \oc8051_golden_model_1.DPH [7]);
  and (_09369_, _09368_, _09367_);
  and (_09370_, _09369_, _09334_);
  nor (_09371_, _02893_, _02585_);
  not (_09372_, _09371_);
  or (_09373_, _09372_, _09370_);
  or (_09374_, _09373_, _09336_);
  and (_09375_, _02777_, _02584_);
  not (_09376_, _09375_);
  or (_09377_, _09371_, _06154_);
  and (_09378_, _09377_, _09376_);
  and (_09379_, _09378_, _09374_);
  or (_09380_, _09144_, _08149_);
  not (_09381_, _08149_);
  or (_09382_, _09381_, _06154_);
  and (_09383_, _09382_, _09375_);
  and (_09384_, _09383_, _09380_);
  not (_09385_, _08822_);
  or (_09386_, _09385_, _09384_);
  or (_09387_, _09386_, _09379_);
  and (_09388_, _09387_, _08823_);
  or (_09389_, _09388_, _08815_);
  or (_09390_, _08814_, _06154_);
  and (_09391_, _09390_, _07092_);
  and (_09392_, _09391_, _09389_);
  nand (_09393_, _06145_, _02977_);
  nor (_09394_, _03107_, _02582_);
  nand (_09395_, _09394_, _09393_);
  or (_09396_, _09395_, _09392_);
  and (_09397_, _02777_, _02581_);
  not (_09398_, _09397_);
  or (_09399_, _09394_, _06154_);
  and (_09400_, _09399_, _09398_);
  and (_09401_, _09400_, _09396_);
  or (_09402_, _09144_, _09381_);
  or (_09403_, _08149_, _06154_);
  and (_09404_, _09403_, _09397_);
  and (_09405_, _09404_, _09402_);
  not (_09406_, _08812_);
  or (_09407_, _09406_, _09405_);
  or (_09408_, _09407_, _09401_);
  and (_09409_, _09408_, _08813_);
  or (_09410_, _09409_, _07882_);
  or (_09411_, _07881_, _06154_);
  and (_09412_, _09411_, _03881_);
  and (_09413_, _09412_, _09410_);
  nand (_09414_, _06145_, _02991_);
  nand (_09415_, _09414_, _08809_);
  or (_09416_, _09415_, _09413_);
  and (_09417_, _09416_, _08811_);
  not (_09418_, _08805_);
  or (_09419_, _09144_, \oc8051_golden_model_1.PSW [7]);
  or (_09420_, _06154_, _07294_);
  and (_09421_, _09420_, _08807_);
  and (_09422_, _09421_, _09419_);
  or (_09423_, _09422_, _09418_);
  or (_09424_, _09423_, _09417_);
  and (_09425_, _09424_, _08806_);
  or (_09426_, _09425_, _07901_);
  or (_09427_, _07900_, _06154_);
  and (_09428_, _09427_, _07120_);
  and (_09429_, _09428_, _09426_);
  nand (_09430_, _06145_, _02994_);
  nand (_09431_, _09430_, _08801_);
  or (_09432_, _09431_, _09429_);
  and (_09433_, _09432_, _08803_);
  not (_09434_, _08797_);
  or (_09435_, _09144_, _07294_);
  or (_09436_, _06154_, \oc8051_golden_model_1.PSW [7]);
  and (_09437_, _09436_, _08799_);
  and (_09438_, _09437_, _09435_);
  or (_09439_, _09438_, _09434_);
  or (_09440_, _09439_, _09433_);
  and (_09441_, _09440_, _08798_);
  or (_09442_, _09441_, _07948_);
  or (_09443_, _07947_, _06154_);
  and (_09444_, _09443_, _08028_);
  and (_09445_, _09444_, _09442_);
  and (_09446_, _08791_, _08027_);
  or (_09447_, _09446_, _03113_);
  or (_09448_, _09447_, _09445_);
  nand (_09449_, _04585_, _03113_);
  and (_09450_, _09449_, _09448_);
  or (_09451_, _09450_, _02592_);
  nand (_09452_, _09138_, _02592_);
  and (_09453_, _09452_, _03549_);
  and (_09454_, _09453_, _09451_);
  not (_09455_, _08795_);
  not (_09456_, _04669_);
  and (_09457_, _05275_, \oc8051_golden_model_1.TCON [2]);
  and (_09458_, _05291_, \oc8051_golden_model_1.ACC [2]);
  nor (_09459_, _09458_, _09457_);
  and (_09460_, _05289_, \oc8051_golden_model_1.PSW [2]);
  not (_09461_, _09460_);
  and (_09462_, _05284_, \oc8051_golden_model_1.IP [2]);
  and (_09463_, _05286_, \oc8051_golden_model_1.B [2]);
  nor (_09464_, _09463_, _09462_);
  and (_09465_, _09464_, _09461_);
  and (_09466_, _09465_, _09459_);
  and (_09467_, _05295_, \oc8051_golden_model_1.SCON [2]);
  and (_09468_, _05297_, \oc8051_golden_model_1.IE [2]);
  nor (_09469_, _09468_, _09467_);
  and (_09470_, _05300_, \oc8051_golden_model_1.P1INREG [2]);
  and (_09471_, _05280_, \oc8051_golden_model_1.P3INREG [2]);
  nor (_09472_, _09471_, _09470_);
  and (_09473_, _04613_, \oc8051_golden_model_1.P0INREG [2]);
  and (_09474_, _05278_, \oc8051_golden_model_1.P2INREG [2]);
  nor (_09475_, _09474_, _09473_);
  and (_09476_, _09475_, _09472_);
  and (_09477_, _09476_, _09469_);
  and (_09478_, _09477_, _09466_);
  and (_09479_, _09478_, _05038_);
  nor (_09480_, _09479_, _09456_);
  not (_09481_, _04595_);
  and (_09482_, _05275_, \oc8051_golden_model_1.TCON [1]);
  and (_09483_, _05291_, \oc8051_golden_model_1.ACC [1]);
  nor (_09484_, _09483_, _09482_);
  and (_09485_, _05289_, \oc8051_golden_model_1.PSW [1]);
  not (_09486_, _09485_);
  and (_09487_, _05284_, \oc8051_golden_model_1.IP [1]);
  and (_09488_, _05286_, \oc8051_golden_model_1.B [1]);
  nor (_09489_, _09488_, _09487_);
  and (_09490_, _09489_, _09486_);
  and (_09491_, _09490_, _09484_);
  and (_09492_, _05295_, \oc8051_golden_model_1.SCON [1]);
  and (_09493_, _05297_, \oc8051_golden_model_1.IE [1]);
  nor (_09494_, _09493_, _09492_);
  and (_09495_, _04613_, \oc8051_golden_model_1.P0INREG [1]);
  and (_09496_, _05278_, \oc8051_golden_model_1.P2INREG [1]);
  nor (_09497_, _09496_, _09495_);
  and (_09498_, _05300_, \oc8051_golden_model_1.P1INREG [1]);
  and (_09499_, _05280_, \oc8051_golden_model_1.P3INREG [1]);
  nor (_09500_, _09499_, _09498_);
  and (_09501_, _09500_, _09497_);
  and (_09502_, _09501_, _09494_);
  and (_09503_, _09502_, _09491_);
  and (_09504_, _09503_, _04940_);
  nor (_09505_, _09504_, _09481_);
  nor (_09506_, _09505_, _09480_);
  and (_09507_, _04603_, _03321_);
  not (_09508_, _09507_);
  and (_09509_, _05280_, \oc8051_golden_model_1.P3INREG [4]);
  and (_09510_, _05295_, \oc8051_golden_model_1.SCON [4]);
  and (_09511_, _05297_, \oc8051_golden_model_1.IE [4]);
  nor (_09512_, _09511_, _09510_);
  and (_09513_, _05289_, \oc8051_golden_model_1.PSW [4]);
  and (_09514_, _05286_, \oc8051_golden_model_1.B [4]);
  nor (_09515_, _09514_, _09513_);
  and (_09516_, _05284_, \oc8051_golden_model_1.IP [4]);
  and (_09517_, _05291_, \oc8051_golden_model_1.ACC [4]);
  nor (_09518_, _09517_, _09516_);
  and (_09519_, _09518_, _09515_);
  and (_09520_, _05278_, \oc8051_golden_model_1.P2INREG [4]);
  and (_09521_, _04613_, \oc8051_golden_model_1.P0INREG [4]);
  nor (_09522_, _09521_, _09520_);
  and (_09523_, _05275_, \oc8051_golden_model_1.TCON [4]);
  and (_09524_, _05300_, \oc8051_golden_model_1.P1INREG [4]);
  nor (_09525_, _09524_, _09523_);
  and (_09526_, _09525_, _09522_);
  and (_09527_, _09526_, _09519_);
  nand (_09528_, _09527_, _09512_);
  nor (_09529_, _09528_, _09509_);
  and (_09530_, _09529_, _05144_);
  nor (_09531_, _09530_, _09508_);
  nor (_09532_, _05499_, _05443_);
  nor (_09533_, _09532_, _09531_);
  and (_09534_, _09533_, _09506_);
  not (_09535_, _04607_);
  and (_09536_, _05284_, \oc8051_golden_model_1.IP [0]);
  and (_09537_, _05291_, \oc8051_golden_model_1.ACC [0]);
  nor (_09538_, _09537_, _09536_);
  and (_09539_, _05289_, \oc8051_golden_model_1.PSW [0]);
  and (_09540_, _05286_, \oc8051_golden_model_1.B [0]);
  nor (_09541_, _09540_, _09539_);
  and (_09542_, _09541_, _09538_);
  and (_09543_, _05295_, \oc8051_golden_model_1.SCON [0]);
  and (_09544_, _05297_, \oc8051_golden_model_1.IE [0]);
  nor (_09545_, _09544_, _09543_);
  and (_09546_, _05275_, \oc8051_golden_model_1.TCON [0]);
  and (_09547_, _05280_, \oc8051_golden_model_1.P3INREG [0]);
  nor (_09548_, _09547_, _09546_);
  and (_09549_, _09548_, _09545_);
  and (_09550_, _05300_, \oc8051_golden_model_1.P1INREG [0]);
  not (_09551_, _09550_);
  and (_09552_, _04613_, \oc8051_golden_model_1.P0INREG [0]);
  and (_09553_, _05278_, \oc8051_golden_model_1.P2INREG [0]);
  nor (_09554_, _09553_, _09552_);
  and (_09555_, _09554_, _09551_);
  and (_09556_, _09555_, _09549_);
  and (_09557_, _09556_, _09542_);
  and (_09558_, _09557_, _04989_);
  nor (_09559_, _09558_, _09535_);
  and (_09560_, _04628_, _03321_);
  not (_09561_, _09560_);
  and (_09562_, _05275_, \oc8051_golden_model_1.TCON [6]);
  and (_09563_, _05291_, \oc8051_golden_model_1.ACC [6]);
  nor (_09564_, _09563_, _09562_);
  and (_09565_, _05289_, \oc8051_golden_model_1.PSW [6]);
  not (_09566_, _09565_);
  and (_09567_, _05284_, \oc8051_golden_model_1.IP [6]);
  and (_09568_, _05286_, \oc8051_golden_model_1.B [6]);
  nor (_09569_, _09568_, _09567_);
  and (_09570_, _09569_, _09566_);
  and (_09571_, _09570_, _09564_);
  and (_09572_, _05295_, \oc8051_golden_model_1.SCON [6]);
  and (_09573_, _05297_, \oc8051_golden_model_1.IE [6]);
  nor (_09574_, _09573_, _09572_);
  and (_09575_, _04613_, \oc8051_golden_model_1.P0INREG [6]);
  and (_09576_, _05278_, \oc8051_golden_model_1.P2INREG [6]);
  nor (_09577_, _09576_, _09575_);
  and (_09578_, _05300_, \oc8051_golden_model_1.P1INREG [6]);
  and (_09579_, _05280_, \oc8051_golden_model_1.P3INREG [6]);
  nor (_09580_, _09579_, _09578_);
  and (_09581_, _09580_, _09577_);
  and (_09582_, _09581_, _09574_);
  and (_09583_, _09582_, _09571_);
  and (_09584_, _09583_, _04736_);
  nor (_09585_, _09584_, _09561_);
  nor (_09586_, _09585_, _09559_);
  not (_09587_, _04615_);
  and (_09588_, _05289_, \oc8051_golden_model_1.PSW [3]);
  and (_09589_, _05286_, \oc8051_golden_model_1.B [3]);
  nor (_09590_, _09589_, _09588_);
  and (_09591_, _05284_, \oc8051_golden_model_1.IP [3]);
  and (_09592_, _05291_, \oc8051_golden_model_1.ACC [3]);
  nor (_09593_, _09592_, _09591_);
  and (_09594_, _09593_, _09590_);
  and (_09595_, _04613_, \oc8051_golden_model_1.P0INREG [3]);
  not (_09596_, _09595_);
  and (_09597_, _05300_, \oc8051_golden_model_1.P1INREG [3]);
  and (_09598_, _05280_, \oc8051_golden_model_1.P3INREG [3]);
  nor (_09599_, _09598_, _09597_);
  and (_09600_, _09599_, _09596_);
  and (_09601_, _05295_, \oc8051_golden_model_1.SCON [3]);
  and (_09602_, _05297_, \oc8051_golden_model_1.IE [3]);
  nor (_09603_, _09602_, _09601_);
  and (_09604_, _05275_, \oc8051_golden_model_1.TCON [3]);
  and (_09605_, _05278_, \oc8051_golden_model_1.P2INREG [3]);
  nor (_09606_, _09605_, _09604_);
  and (_09607_, _09606_, _09603_);
  and (_09608_, _09607_, _09600_);
  and (_09609_, _09608_, _09594_);
  and (_09610_, _09609_, _04891_);
  nor (_09611_, _09610_, _09587_);
  and (_09612_, _04590_, _03321_);
  not (_09613_, _09612_);
  and (_09614_, _05295_, \oc8051_golden_model_1.SCON [5]);
  not (_09615_, _09614_);
  and (_09616_, _05275_, \oc8051_golden_model_1.TCON [5]);
  and (_09617_, _05297_, \oc8051_golden_model_1.IE [5]);
  nor (_09618_, _09617_, _09616_);
  and (_09619_, _09618_, _09615_);
  and (_09620_, _05284_, \oc8051_golden_model_1.IP [5]);
  and (_09621_, _05286_, \oc8051_golden_model_1.B [5]);
  nor (_09622_, _09621_, _09620_);
  and (_09623_, _05289_, \oc8051_golden_model_1.PSW [5]);
  and (_09624_, _05291_, \oc8051_golden_model_1.ACC [5]);
  nor (_09625_, _09624_, _09623_);
  and (_09626_, _09625_, _09622_);
  and (_09627_, _04613_, \oc8051_golden_model_1.P0INREG [5]);
  and (_09628_, _05278_, \oc8051_golden_model_1.P2INREG [5]);
  nor (_09629_, _09628_, _09627_);
  and (_09630_, _05300_, \oc8051_golden_model_1.P1INREG [5]);
  and (_09631_, _05280_, \oc8051_golden_model_1.P3INREG [5]);
  nor (_09632_, _09631_, _09630_);
  and (_09633_, _09632_, _09629_);
  and (_09634_, _09633_, _09626_);
  and (_09635_, _09634_, _09619_);
  and (_09636_, _09635_, _04840_);
  nor (_09637_, _09636_, _09613_);
  nor (_09638_, _09637_, _09611_);
  and (_09639_, _09638_, _09586_);
  and (_09640_, _09639_, _09534_);
  not (_09641_, _09640_);
  or (_09642_, _09641_, _08964_);
  or (_09643_, _09640_, _06145_);
  and (_09644_, _09643_, _02993_);
  and (_09645_, _09644_, _09642_);
  or (_09646_, _09645_, _09455_);
  or (_09647_, _09646_, _09454_);
  and (_09648_, _09647_, _08796_);
  or (_09649_, _09648_, _08772_);
  not (_09650_, _07143_);
  nand (_09651_, _08772_, _09138_);
  and (_09652_, _09651_, _09650_);
  and (_09653_, _09652_, _09649_);
  and (_09654_, _08791_, _07143_);
  or (_09655_, _09654_, _02854_);
  or (_09656_, _09655_, _09653_);
  nand (_09657_, _04585_, _02854_);
  and (_09658_, _09657_, _09656_);
  or (_09659_, _09658_, _02575_);
  nand (_09660_, _09138_, _02575_);
  and (_09661_, _09660_, _03134_);
  and (_09662_, _09661_, _09659_);
  or (_09663_, _09640_, _08964_);
  nand (_09664_, _09640_, _06146_);
  and (_09665_, _09664_, _09663_);
  and (_09666_, _09665_, _02990_);
  and (_09667_, _06085_, _05753_);
  not (_09668_, _09667_);
  or (_09669_, _09668_, _09666_);
  or (_09670_, _09669_, _09662_);
  or (_09671_, _09667_, _08791_);
  and (_09672_, _09671_, _03138_);
  and (_09673_, _09672_, _09670_);
  nand (_09674_, _06154_, _03133_);
  nor (_09675_, _08143_, _08138_);
  nand (_09676_, _09675_, _09674_);
  or (_09677_, _09676_, _09673_);
  or (_09678_, _09675_, _08791_);
  and (_09679_, _09678_, _05219_);
  and (_09680_, _09679_, _09677_);
  nor (_09681_, _05219_, _02743_);
  or (_09682_, _09681_, _02572_);
  or (_09683_, _09682_, _09680_);
  nand (_09684_, _09138_, _02572_);
  and (_09685_, _09684_, _03142_);
  and (_09686_, _09685_, _09683_);
  and (_09687_, _09665_, _02778_);
  and (_09688_, _05216_, _06112_);
  not (_09689_, _09688_);
  or (_09690_, _09689_, _09687_);
  or (_09691_, _09690_, _09686_);
  or (_09692_, _09688_, _08791_);
  and (_09693_, _09692_, _02853_);
  and (_09694_, _09693_, _09691_);
  nand (_09695_, _06154_, _02852_);
  nor (_09696_, _08167_, _08160_);
  nand (_09697_, _09696_, _09695_);
  or (_09698_, _09697_, _09694_);
  not (_09699_, _02982_);
  or (_09700_, _09696_, _08791_);
  and (_09701_, _09700_, _09699_);
  and (_09702_, _09701_, _09698_);
  nor (_09703_, _09699_, _02743_);
  or (_09704_, _09703_, _02568_);
  or (_09705_, _09704_, _09702_);
  and (_09706_, _02777_, _02567_);
  not (_09707_, _09706_);
  nand (_09708_, _09138_, _02568_);
  and (_09709_, _09708_, _09707_);
  and (_09710_, _09709_, _09705_);
  and (_09711_, _08791_, _09706_);
  or (_09712_, _09711_, _09710_);
  or (_09713_, _09712_, _34450_);
  or (_09714_, _34446_, \oc8051_golden_model_1.PC [15]);
  and (_09715_, _09714_, _35583_);
  and (_35629_[15], _09715_, _09713_);
  not (_09716_, _08143_);
  not (_09717_, _07844_);
  nor (_09718_, _08129_, _07843_);
  nor (_09719_, _09718_, _08074_);
  nand (_09720_, _09719_, _09717_);
  and (_09721_, _07702_, _04660_);
  and (_09722_, _07707_, \oc8051_golden_model_1.ACC [7]);
  nor (_09723_, _09722_, _08052_);
  not (_09724_, _09723_);
  or (_09725_, _09724_, _09721_);
  and (_09726_, _09725_, _07946_);
  and (_09727_, _07335_, \oc8051_golden_model_1.ACC [7]);
  or (_09728_, _09727_, _07940_);
  and (_09729_, _07332_, _05426_);
  or (_09730_, _09729_, _07917_);
  or (_09731_, _09730_, _09728_);
  not (_09732_, _03513_);
  and (_09733_, _07243_, _05208_);
  nor (_09734_, _07247_, _05719_);
  or (_09735_, _09734_, _07311_);
  or (_09736_, _09735_, _09733_);
  and (_09737_, _09736_, _09732_);
  or (_09738_, _09737_, _07241_);
  nor (_09739_, _04658_, _07294_);
  and (_09740_, _05722_, _04658_);
  or (_09741_, _09740_, _09739_);
  and (_09742_, _09741_, _03107_);
  and (_09743_, _05706_, _04658_);
  or (_09744_, _09743_, _09739_);
  and (_09745_, _09744_, _02524_);
  not (_09746_, _04658_);
  nor (_09747_, _09746_, _04585_);
  or (_09748_, _09747_, _09739_);
  or (_09749_, _09748_, _03860_);
  and (_09750_, _07343_, _07338_);
  nor (_09751_, _09750_, _07336_);
  not (_09752_, _09751_);
  and (_09753_, _07919_, _07338_);
  not (_09754_, _09753_);
  nor (_09755_, _09754_, _07391_);
  nor (_09756_, _09755_, _09752_);
  or (_09757_, _09729_, _07330_);
  or (_09758_, _09757_, _09756_);
  not (_09759_, _02901_);
  nor (_09760_, _09640_, _09276_);
  and (_09761_, _05278_, \oc8051_golden_model_1.P2 [2]);
  and (_09762_, _05280_, \oc8051_golden_model_1.P3 [2]);
  nor (_09763_, _09762_, _09761_);
  and (_09764_, _04613_, \oc8051_golden_model_1.P0 [2]);
  and (_09765_, _05300_, \oc8051_golden_model_1.P1 [2]);
  nor (_09766_, _09765_, _09764_);
  and (_09767_, _09766_, _09763_);
  and (_09768_, _09767_, _09469_);
  and (_09769_, _09768_, _09466_);
  and (_09770_, _09769_, _05038_);
  nor (_09771_, _09770_, _09456_);
  and (_09772_, _05278_, \oc8051_golden_model_1.P2 [1]);
  and (_09773_, _05280_, \oc8051_golden_model_1.P3 [1]);
  nor (_09774_, _09773_, _09772_);
  and (_09775_, _04613_, \oc8051_golden_model_1.P0 [1]);
  and (_09776_, _05300_, \oc8051_golden_model_1.P1 [1]);
  nor (_09777_, _09776_, _09775_);
  and (_09778_, _09777_, _09774_);
  and (_09779_, _09778_, _09494_);
  and (_09780_, _09779_, _09491_);
  and (_09781_, _09780_, _04940_);
  nor (_09782_, _09781_, _09481_);
  nor (_09783_, _09782_, _09771_);
  and (_09784_, _05280_, \oc8051_golden_model_1.P3 [4]);
  not (_09785_, _09784_);
  and (_09786_, _05278_, \oc8051_golden_model_1.P2 [4]);
  nor (_09787_, _09786_, _09523_);
  and (_09788_, _09787_, _09785_);
  and (_09789_, _04613_, \oc8051_golden_model_1.P0 [4]);
  and (_09790_, _05300_, \oc8051_golden_model_1.P1 [4]);
  nor (_09791_, _09790_, _09789_);
  and (_09792_, _09791_, _09512_);
  and (_09793_, _09792_, _09788_);
  and (_09794_, _09793_, _09519_);
  and (_09795_, _09794_, _05144_);
  nor (_09796_, _09508_, _09795_);
  nor (_09797_, _09796_, _05470_);
  and (_09798_, _09797_, _09783_);
  and (_09799_, _04613_, \oc8051_golden_model_1.P0 [0]);
  and (_09800_, _05300_, \oc8051_golden_model_1.P1 [0]);
  nor (_09801_, _09800_, _09799_);
  and (_09802_, _05280_, \oc8051_golden_model_1.P3 [0]);
  and (_09803_, _05278_, \oc8051_golden_model_1.P2 [0]);
  or (_09804_, _09803_, _09802_);
  nor (_09805_, _09804_, _09546_);
  and (_09806_, _09805_, _09542_);
  and (_09807_, _09806_, _09545_);
  and (_09808_, _09807_, _09801_);
  and (_09809_, _09808_, _04989_);
  nor (_09810_, _09809_, _09535_);
  and (_09811_, _05278_, \oc8051_golden_model_1.P2 [6]);
  and (_09812_, _05280_, \oc8051_golden_model_1.P3 [6]);
  nor (_09813_, _09812_, _09811_);
  and (_09814_, _04613_, \oc8051_golden_model_1.P0 [6]);
  and (_09815_, _05300_, \oc8051_golden_model_1.P1 [6]);
  nor (_09816_, _09815_, _09814_);
  and (_09817_, _09816_, _09813_);
  and (_09818_, _09817_, _09574_);
  and (_09819_, _09818_, _09571_);
  and (_09820_, _09819_, _04736_);
  nor (_09821_, _09561_, _09820_);
  nor (_09822_, _09821_, _09810_);
  and (_09823_, _05280_, \oc8051_golden_model_1.P3 [3]);
  not (_09824_, _09823_);
  and (_09825_, _05278_, \oc8051_golden_model_1.P2 [3]);
  nor (_09826_, _09825_, _09604_);
  and (_09827_, _09826_, _09824_);
  and (_09828_, _04613_, \oc8051_golden_model_1.P0 [3]);
  and (_09829_, _05300_, \oc8051_golden_model_1.P1 [3]);
  nor (_09830_, _09829_, _09828_);
  and (_09831_, _09830_, _09603_);
  and (_09832_, _09831_, _09827_);
  and (_09833_, _09832_, _09594_);
  and (_09834_, _09833_, _04891_);
  nor (_09835_, _09834_, _09587_);
  and (_09836_, _05278_, \oc8051_golden_model_1.P2 [5]);
  and (_09837_, _05280_, \oc8051_golden_model_1.P3 [5]);
  nor (_09838_, _09837_, _09836_);
  and (_09839_, _04613_, \oc8051_golden_model_1.P0 [5]);
  and (_09840_, _05300_, \oc8051_golden_model_1.P1 [5]);
  nor (_09841_, _09840_, _09839_);
  and (_09842_, _09841_, _09838_);
  and (_09843_, _09842_, _09626_);
  and (_09844_, _09843_, _09619_);
  and (_09845_, _09844_, _04840_);
  nor (_09846_, _09613_, _09845_);
  nor (_09847_, _09846_, _09835_);
  and (_09848_, _09847_, _09822_);
  and (_09849_, _09848_, _09798_);
  and (_09850_, _02925_, \oc8051_golden_model_1.PSW [7]);
  and (_09851_, _09850_, _09849_);
  nor (_09852_, _05289_, _07294_);
  and (_09853_, _05444_, _05289_);
  or (_09854_, _09853_, _09852_);
  or (_09855_, _09852_, _05471_);
  and (_09856_, _09855_, _02790_);
  and (_09857_, _09856_, _09854_);
  not (_09858_, _02972_);
  and (_09859_, _09217_, _09858_);
  and (_09860_, _09245_, _09242_);
  nor (_09861_, _09239_, _09236_);
  nor (_09862_, _09237_, _09861_);
  or (_09863_, _09862_, _09248_);
  or (_09864_, _09863_, _09860_);
  and (_09865_, _09864_, _09235_);
  or (_09866_, _09225_, _09221_);
  and (_09867_, _09866_, _04586_);
  nor (_09868_, _09231_, _09228_);
  nor (_09869_, _09229_, _09868_);
  and (_09870_, _09869_, _09227_);
  or (_09871_, _09870_, _09867_);
  or (_09872_, _09871_, _09865_);
  nor (_09873_, _09252_, _02972_);
  and (_09874_, _09873_, _09872_);
  or (_09875_, _09874_, _09859_);
  and (_09876_, _05439_, _04658_);
  nor (_09877_, _09876_, _09739_);
  nand (_09878_, _09877_, _02932_);
  not (_09879_, _07402_);
  and (_09880_, _04658_, \oc8051_golden_model_1.ACC [7]);
  or (_09881_, _09880_, _09739_);
  and (_09882_, _09881_, _02837_);
  nor (_09883_, _02837_, _07294_);
  or (_09884_, _09883_, _02932_);
  or (_09885_, _09884_, _09882_);
  and (_09886_, _09885_, _09879_);
  and (_09887_, _09886_, _09878_);
  nor (_09888_, _07444_, \oc8051_golden_model_1.PSW [7]);
  not (_09889_, _09888_);
  nor (_09890_, _09889_, _07454_);
  not (_09891_, _09890_);
  and (_09892_, _09891_, _02978_);
  or (_09893_, _09892_, _07431_);
  and (_09894_, _09893_, _02798_);
  or (_09895_, _09894_, _09887_);
  or (_09896_, _09854_, _03186_);
  and (_09897_, _09896_, _03693_);
  and (_09898_, _09897_, _09895_);
  and (_09899_, _09748_, _02930_);
  or (_09900_, _09899_, _02928_);
  or (_09901_, _09900_, _09898_);
  or (_09902_, _09881_, _02943_);
  nand (_09903_, _07431_, _02794_);
  and (_09904_, _09903_, _09902_);
  and (_09905_, _09904_, _09901_);
  not (_09906_, _09217_);
  and (_09907_, _05308_, _05289_);
  nor (_09908_, _09907_, _09852_);
  nor (_09909_, _09908_, _02927_);
  or (_09910_, _09909_, _09906_);
  or (_09911_, _09910_, _09905_);
  and (_09912_, _09911_, _09875_);
  and (_09913_, _08993_, _08991_);
  nand (_09914_, _08986_, _08988_);
  nand (_09915_, _09914_, _08985_);
  or (_09916_, _09915_, _08997_);
  or (_09917_, _09916_, _09913_);
  and (_09918_, _09917_, _08984_);
  nand (_09919_, _08977_, _08972_);
  nor (_09920_, _08982_, _09919_);
  nor (_09921_, _08976_, _05483_);
  or (_09922_, _09921_, _09920_);
  or (_09923_, _09922_, _09918_);
  nor (_09924_, _09000_, _09858_);
  and (_09925_, _09924_, _09923_);
  or (_09926_, _09925_, _09912_);
  nor (_09927_, _02979_, _02944_);
  and (_09928_, _09927_, _09926_);
  not (_09929_, _07682_);
  nor (_09930_, _07683_, _09929_);
  or (_09931_, _09930_, _07640_);
  and (_09932_, _09931_, _07681_);
  and (_09933_, _07680_, _07655_);
  or (_09934_, _09933_, _07613_);
  or (_09935_, _09934_, _09932_);
  and (_09936_, _09935_, _09007_);
  and (_09937_, _07674_, _07661_);
  or (_09938_, _09937_, _07574_);
  and (_09939_, _09938_, _09006_);
  nor (_09940_, _05466_, \oc8051_golden_model_1.ACC [7]);
  and (_09941_, _07558_, _07545_);
  or (_09942_, _09941_, _09940_);
  or (_09943_, _09942_, _09939_);
  or (_09944_, _09943_, _09936_);
  nor (_09945_, _09008_, _03397_);
  and (_09946_, _09945_, _09944_);
  or (_09947_, _02889_, \oc8051_golden_model_1.ACC [6]);
  nor (_09948_, _09947_, _07845_);
  nor (_09949_, _02743_, \oc8051_golden_model_1.ACC [7]);
  or (_09950_, _09949_, _09948_);
  nand (_09951_, _03179_, \oc8051_golden_model_1.ACC [5]);
  nor (_09952_, _03179_, \oc8051_golden_model_1.ACC [5]);
  nor (_09953_, _03620_, \oc8051_golden_model_1.ACC [4]);
  or (_09954_, _09953_, _09952_);
  and (_09955_, _09954_, _09951_);
  and (_09956_, _09955_, _08836_);
  or (_09957_, _09956_, _09950_);
  nor (_09958_, _03742_, \oc8051_golden_model_1.ACC [1]);
  and (_09959_, _03742_, \oc8051_golden_model_1.ACC [1]);
  and (_09960_, _02835_, \oc8051_golden_model_1.ACC [0]);
  nor (_09961_, _09960_, _09959_);
  or (_09962_, _09961_, _09958_);
  and (_09963_, _09962_, _08833_);
  or (_09964_, _02774_, _02605_);
  and (_09965_, _02774_, _02605_);
  nor (_09966_, _03320_, \oc8051_golden_model_1.ACC [2]);
  or (_09967_, _09966_, _09965_);
  and (_09968_, _09967_, _09964_);
  or (_09969_, _09968_, _09963_);
  and (_09970_, _09969_, _08837_);
  or (_09971_, _09970_, _09957_);
  nor (_09972_, _08839_, _08969_);
  and (_09973_, _09972_, _09971_);
  or (_09974_, _09973_, _08827_);
  or (_09975_, _09974_, _09946_);
  or (_09976_, _09975_, _09928_);
  and (_09977_, _08827_, \oc8051_golden_model_1.PSW [7]);
  nor (_09978_, _09977_, _02790_);
  and (_09979_, _09978_, _09976_);
  nor (_09980_, _09979_, _09857_);
  nor (_09981_, _09980_, _02925_);
  or (_09982_, _09981_, _09851_);
  nor (_09983_, _06195_, _02902_);
  and (_09984_, _09983_, _09982_);
  or (_09985_, _09984_, _09760_);
  and (_09986_, _09985_, _09759_);
  or (_09987_, _09849_, \oc8051_golden_model_1.PSW [7]);
  nand (_09988_, _09987_, _02901_);
  and (_09989_, _03009_, _02782_);
  nor (_09990_, _09989_, _07399_);
  nand (_09991_, _09990_, _09988_);
  or (_09992_, _09991_, _09986_);
  and (_09993_, _07255_, _07250_);
  nor (_09994_, _09993_, _07248_);
  not (_09995_, _09994_);
  and (_09996_, _07256_, _07250_);
  not (_09997_, _09996_);
  nor (_09998_, _09997_, _07529_);
  nor (_09999_, _09998_, _09995_);
  or (_10000_, _09999_, _09733_);
  nor (_10001_, _10000_, _09990_);
  nor (_10002_, _10001_, _03419_);
  and (_10003_, _10002_, _09992_);
  and (_10004_, _10000_, _03419_);
  or (_10005_, _10004_, _07329_);
  or (_10006_, _10005_, _10003_);
  and (_10007_, _10006_, _09758_);
  or (_10008_, _10007_, _02898_);
  and (_10009_, _07970_, _07965_);
  nor (_10010_, _10009_, _07963_);
  not (_10011_, _10010_);
  nor (_10012_, _07984_, _07979_);
  nor (_10013_, _10012_, _07978_);
  and (_10014_, _07986_, _07980_);
  and (_10015_, _07998_, _07992_);
  and (_10016_, _08006_, _02658_);
  nor (_10017_, _10016_, _08003_);
  or (_10018_, _10017_, _08002_);
  nand (_10019_, _10018_, _10015_);
  not (_10020_, _07990_);
  nand (_10021_, _07996_, _07992_);
  and (_10022_, _10021_, _10020_);
  and (_10023_, _10022_, _10019_);
  not (_10024_, _10023_);
  and (_10025_, _10024_, _10014_);
  nor (_10026_, _10025_, _10013_);
  and (_10027_, _07971_, _07965_);
  not (_10028_, _10027_);
  nor (_10029_, _10028_, _10026_);
  nor (_10030_, _10029_, _10011_);
  not (_10031_, _05466_);
  and (_10032_, _07959_, _10031_);
  or (_10033_, _10032_, _02899_);
  or (_10034_, _10033_, _10030_);
  and (_10035_, _10034_, _07541_);
  and (_10036_, _10035_, _10008_);
  and (_10037_, _07714_, _07710_);
  nor (_10038_, _10037_, _07708_);
  not (_10039_, _10038_);
  and (_10040_, _08031_, _07710_);
  not (_10041_, _10040_);
  nor (_10042_, _10041_, _07774_);
  nor (_10043_, _10042_, _10039_);
  or (_10044_, _10043_, _09721_);
  and (_10045_, _10044_, _07540_);
  or (_10046_, _10045_, _03861_);
  or (_10047_, _10046_, _10036_);
  and (_10048_, _10047_, _09749_);
  or (_10049_, _10048_, _03850_);
  and (_10050_, _05426_, _04658_);
  or (_10051_, _09739_, _06726_);
  or (_10052_, _10051_, _10050_);
  and (_10053_, _10052_, _02970_);
  and (_10054_, _10053_, _10049_);
  or (_10055_, _10054_, _09745_);
  nor (_10056_, _06731_, _02894_);
  and (_10057_, _10056_, _10055_);
  nor (_10058_, _09849_, _07294_);
  and (_10059_, _10058_, _02894_);
  or (_10060_, _10059_, _02974_);
  or (_10061_, _10060_, _10057_);
  and (_10062_, _05517_, _04658_);
  or (_10063_, _10062_, _09739_);
  or (_10064_, _10063_, _05261_);
  and (_10065_, _10064_, _10061_);
  or (_10066_, _10065_, _02893_);
  not (_10067_, _02893_);
  nand (_10068_, _09849_, _07294_);
  or (_10069_, _10068_, _10067_);
  and (_10070_, _10069_, _10066_);
  or (_10071_, _10070_, _02977_);
  and (_10072_, _05259_, _04658_);
  or (_10073_, _09739_, _07092_);
  or (_10074_, _10073_, _10072_);
  and (_10075_, _10074_, _07104_);
  and (_10076_, _10075_, _10071_);
  or (_10077_, _10076_, _09742_);
  and (_10078_, _10077_, _03095_);
  or (_10079_, _09739_, _04690_);
  and (_10080_, _09881_, _03094_);
  and (_10081_, _10063_, _02991_);
  or (_10082_, _10081_, _10080_);
  and (_10083_, _10082_, _10079_);
  or (_10084_, _10083_, _02994_);
  or (_10085_, _10084_, _10078_);
  nor (_10086_, _05257_, _09746_);
  or (_10087_, _10086_, _09739_);
  or (_10088_, _10087_, _07120_);
  and (_10089_, _10088_, _07118_);
  and (_10090_, _10089_, _10085_);
  nor (_10091_, _05721_, _09746_);
  or (_10092_, _10091_, _09739_);
  and (_10093_, _10092_, _03099_);
  nor (_10094_, _07239_, _02911_);
  nor (_10095_, _10094_, _07241_);
  or (_10096_, _10095_, _10093_);
  or (_10097_, _10096_, _10090_);
  and (_10098_, _10097_, _09738_);
  and (_10099_, _09736_, _03513_);
  or (_10100_, _10099_, _07236_);
  or (_10101_, _10100_, _10098_);
  and (_10102_, _10101_, _09731_);
  or (_10103_, _10102_, _03103_);
  nor (_10104_, _07962_, _05719_);
  or (_10105_, _10104_, _08021_);
  or (_10106_, _10105_, _10032_);
  or (_10107_, _10106_, _03104_);
  and (_10108_, _10107_, _08029_);
  and (_10109_, _10108_, _10103_);
  or (_10110_, _10109_, _09726_);
  and (_10111_, _10110_, _08028_);
  nand (_10112_, _08027_, \oc8051_golden_model_1.ACC [7]);
  nand (_10113_, _10112_, _07193_);
  or (_10114_, _10113_, _10111_);
  and (_10115_, _07229_, _07196_);
  nor (_10116_, _07197_, _07195_);
  nor (_10117_, _10116_, _07194_);
  or (_10118_, _10117_, _07193_);
  or (_10119_, _10118_, _10115_);
  and (_10120_, _10119_, _10114_);
  or (_10121_, _10120_, _07183_);
  and (_10122_, _07178_, _07147_);
  nor (_10123_, _07148_, _07146_);
  nor (_10124_, _10123_, _07145_);
  or (_10125_, _10124_, _08792_);
  or (_10126_, _10125_, _10122_);
  and (_10127_, _10126_, _02857_);
  and (_10128_, _10127_, _10121_);
  not (_10129_, _07542_);
  not (_10130_, _07543_);
  and (_10131_, _08096_, _10130_);
  nor (_10132_, _10131_, _03125_);
  and (_10133_, _10132_, _10129_);
  or (_10134_, _10133_, _08073_);
  or (_10135_, _10134_, _10128_);
  and (_10136_, _10135_, _09720_);
  and (_10137_, _10136_, _03138_);
  nor (_10138_, _09877_, _03138_);
  or (_10139_, _10138_, _10137_);
  and (_10140_, _10139_, _09716_);
  and (_10141_, _08143_, \oc8051_golden_model_1.ACC [0]);
  or (_10142_, _10141_, _10140_);
  and (_10143_, _10142_, _03142_);
  nor (_10144_, _09908_, _03142_);
  or (_10145_, _10144_, _10143_);
  nor (_10146_, _10145_, _02852_);
  and (_10147_, _05196_, _04658_);
  nor (_10148_, _10147_, _09739_);
  and (_10149_, _10148_, _02852_);
  nor (_10150_, _10149_, _10146_);
  or (_10151_, _10150_, _34450_);
  or (_10152_, _34446_, \oc8051_golden_model_1.PSW [7]);
  and (_10153_, _10152_, _35583_);
  and (_35630_[7], _10153_, _10151_);
  and (_35628_[7], \oc8051_golden_model_1.PCON [7], _35583_);
  and (_35631_[7], \oc8051_golden_model_1.SBUF [7], _35583_);
  and (_35632_[7], \oc8051_golden_model_1.SCON [7], _35583_);
  not (_10154_, \oc8051_golden_model_1.SP [7]);
  nor (_10155_, _04667_, _10154_);
  and (_10156_, _05196_, _04667_);
  nor (_10157_, _10156_, _10155_);
  nor (_10158_, _10157_, _02853_);
  not (_10159_, _03113_);
  not (_10160_, _08809_);
  and (_10161_, _05722_, _04667_);
  nor (_10162_, _10161_, _10155_);
  nor (_10163_, _10162_, _07104_);
  not (_10164_, _04667_);
  nor (_10165_, _10164_, _04585_);
  nor (_10166_, _10165_, _10155_);
  nor (_10167_, _10166_, _03860_);
  or (_10168_, _10167_, _03850_);
  nor (_10169_, _02837_, _10154_);
  and (_10170_, _04667_, \oc8051_golden_model_1.ACC [7]);
  nor (_10171_, _10170_, _10155_);
  nor (_10172_, _10171_, _09167_);
  or (_10173_, _10172_, _10169_);
  and (_10174_, _10173_, _02546_);
  and (_10175_, _04235_, \oc8051_golden_model_1.SP [4]);
  and (_10176_, _10175_, \oc8051_golden_model_1.SP [5]);
  and (_10177_, _10176_, \oc8051_golden_model_1.SP [6]);
  nor (_10178_, _10177_, \oc8051_golden_model_1.SP [7]);
  and (_10179_, _10177_, \oc8051_golden_model_1.SP [7]);
  nor (_10180_, _10179_, _10178_);
  and (_10181_, _10180_, _02804_);
  nor (_10182_, _10181_, _10174_);
  nor (_10183_, _10182_, _02932_);
  and (_10184_, _05439_, _04667_);
  nor (_10185_, _10184_, _10155_);
  nor (_10186_, _10185_, _06162_);
  or (_10187_, _10186_, _10183_);
  and (_10188_, _10187_, _02540_);
  not (_10189_, _10180_);
  nor (_10190_, _10189_, _02540_);
  or (_10191_, _10190_, _10188_);
  and (_10192_, _10191_, _03693_);
  not (_10193_, \oc8051_golden_model_1.SP [6]);
  not (_10194_, \oc8051_golden_model_1.SP [5]);
  not (_10195_, \oc8051_golden_model_1.SP [4]);
  and (_10196_, _05344_, _10195_);
  and (_10197_, _10196_, _10194_);
  and (_10198_, _10197_, _10193_);
  and (_10199_, _10198_, _02787_);
  nor (_10200_, _10199_, \oc8051_golden_model_1.SP [7]);
  and (_10201_, _10199_, \oc8051_golden_model_1.SP [7]);
  nor (_10202_, _10201_, _10200_);
  and (_10203_, _10202_, _10164_);
  nor (_10204_, _10203_, _10165_);
  nor (_10205_, _10204_, _03693_);
  or (_10206_, _10205_, _10192_);
  and (_10207_, _10206_, _02943_);
  nor (_10208_, _10171_, _02943_);
  or (_10209_, _10208_, _10207_);
  and (_10210_, _10209_, _03932_);
  not (_10211_, _04133_);
  and (_10212_, _10177_, \oc8051_golden_model_1.SP [0]);
  nor (_10213_, _10212_, _10154_);
  and (_10214_, _10212_, _10154_);
  nor (_10215_, _10214_, _10213_);
  nor (_10216_, _10215_, _03932_);
  nor (_10217_, _10216_, _10211_);
  not (_10218_, _10217_);
  nor (_10219_, _10218_, _10210_);
  nor (_10220_, _10180_, _04133_);
  or (_10221_, _10220_, _03861_);
  nor (_10222_, _10221_, _10219_);
  nor (_10223_, _10222_, _10168_);
  and (_10224_, _05426_, _04667_);
  nor (_10225_, _10155_, _06726_);
  not (_10226_, _10225_);
  nor (_10227_, _10226_, _10224_);
  or (_10228_, _10227_, _02524_);
  nor (_10229_, _10228_, _10223_);
  and (_10230_, _05706_, _04667_);
  nor (_10231_, _10230_, _10155_);
  nor (_10232_, _10231_, _02970_);
  or (_10233_, _10232_, _02974_);
  or (_10234_, _10233_, _10229_);
  and (_10235_, _05517_, _04667_);
  nor (_10236_, _10235_, _10155_);
  nand (_10237_, _10236_, _02974_);
  and (_10238_, _10237_, _10234_);
  nor (_10239_, _10238_, _02585_);
  and (_10240_, _10189_, _02585_);
  nor (_10241_, _10240_, _10239_);
  and (_10242_, _10241_, _07092_);
  and (_10243_, _05259_, _04667_);
  nor (_10244_, _10243_, _10155_);
  nor (_10245_, _10244_, _07092_);
  or (_10246_, _10245_, _10242_);
  and (_10247_, _10246_, _07104_);
  nor (_10248_, _10247_, _10163_);
  nor (_10249_, _10248_, _02991_);
  not (_10250_, _10155_);
  and (_10251_, _10250_, _04689_);
  or (_10252_, _10251_, _03881_);
  nor (_10253_, _10252_, _10236_);
  nor (_10254_, _10253_, _10249_);
  nor (_10255_, _10254_, _10160_);
  and (_10256_, _10180_, _02594_);
  nor (_10257_, _10256_, _02994_);
  or (_10258_, _10171_, _06161_);
  or (_10259_, _10258_, _10251_);
  nand (_10260_, _10259_, _10257_);
  nor (_10261_, _10260_, _10255_);
  nor (_10262_, _05257_, _10164_);
  or (_10263_, _10155_, _07120_);
  nor (_10264_, _10263_, _10262_);
  nor (_10265_, _10264_, _10261_);
  and (_10266_, _10265_, _07118_);
  nor (_10267_, _05721_, _10164_);
  nor (_10268_, _10267_, _10155_);
  nor (_10269_, _10268_, _07118_);
  or (_10270_, _10269_, _10266_);
  and (_10271_, _10270_, _10159_);
  nor (_10272_, _10198_, \oc8051_golden_model_1.SP [7]);
  and (_10273_, _10198_, \oc8051_golden_model_1.SP [7]);
  nor (_10274_, _10273_, _10272_);
  and (_10275_, _10274_, _03113_);
  or (_10276_, _10275_, _02592_);
  nor (_10277_, _10276_, _10271_);
  and (_10278_, _10189_, _02592_);
  nor (_10279_, _10278_, _10277_);
  and (_10280_, _10279_, _02855_);
  and (_10281_, _10274_, _02854_);
  or (_10282_, _10281_, _10280_);
  and (_10283_, _10282_, _03138_);
  nor (_10284_, _10185_, _03138_);
  or (_10285_, _10284_, _04331_);
  nor (_10286_, _10285_, _10283_);
  nor (_10287_, _10180_, _03907_);
  nor (_10288_, _10287_, _02852_);
  not (_10289_, _10288_);
  nor (_10290_, _10289_, _10286_);
  nor (_10291_, _10290_, _10158_);
  nand (_10292_, _10291_, _34446_);
  or (_10293_, _34446_, \oc8051_golden_model_1.SP [7]);
  and (_10294_, _10293_, _35583_);
  and (_35633_[7], _10294_, _10292_);
  and (_35634_[7], \oc8051_golden_model_1.TCON [7], _35583_);
  and (_35635_[7], \oc8051_golden_model_1.TH0 [7], _35583_);
  and (_35636_[7], \oc8051_golden_model_1.TH1 [7], _35583_);
  and (_35637_[7], \oc8051_golden_model_1.TL0 [7], _35583_);
  and (_35638_[7], \oc8051_golden_model_1.TL1 [7], _35583_);
  and (_35639_[7], \oc8051_golden_model_1.TMOD [7], _35583_);
  and (_10295_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [15]);
  not (_10296_, _03123_);
  and (_10297_, _07193_, _10296_);
  and (_10298_, _10297_, _03549_);
  and (_10299_, _09859_, _03932_);
  and (_10300_, _09199_, _03693_);
  and (_10301_, _09210_, _02943_);
  and (_10302_, _10301_, _09212_);
  and (_10303_, _10302_, _10300_);
  and (_10304_, _10303_, _10299_);
  and (_10305_, _09319_, _05267_);
  and (_10306_, _10305_, _10304_);
  and (_10307_, _09667_, _03134_);
  and (_10308_, _09305_, _08194_);
  nor (_10309_, _03113_, _02592_);
  nor (_10310_, _02982_, _02568_);
  and (_10311_, _10310_, _10309_);
  nor (_10312_, _03806_, _04087_);
  and (_10313_, _10312_, _10311_);
  nor (_10314_, _07807_, _02979_);
  nor (_10315_, _02974_, _02575_);
  nand (_10316_, _07431_, _02574_);
  and (_10317_, _10316_, _10315_);
  and (_10318_, _10317_, _10314_);
  nor (_10319_, _09290_, _03418_);
  and (_10320_, _10319_, _05324_);
  and (_10321_, _10320_, _10318_);
  and (_10322_, _10321_, _10313_);
  and (_10323_, _09014_, _06162_);
  and (_10324_, _10323_, _09018_);
  nor (_10325_, _08824_, _02524_);
  and (_10326_, _09315_, _10325_);
  and (_10327_, _10326_, _10324_);
  nor (_10328_, _09706_, _34450_);
  nor (_10329_, _08027_, _02944_);
  and (_10330_, _10329_, _10328_);
  and (_10331_, _09298_, _02499_);
  and (_10332_, _09371_, _09335_);
  and (_10333_, _10332_, _10331_);
  and (_10334_, _10333_, _10330_);
  and (_10335_, _10334_, _10327_);
  and (_10336_, _10335_, _10322_);
  and (_10337_, _10336_, _10308_);
  and (_10338_, _10337_, _10307_);
  and (_10339_, _10338_, _10306_);
  and (_10340_, _10339_, _10298_);
  and (_10341_, _09267_, _08828_);
  nor (_10342_, _02902_, _09277_);
  and (_10343_, _10342_, _09273_);
  and (_10344_, _10343_, _10341_);
  and (_10345_, _10344_, _09759_);
  and (_10346_, _02522_, _03003_);
  nand (_10347_, _10346_, _02782_);
  and (_10348_, _10347_, _07400_);
  and (_10349_, _10348_, _10345_);
  and (_10350_, _08822_, _09376_);
  and (_10351_, _10350_, _08814_);
  and (_10352_, _09394_, _07092_);
  not (_10353_, _02594_);
  and (_10354_, _03095_, _10353_);
  and (_10355_, _08812_, _09398_);
  and (_10356_, _10355_, _07881_);
  and (_10357_, _10356_, _10354_);
  and (_10358_, _10357_, _10352_);
  and (_10359_, _10358_, _10351_);
  and (_10360_, _10359_, _10349_);
  and (_10361_, _10360_, _10340_);
  or (_10362_, _09156_, _07425_);
  and (_10363_, _10362_, \oc8051_golden_model_1.DPH [7]);
  nor (_10364_, _09156_, _02804_);
  and (_10365_, _09163_, \oc8051_golden_model_1.XRAM_ADDR [15]);
  and (_10366_, _10365_, _09168_);
  and (_10367_, _10366_, _10364_);
  and (_10368_, _10367_, _02543_);
  or (_10369_, _10368_, _10363_);
  and (_10370_, _09688_, _03142_);
  and (_10371_, _09696_, _02853_);
  and (_10372_, _03907_, _03138_);
  and (_10373_, _09675_, _10372_);
  and (_10374_, _10373_, _10371_);
  and (_10375_, _10374_, _10370_);
  and (_10376_, _08800_, _08797_);
  and (_10377_, _10376_, _07947_);
  and (_10378_, _03100_, _02590_);
  and (_10379_, _08808_, _08805_);
  and (_10380_, _10379_, _07900_);
  and (_10381_, _10380_, _10378_);
  and (_10382_, _10381_, _10377_);
  and (_10383_, _10382_, _10375_);
  and (_10384_, _10383_, _10369_);
  and (_10385_, _10384_, _10361_);
  or (_10386_, _10385_, _10295_);
  and (_35640_[15], _10386_, _35583_);
  and (_10387_, _34450_, \oc8051_golden_model_1.XRAM_DATA_OUT [7]);
  nor (_10388_, _09162_, _09156_);
  nor (_10389_, _10388_, _05719_);
  and (_10390_, _10389_, _34446_);
  or (_10391_, _10390_, _10387_);
  and (_35642_[7], _10391_, _35583_);
  and (_10392_, _34450_, \oc8051_golden_model_1.P0INREG [7]);
  or (_10393_, _10392_, _00514_);
  and (_35620_[7], _10393_, _35583_);
  and (_10394_, _34450_, \oc8051_golden_model_1.P1INREG [7]);
  or (_10395_, _10394_, _00501_);
  and (_35622_[7], _10395_, _35583_);
  and (_10396_, _34450_, \oc8051_golden_model_1.P2INREG [7]);
  or (_10397_, _10396_, _00604_);
  and (_35624_[7], _10397_, _35583_);
  and (_10398_, _34450_, \oc8051_golden_model_1.P3INREG [7]);
  or (_10399_, _10398_, _00696_);
  and (_35626_[7], _10399_, _35583_);
  and (_35641_[7], \oc8051_golden_model_1.XRAM_DATA_IN [7], _35583_);
  nor (_10400_, _04348_, _04174_);
  nor (_10401_, _10400_, _04498_);
  nor (_10402_, _04174_, _03920_);
  nor (_10403_, _10402_, _04175_);
  and (_10404_, _10403_, _04173_);
  and (_10405_, _10404_, _10401_);
  or (_10406_, _10405_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor (_10407_, _04512_, _04080_);
  not (_10408_, _10407_);
  not (_10409_, _03925_);
  and (_10410_, _10407_, _04505_);
  and (_10411_, _10407_, _04508_);
  or (_10412_, _10411_, _10410_);
  or (_10413_, _10412_, _10409_);
  or (_10414_, _10413_, _10408_);
  and (_10415_, _10414_, _10406_);
  nor (_10416_, _04520_, _04079_);
  nor (_10417_, _10416_, _04521_);
  nor (_10418_, _04520_, _04497_);
  nor (_10419_, _10418_, _04525_);
  and (_10420_, _10419_, _04519_);
  nand (_10421_, _10420_, _10417_);
  nand (_10422_, _02572_, _02225_);
  nor (_10423_, _05036_, \oc8051_golden_model_1.ACC [0]);
  nand (_10424_, _10423_, _05736_);
  nor (_10425_, _05036_, _05647_);
  and (_10426_, _05036_, _05647_);
  nor (_10427_, _10426_, _10425_);
  and (_10428_, _10427_, _05225_);
  nor (_10429_, _09809_, _04607_);
  or (_10430_, _10429_, _05270_);
  and (_10431_, _05327_, _03823_);
  and (_10432_, _02804_, \oc8051_golden_model_1.PC [0]);
  and (_10433_, _02546_, \oc8051_golden_model_1.ACC [0]);
  or (_10434_, _10433_, _10432_);
  and (_10435_, _10434_, _05325_);
  or (_10436_, _10435_, _10431_);
  and (_10437_, _10436_, _03992_);
  nor (_10438_, _05036_, _03992_);
  or (_10439_, _10438_, _10437_);
  and (_10440_, _10439_, _05310_);
  nand (_10441_, _09809_, _09535_);
  and (_10442_, _10441_, _03810_);
  or (_10443_, _10442_, _04239_);
  or (_10444_, _10443_, _10440_);
  nor (_10445_, _02540_, \oc8051_golden_model_1.PC [0]);
  nor (_10446_, _10445_, _03818_);
  and (_10447_, _10446_, _10444_);
  and (_10448_, _03818_, _03805_);
  or (_10449_, _10448_, _03827_);
  or (_10450_, _10449_, _10447_);
  and (_10451_, _10450_, _10430_);
  or (_10452_, _10451_, _02795_);
  nand (_10453_, _07651_, _02795_);
  and (_10454_, _10453_, _02793_);
  and (_10455_, _10454_, _10452_);
  nor (_10456_, _09810_, _02793_);
  and (_10457_, _10456_, _10441_);
  or (_10458_, _10457_, _10455_);
  and (_10459_, _10458_, _02533_);
  or (_10460_, _02533_, _02225_);
  nand (_10461_, _02922_, _10460_);
  or (_10462_, _10461_, _10459_);
  nand (_10463_, _07651_, _02923_);
  and (_10464_, _10463_, _10462_);
  or (_10465_, _10464_, _03842_);
  or (_10466_, _05889_, _02858_);
  nand (_10467_, _10466_, _07650_);
  or (_10468_, _10467_, _05349_);
  and (_10469_, _10468_, _04289_);
  and (_10470_, _10469_, _10465_);
  nor (_10471_, _09558_, _04607_);
  and (_10472_, _04607_, \oc8051_golden_model_1.PSW [7]);
  nor (_10473_, _10472_, _10471_);
  nor (_10474_, _10473_, _04289_);
  or (_10475_, _10474_, _02518_);
  or (_10476_, _10475_, _10470_);
  and (_10477_, _02518_, _02225_);
  nor (_10478_, _10477_, _03862_);
  and (_10479_, _10478_, _10476_);
  and (_10480_, _03862_, _03805_);
  or (_10481_, _10480_, _03851_);
  or (_10482_, _10481_, _10479_);
  or (_10483_, _06114_, _03852_);
  and (_10484_, _10483_, _05512_);
  and (_10485_, _10484_, _10482_);
  and (_10486_, _05256_, _03805_);
  and (_10487_, _05619_, \oc8051_golden_model_1.TCON [0]);
  and (_10488_, _05635_, \oc8051_golden_model_1.ACC [0]);
  nor (_10489_, _10488_, _10487_);
  and (_10490_, _05631_, \oc8051_golden_model_1.PSW [0]);
  and (_10491_, _05626_, \oc8051_golden_model_1.B [0]);
  nor (_10492_, _10491_, _10490_);
  and (_10493_, _10492_, _10489_);
  and (_10494_, _05639_, \oc8051_golden_model_1.P0INREG [0]);
  and (_10495_, _05650_, \oc8051_golden_model_1.SBUF [0]);
  nor (_10496_, _10495_, _10494_);
  and (_10497_, _05645_, \oc8051_golden_model_1.P1INREG [0]);
  and (_10498_, _05642_, \oc8051_golden_model_1.SCON [0]);
  nor (_10499_, _10498_, _10497_);
  and (_10500_, _10499_, _10496_);
  and (_10501_, _05686_, \oc8051_golden_model_1.TH0 [0]);
  not (_10502_, _10501_);
  and (_10503_, _05665_, \oc8051_golden_model_1.P2INREG [0]);
  and (_10504_, _05659_, \oc8051_golden_model_1.IE [0]);
  nor (_10505_, _10504_, _10503_);
  and (_10506_, _05662_, \oc8051_golden_model_1.P3INREG [0]);
  and (_10507_, _05667_, \oc8051_golden_model_1.IP [0]);
  nor (_10508_, _10507_, _10506_);
  and (_10509_, _10508_, _10505_);
  and (_10510_, _10509_, _10502_);
  and (_10511_, _10510_, _10500_);
  and (_10512_, _10511_, _10493_);
  and (_10513_, _05681_, \oc8051_golden_model_1.DPH [0]);
  and (_10514_, _05695_, \oc8051_golden_model_1.TMOD [0]);
  nor (_10515_, _10514_, _10513_);
  and (_10516_, _05698_, \oc8051_golden_model_1.TL0 [0]);
  and (_10517_, _05700_, \oc8051_golden_model_1.TL1 [0]);
  nor (_10518_, _10517_, _10516_);
  and (_10519_, _10518_, _10515_);
  and (_10520_, _05684_, \oc8051_golden_model_1.SP [0]);
  and (_10521_, _05656_, \oc8051_golden_model_1.TH1 [0]);
  nor (_10522_, _10521_, _10520_);
  and (_10523_, _05677_, \oc8051_golden_model_1.DPL [0]);
  and (_10524_, _05692_, \oc8051_golden_model_1.PCON [0]);
  nor (_10525_, _10524_, _10523_);
  and (_10526_, _10525_, _10522_);
  and (_10527_, _10526_, _10519_);
  and (_10528_, _10527_, _10512_);
  not (_10529_, _10528_);
  nor (_10530_, _10529_, _10486_);
  nor (_10531_, _10530_, _05512_);
  or (_10532_, _10531_, _05516_);
  or (_10533_, _10532_, _10485_);
  and (_10534_, _05516_, _02835_);
  nor (_10535_, _10534_, _03874_);
  and (_10536_, _10535_, _10533_);
  and (_10537_, _03874_, _05647_);
  or (_10538_, _10537_, _02585_);
  or (_10539_, _10538_, _10536_);
  and (_10540_, _02585_, _02225_);
  nor (_10541_, _10540_, _05225_);
  and (_10542_, _10541_, _10539_);
  or (_10543_, _10542_, _10428_);
  and (_10544_, _10543_, _05224_);
  and (_10545_, _05036_, \oc8051_golden_model_1.ACC [0]);
  nor (_10546_, _10545_, _10423_);
  and (_10547_, _10546_, _05223_);
  or (_10548_, _10547_, _05221_);
  or (_10549_, _10548_, _10544_);
  or (_10550_, _10426_, _05222_);
  and (_10551_, _10550_, _05220_);
  and (_10552_, _10551_, _10549_);
  and (_10553_, _10545_, _03880_);
  or (_10554_, _10553_, _02594_);
  or (_10555_, _10554_, _10552_);
  and (_10556_, _02594_, _02225_);
  nor (_10557_, _10556_, _05732_);
  and (_10558_, _10557_, _10555_);
  nor (_10559_, _10425_, _05737_);
  or (_10560_, _10559_, _05736_);
  or (_10561_, _10560_, _10558_);
  and (_10562_, _10561_, _10424_);
  or (_10563_, _10562_, _02592_);
  nand (_10564_, _02592_, _02225_);
  and (_10565_, _10564_, _06085_);
  and (_10566_, _10565_, _10563_);
  nor (_10567_, _06085_, _03805_);
  or (_10568_, _10567_, _10566_);
  and (_10569_, _10568_, _05753_);
  and (_10570_, _05889_, _03898_);
  or (_10571_, _10570_, _03900_);
  or (_10572_, _10571_, _10569_);
  nand (_10573_, _05036_, _03900_);
  and (_10574_, _10573_, _05219_);
  and (_10575_, _10574_, _10572_);
  and (_10576_, _02988_, _02225_);
  or (_10577_, _10576_, _02572_);
  or (_10578_, _10577_, _10575_);
  and (_10579_, _10578_, _10422_);
  or (_10580_, _10579_, _02780_);
  or (_10581_, _10471_, _02781_);
  and (_10582_, _10581_, _05216_);
  and (_10583_, _10582_, _10580_);
  and (_10584_, _06105_, _03823_);
  or (_10585_, _10584_, _10583_);
  and (_10586_, _10585_, _06112_);
  and (_10587_, _05889_, _03912_);
  or (_10588_, _10587_, _03914_);
  or (_10589_, _10588_, _10586_);
  nand (_10590_, _05036_, _03914_);
  and (_10591_, _10590_, _04519_);
  and (_10592_, _10591_, _10589_);
  or (_10593_, _10592_, _10421_);
  and (_10594_, _10593_, _10415_);
  and (_10595_, _04513_, _04505_);
  nor (_10596_, _10595_, _04514_);
  and (_10597_, _04513_, _03925_);
  and (_10598_, _10597_, _10596_);
  nand (_10599_, _08936_, _02988_);
  or (_10600_, _09067_, _02988_);
  and (_10601_, _10600_, _10599_);
  and (_10602_, _10601_, _04513_);
  and (_10603_, _10602_, _10598_);
  or (_35643_, _10603_, _10594_);
  or (_10604_, _10405_, \oc8051_golden_model_1.IRAM[0] [1]);
  and (_10605_, _10604_, _10414_);
  nor (_10606_, _05329_, _05201_);
  and (_10607_, _10606_, _03581_);
  nor (_10608_, _04987_, _02477_);
  and (_10609_, _04987_, _02477_);
  nor (_10610_, _10609_, _10608_);
  and (_10611_, _10610_, _05223_);
  and (_10612_, _04987_, _03660_);
  nor (_10613_, _04987_, _03660_);
  nor (_10614_, _10613_, _10612_);
  and (_10615_, _10614_, _05225_);
  not (_10616_, _09782_);
  nand (_10617_, _09781_, _09481_);
  and (_10618_, _10617_, _02792_);
  and (_10619_, _10618_, _10616_);
  nor (_10620_, _09781_, _04595_);
  or (_10621_, _10620_, _05270_);
  nor (_10622_, _05432_, _05037_);
  nor (_10623_, _10622_, _03992_);
  nand (_10624_, _10606_, _05327_);
  and (_10625_, _02804_, _02198_);
  and (_10626_, _02546_, \oc8051_golden_model_1.ACC [1]);
  nor (_10627_, _10626_, _10625_);
  and (_10628_, _10627_, _05325_);
  nor (_10629_, _10628_, _03811_);
  and (_10630_, _10629_, _10624_);
  or (_10631_, _10630_, _03810_);
  or (_10632_, _10631_, _10623_);
  or (_10633_, _10617_, _05310_);
  and (_10634_, _10633_, _10632_);
  or (_10635_, _10634_, _04239_);
  nor (_10636_, _02540_, _02198_);
  nor (_10637_, _10636_, _03818_);
  and (_10638_, _10637_, _10635_);
  and (_10639_, _03990_, _03818_);
  or (_10640_, _10639_, _03827_);
  or (_10641_, _10640_, _10638_);
  and (_10642_, _10641_, _10621_);
  or (_10643_, _10642_, _02795_);
  nand (_10644_, _07638_, _02795_);
  and (_10645_, _10644_, _02793_);
  and (_10646_, _10645_, _10643_);
  or (_10647_, _10646_, _10619_);
  and (_10648_, _10647_, _02533_);
  or (_10649_, _02533_, \oc8051_golden_model_1.PC [1]);
  nand (_10650_, _02922_, _10649_);
  or (_10651_, _10650_, _10648_);
  nand (_10652_, _07638_, _02923_);
  and (_10653_, _10652_, _10651_);
  or (_10654_, _10653_, _03842_);
  and (_10655_, _06113_, _02743_);
  or (_10656_, _10655_, _07637_);
  or (_10657_, _10656_, _05349_);
  and (_10658_, _10657_, _04289_);
  and (_10659_, _10658_, _10654_);
  nor (_10660_, _09504_, _04595_);
  and (_10661_, _04595_, \oc8051_golden_model_1.PSW [7]);
  nor (_10662_, _10661_, _10660_);
  nor (_10663_, _10662_, _04289_);
  or (_10664_, _10663_, _02518_);
  or (_10665_, _10664_, _10659_);
  and (_10666_, _02518_, \oc8051_golden_model_1.PC [1]);
  nor (_10667_, _10666_, _03862_);
  and (_10668_, _10667_, _10665_);
  and (_10669_, _03990_, _03862_);
  or (_10670_, _10669_, _03851_);
  or (_10671_, _10670_, _10668_);
  or (_10672_, _06113_, _03852_);
  and (_10673_, _10672_, _05512_);
  and (_10674_, _10673_, _10671_);
  nor (_10675_, _05517_, _03989_);
  and (_10676_, _05619_, \oc8051_golden_model_1.TCON [1]);
  and (_10677_, _05635_, \oc8051_golden_model_1.ACC [1]);
  nor (_10678_, _10677_, _10676_);
  and (_10679_, _05631_, \oc8051_golden_model_1.PSW [1]);
  and (_10680_, _05626_, \oc8051_golden_model_1.B [1]);
  nor (_10681_, _10680_, _10679_);
  and (_10682_, _10681_, _10678_);
  and (_10683_, _05639_, \oc8051_golden_model_1.P0INREG [1]);
  and (_10684_, _05650_, \oc8051_golden_model_1.SBUF [1]);
  nor (_10685_, _10684_, _10683_);
  and (_10686_, _05645_, \oc8051_golden_model_1.P1INREG [1]);
  and (_10687_, _05642_, \oc8051_golden_model_1.SCON [1]);
  nor (_10688_, _10687_, _10686_);
  and (_10689_, _10688_, _10685_);
  and (_10690_, _05686_, \oc8051_golden_model_1.TH0 [1]);
  not (_10691_, _10690_);
  and (_10692_, _05665_, \oc8051_golden_model_1.P2INREG [1]);
  and (_10693_, _05659_, \oc8051_golden_model_1.IE [1]);
  nor (_10694_, _10693_, _10692_);
  and (_10695_, _05662_, \oc8051_golden_model_1.P3INREG [1]);
  and (_10696_, _05667_, \oc8051_golden_model_1.IP [1]);
  nor (_10697_, _10696_, _10695_);
  and (_10698_, _10697_, _10694_);
  and (_10699_, _10698_, _10691_);
  and (_10700_, _10699_, _10689_);
  and (_10701_, _10700_, _10682_);
  and (_10702_, _05681_, \oc8051_golden_model_1.DPH [1]);
  and (_10703_, _05695_, \oc8051_golden_model_1.TMOD [1]);
  nor (_10704_, _10703_, _10702_);
  and (_10705_, _05698_, \oc8051_golden_model_1.TL0 [1]);
  and (_10706_, _05700_, \oc8051_golden_model_1.TL1 [1]);
  nor (_10707_, _10706_, _10705_);
  and (_10708_, _10707_, _10704_);
  and (_10709_, _05684_, \oc8051_golden_model_1.SP [1]);
  and (_10710_, _05656_, \oc8051_golden_model_1.TH1 [1]);
  nor (_10711_, _10710_, _10709_);
  and (_10712_, _05677_, \oc8051_golden_model_1.DPL [1]);
  and (_10713_, _05692_, \oc8051_golden_model_1.PCON [1]);
  nor (_10714_, _10713_, _10712_);
  and (_10715_, _10714_, _10711_);
  and (_10716_, _10715_, _10708_);
  and (_10717_, _10716_, _10701_);
  not (_10718_, _10717_);
  nor (_10719_, _10718_, _10675_);
  nor (_10720_, _10719_, _05512_);
  or (_10721_, _10720_, _05516_);
  or (_10722_, _10721_, _10674_);
  and (_10723_, _05516_, _03742_);
  nor (_10724_, _10723_, _03874_);
  and (_10725_, _10724_, _10722_);
  and (_10726_, _03874_, _05675_);
  or (_10727_, _10726_, _02585_);
  or (_10728_, _10727_, _10725_);
  and (_10729_, _02585_, \oc8051_golden_model_1.PC [1]);
  nor (_10730_, _10729_, _05225_);
  and (_10731_, _10730_, _10728_);
  or (_10732_, _10731_, _10615_);
  and (_10733_, _10732_, _05224_);
  or (_10734_, _10733_, _10611_);
  and (_10735_, _10734_, _05222_);
  and (_10736_, _10613_, _05221_);
  or (_10737_, _10736_, _10735_);
  and (_10738_, _10737_, _05220_);
  and (_10739_, _10608_, _03880_);
  or (_10740_, _10739_, _02594_);
  or (_10741_, _10740_, _10738_);
  and (_10742_, _02594_, \oc8051_golden_model_1.PC [1]);
  nor (_10743_, _10742_, _05732_);
  and (_10744_, _10743_, _10741_);
  nor (_10745_, _10612_, _05737_);
  or (_10746_, _10745_, _05736_);
  or (_10747_, _10746_, _10744_);
  nand (_10748_, _10609_, _05736_);
  and (_10749_, _10748_, _05741_);
  and (_10750_, _10749_, _10747_);
  not (_10751_, _03236_);
  not (_10752_, _03229_);
  and (_10753_, _06083_, _10752_);
  and (_10754_, _10753_, _10751_);
  nand (_10755_, _02592_, _02198_);
  nand (_10756_, _03857_, _02571_);
  and (_10757_, _10756_, _10755_);
  nand (_10758_, _10757_, _10754_);
  or (_10759_, _10758_, _10750_);
  not (_10760_, _06085_);
  nand (_10761_, _10606_, _10760_);
  and (_10762_, _10761_, _05753_);
  and (_10763_, _10762_, _10759_);
  or (_10764_, _06115_, _05890_);
  and (_10765_, _10764_, _03898_);
  or (_10766_, _10765_, _10763_);
  and (_10767_, _10766_, _06080_);
  nor (_10768_, _10622_, _06080_);
  or (_10769_, _10768_, _02988_);
  or (_10770_, _10769_, _10767_);
  nand (_10771_, _02988_, _08909_);
  and (_10772_, _10771_, _05218_);
  and (_10773_, _10772_, _10770_);
  and (_10774_, _02572_, _02198_);
  or (_10775_, _02780_, _10774_);
  or (_10776_, _10775_, _10773_);
  nor (_10777_, _10660_, _02781_);
  and (_10778_, _03009_, _02567_);
  not (_10779_, _05215_);
  or (_10780_, _10779_, _10778_);
  nor (_10781_, _10780_, _10777_);
  and (_10782_, _10781_, _10776_);
  and (_10783_, _10780_, _10606_);
  nor (_10784_, _10783_, _10782_);
  nor (_10785_, _10784_, _03581_);
  or (_10786_, _10785_, _10607_);
  and (_10787_, _10786_, _06112_);
  nor (_10788_, _06115_, _05890_);
  and (_10789_, _10788_, _03912_);
  or (_10790_, _10789_, _03914_);
  or (_10791_, _10790_, _10787_);
  not (_10792_, _03914_);
  or (_10793_, _10622_, _10792_);
  and (_10794_, _10793_, _04519_);
  and (_10795_, _10794_, _10791_);
  or (_10796_, _10795_, _10421_);
  and (_10797_, _10796_, _10605_);
  nand (_10798_, _08874_, _02988_);
  or (_10799_, _09061_, _02988_);
  and (_10800_, _10799_, _10798_);
  and (_10801_, _10800_, _04513_);
  and (_10802_, _10801_, _10598_);
  or (_35644_, _10802_, _10797_);
  or (_10803_, _10405_, \oc8051_golden_model_1.IRAM[0] [2]);
  and (_10804_, _10803_, _10414_);
  nor (_10805_, _05201_, _04414_);
  nor (_10806_, _10805_, _07273_);
  and (_10807_, _10806_, _06105_);
  and (_10808_, _05890_, _05980_);
  nor (_10809_, _05890_, _05980_);
  or (_10810_, _10809_, _10808_);
  and (_10811_, _10810_, _03898_);
  nor (_10812_, _05085_, _03223_);
  and (_10813_, _10812_, _05221_);
  not (_10814_, _09771_);
  nand (_10815_, _09770_, _09456_);
  and (_10816_, _10815_, _02792_);
  and (_10817_, _10816_, _10814_);
  nor (_10818_, _09770_, _04669_);
  or (_10819_, _10818_, _05270_);
  or (_10820_, _10815_, _05310_);
  and (_10821_, _05085_, _04987_);
  and (_10822_, _10821_, _05431_);
  nor (_10823_, _05432_, _05085_);
  nor (_10824_, _10823_, _10822_);
  nor (_10825_, _10824_, _03992_);
  and (_10826_, _05329_, _04413_);
  nor (_10827_, _05329_, _04413_);
  or (_10828_, _10827_, _10826_);
  or (_10829_, _10828_, _05325_);
  and (_10830_, _02555_, _02804_);
  and (_10831_, _02546_, \oc8051_golden_model_1.ACC [2]);
  nor (_10832_, _10831_, _10830_);
  and (_10833_, _10832_, _05325_);
  nor (_10834_, _10833_, _03811_);
  and (_10835_, _10834_, _10829_);
  or (_10836_, _10835_, _03810_);
  or (_10837_, _10836_, _10825_);
  and (_10838_, _10837_, _10820_);
  or (_10839_, _10838_, _04239_);
  nor (_10840_, _02555_, _02540_);
  nor (_10841_, _10840_, _03818_);
  and (_10842_, _10841_, _10839_);
  and (_10843_, _04414_, _03818_);
  or (_10844_, _10843_, _03827_);
  or (_10845_, _10844_, _10842_);
  and (_10846_, _10845_, _10819_);
  or (_10847_, _10846_, _02795_);
  nand (_10848_, _07625_, _02795_);
  and (_10849_, _10848_, _02793_);
  and (_10850_, _10849_, _10847_);
  or (_10851_, _10850_, _10817_);
  and (_10852_, _10851_, _02533_);
  or (_10853_, _02600_, _02533_);
  nand (_10854_, _02922_, _10853_);
  or (_10855_, _10854_, _10852_);
  nand (_10856_, _07625_, _02923_);
  and (_10857_, _10856_, _10855_);
  or (_10858_, _10857_, _03842_);
  and (_10859_, _06117_, _02743_);
  or (_10860_, _10859_, _07624_);
  or (_10861_, _10860_, _05349_);
  and (_10862_, _10861_, _04289_);
  and (_10863_, _10862_, _10858_);
  nor (_10864_, _09479_, _04669_);
  and (_10865_, _04669_, \oc8051_golden_model_1.PSW [7]);
  nor (_10866_, _10865_, _10864_);
  nor (_10867_, _10866_, _04289_);
  or (_10868_, _10867_, _02518_);
  or (_10869_, _10868_, _10863_);
  and (_10870_, _02600_, _02518_);
  nor (_10871_, _10870_, _03862_);
  and (_10872_, _10871_, _10869_);
  and (_10873_, _04414_, _03862_);
  or (_10874_, _10873_, _03851_);
  or (_10875_, _10874_, _10872_);
  or (_10876_, _06117_, _03852_);
  and (_10877_, _10876_, _05512_);
  and (_10878_, _10877_, _10875_);
  nor (_10879_, _05517_, _04413_);
  not (_10880_, _10879_);
  and (_10881_, _05684_, \oc8051_golden_model_1.SP [2]);
  and (_10882_, _05639_, \oc8051_golden_model_1.P0INREG [2]);
  and (_10883_, _05677_, \oc8051_golden_model_1.DPL [2]);
  or (_10884_, _10883_, _10882_);
  nor (_10885_, _10884_, _10881_);
  and (_10886_, _05698_, \oc8051_golden_model_1.TL0 [2]);
  and (_10887_, _05700_, \oc8051_golden_model_1.TL1 [2]);
  and (_10888_, _05656_, \oc8051_golden_model_1.TH1 [2]);
  or (_10889_, _10888_, _10887_);
  nor (_10890_, _10889_, _10886_);
  and (_10891_, _10890_, _10885_);
  and (_10892_, _05659_, \oc8051_golden_model_1.IE [2]);
  and (_10893_, _05662_, \oc8051_golden_model_1.P3INREG [2]);
  and (_10894_, _05667_, \oc8051_golden_model_1.IP [2]);
  and (_10895_, _05631_, \oc8051_golden_model_1.PSW [2]);
  and (_10896_, _05626_, \oc8051_golden_model_1.B [2]);
  and (_10897_, _05635_, \oc8051_golden_model_1.ACC [2]);
  or (_10898_, _10897_, _10896_);
  or (_10899_, _10898_, _10895_);
  or (_10900_, _10899_, _10894_);
  or (_10901_, _10900_, _10893_);
  nor (_10902_, _10901_, _10892_);
  and (_10903_, _05686_, \oc8051_golden_model_1.TH0 [2]);
  and (_10904_, _05645_, \oc8051_golden_model_1.P1INREG [2]);
  and (_10905_, _05642_, \oc8051_golden_model_1.SCON [2]);
  and (_10906_, _05650_, \oc8051_golden_model_1.SBUF [2]);
  and (_10907_, _05665_, \oc8051_golden_model_1.P2INREG [2]);
  or (_10908_, _10907_, _10906_);
  or (_10909_, _10908_, _10905_);
  or (_10910_, _10909_, _10904_);
  nor (_10911_, _10910_, _10903_);
  and (_10912_, _05619_, \oc8051_golden_model_1.TCON [2]);
  and (_10913_, _05695_, \oc8051_golden_model_1.TMOD [2]);
  nor (_10914_, _10913_, _10912_);
  and (_10915_, _05681_, \oc8051_golden_model_1.DPH [2]);
  and (_10916_, _05692_, \oc8051_golden_model_1.PCON [2]);
  nor (_10917_, _10916_, _10915_);
  and (_10918_, _10917_, _10914_);
  and (_10919_, _10918_, _10911_);
  and (_10920_, _10919_, _10902_);
  and (_10921_, _10920_, _10891_);
  and (_10922_, _10921_, _10880_);
  nor (_10923_, _10922_, _05512_);
  or (_10924_, _10923_, _05516_);
  or (_10925_, _10924_, _10878_);
  and (_10926_, _05516_, _03320_);
  nor (_10927_, _10926_, _03874_);
  and (_10928_, _10927_, _10925_);
  and (_10929_, _03874_, _05690_);
  or (_10930_, _10929_, _02585_);
  or (_10931_, _10930_, _10928_);
  and (_10932_, _02585_, _02600_);
  nor (_10933_, _10932_, _05225_);
  and (_10934_, _10933_, _10931_);
  and (_10935_, _05085_, _03223_);
  nor (_10936_, _10935_, _10812_);
  and (_10937_, _10936_, _05225_);
  or (_10938_, _10937_, _05223_);
  or (_10939_, _10938_, _10934_);
  nor (_10940_, _05085_, _06908_);
  and (_10941_, _05085_, _06908_);
  nor (_10942_, _10941_, _10940_);
  or (_10943_, _10942_, _05224_);
  and (_10944_, _10943_, _05222_);
  and (_10945_, _10944_, _10939_);
  or (_10946_, _10945_, _10813_);
  and (_10947_, _10946_, _05220_);
  and (_10948_, _10940_, _03880_);
  or (_10949_, _10948_, _02594_);
  or (_10950_, _10949_, _10947_);
  and (_10951_, _02594_, _02600_);
  nor (_10952_, _10951_, _05732_);
  and (_10953_, _10952_, _10950_);
  nor (_10954_, _10935_, _05737_);
  or (_10955_, _10954_, _05736_);
  or (_10956_, _10955_, _10953_);
  nand (_10957_, _10941_, _05736_);
  and (_10958_, _10957_, _05741_);
  and (_10959_, _10958_, _10956_);
  nand (_10960_, _02592_, _02555_);
  nand (_10961_, _06085_, _10960_);
  or (_10962_, _10961_, _10959_);
  or (_10963_, _10828_, _06085_);
  and (_10964_, _10963_, _05753_);
  and (_10965_, _10964_, _10962_);
  or (_10966_, _10965_, _10811_);
  and (_10967_, _10966_, _06080_);
  nor (_10968_, _10824_, _06080_);
  or (_10969_, _10968_, _02988_);
  or (_10970_, _10969_, _10967_);
  nand (_10971_, _08907_, _02988_);
  and (_10972_, _10971_, _05218_);
  and (_10973_, _10972_, _10970_);
  and (_10974_, _02572_, _02555_);
  or (_10975_, _02780_, _10974_);
  or (_10976_, _10975_, _10973_);
  or (_10977_, _10864_, _02781_);
  and (_10978_, _10977_, _05216_);
  and (_10979_, _10978_, _10976_);
  or (_10980_, _10979_, _10807_);
  and (_10981_, _10980_, _06112_);
  or (_10982_, _06115_, _06117_);
  nor (_10983_, _07362_, _06112_);
  and (_10984_, _10983_, _10982_);
  or (_10985_, _10984_, _03914_);
  or (_10986_, _10985_, _10981_);
  nor (_10987_, _05086_, _05037_);
  nor (_10988_, _10987_, _05087_);
  or (_10989_, _10988_, _10792_);
  and (_10990_, _10989_, _04519_);
  and (_10991_, _10990_, _10986_);
  or (_10992_, _10991_, _10421_);
  and (_10993_, _10992_, _10804_);
  nand (_10994_, _08866_, _02988_);
  or (_10995_, _09054_, _02988_);
  and (_10996_, _10995_, _10994_);
  and (_10997_, _10996_, _04513_);
  and (_10998_, _10997_, _10598_);
  or (_35645_, _10998_, _10993_);
  or (_10999_, _10405_, \oc8051_golden_model_1.IRAM[0] [3]);
  and (_11000_, _10999_, _10414_);
  or (_11001_, _07273_, _07272_);
  nor (_11002_, _05216_, _05203_);
  and (_11003_, _11002_, _11001_);
  nor (_11004_, _10808_, _05935_);
  or (_11005_, _11004_, _05982_);
  and (_11006_, _11005_, _03898_);
  nor (_11007_, _04938_, _03087_);
  and (_11008_, _11007_, _05221_);
  nor (_11009_, _09834_, _04615_);
  or (_11010_, _11009_, _05270_);
  nand (_11011_, _09834_, _09587_);
  or (_11012_, _11011_, _05310_);
  nor (_11013_, _10822_, _04938_);
  nor (_11014_, _11013_, _05434_);
  nor (_11015_, _11014_, _03992_);
  nor (_11016_, _10826_, _04226_);
  or (_11017_, _11016_, _05331_);
  or (_11018_, _11017_, _05325_);
  and (_11019_, _02620_, _02804_);
  and (_11020_, _02546_, \oc8051_golden_model_1.ACC [3]);
  nor (_11021_, _11020_, _11019_);
  and (_11022_, _11021_, _05325_);
  nor (_11023_, _11022_, _03811_);
  and (_11024_, _11023_, _11018_);
  or (_11025_, _11024_, _03810_);
  or (_11026_, _11025_, _11015_);
  and (_11027_, _11026_, _11012_);
  or (_11028_, _11027_, _04239_);
  nor (_11029_, _02620_, _02540_);
  nor (_11030_, _11029_, _03818_);
  and (_11031_, _11030_, _11028_);
  and (_11032_, _07272_, _03818_);
  or (_11033_, _11032_, _03827_);
  or (_11034_, _11033_, _11031_);
  and (_11035_, _11034_, _11010_);
  or (_11036_, _11035_, _02795_);
  nand (_11037_, _07611_, _02795_);
  and (_11038_, _11037_, _02793_);
  and (_11039_, _11038_, _11036_);
  not (_11040_, _09835_);
  and (_11041_, _11011_, _11040_);
  and (_11042_, _11041_, _02792_);
  or (_11043_, _11042_, _11039_);
  and (_11044_, _11043_, _02533_);
  or (_11045_, _02641_, _02533_);
  nand (_11046_, _02922_, _11045_);
  or (_11047_, _11046_, _11044_);
  nand (_11048_, _07611_, _02923_);
  and (_11049_, _11048_, _11047_);
  or (_11050_, _11049_, _03842_);
  or (_11051_, _05935_, _02858_);
  nand (_11052_, _11051_, _07610_);
  or (_11053_, _11052_, _05349_);
  and (_11054_, _11053_, _04289_);
  and (_11055_, _11054_, _11050_);
  and (_11056_, _04615_, \oc8051_golden_model_1.PSW [7]);
  nor (_11057_, _09610_, _04615_);
  nor (_11058_, _11057_, _11056_);
  nor (_11059_, _11058_, _04289_);
  or (_11060_, _11059_, _02518_);
  or (_11061_, _11060_, _11055_);
  and (_11062_, _02641_, _02518_);
  nor (_11063_, _11062_, _03862_);
  and (_11064_, _11063_, _11061_);
  and (_11065_, _07272_, _03862_);
  or (_11066_, _11065_, _03851_);
  or (_11067_, _11066_, _11064_);
  or (_11068_, _06116_, _03852_);
  and (_11069_, _11068_, _05512_);
  and (_11070_, _11069_, _11067_);
  nor (_11071_, _05517_, _04226_);
  not (_11072_, _11071_);
  and (_11073_, _05692_, \oc8051_golden_model_1.PCON [3]);
  and (_11074_, _05684_, \oc8051_golden_model_1.SP [3]);
  and (_11075_, _05639_, \oc8051_golden_model_1.P0INREG [3]);
  and (_11076_, _05677_, \oc8051_golden_model_1.DPL [3]);
  or (_11077_, _11076_, _11075_);
  or (_11078_, _11077_, _11074_);
  nor (_11079_, _11078_, _11073_);
  and (_11080_, _05698_, \oc8051_golden_model_1.TL0 [3]);
  and (_11081_, _05700_, \oc8051_golden_model_1.TL1 [3]);
  and (_11082_, _05656_, \oc8051_golden_model_1.TH1 [3]);
  or (_11083_, _11082_, _11081_);
  nor (_11084_, _11083_, _11080_);
  and (_11085_, _05686_, \oc8051_golden_model_1.TH0 [3]);
  and (_11086_, _05645_, \oc8051_golden_model_1.P1INREG [3]);
  and (_11087_, _05642_, \oc8051_golden_model_1.SCON [3]);
  and (_11088_, _05650_, \oc8051_golden_model_1.SBUF [3]);
  and (_11089_, _05665_, \oc8051_golden_model_1.P2INREG [3]);
  or (_11090_, _11089_, _11088_);
  or (_11091_, _11090_, _11087_);
  or (_11092_, _11091_, _11086_);
  nor (_11093_, _11092_, _11085_);
  and (_11094_, _11093_, _11084_);
  and (_11095_, _05659_, \oc8051_golden_model_1.IE [3]);
  and (_11096_, _05662_, \oc8051_golden_model_1.P3INREG [3]);
  and (_11097_, _05667_, \oc8051_golden_model_1.IP [3]);
  and (_11098_, _05631_, \oc8051_golden_model_1.PSW [3]);
  and (_11099_, _05626_, \oc8051_golden_model_1.B [3]);
  and (_11100_, _05635_, \oc8051_golden_model_1.ACC [3]);
  or (_11101_, _11100_, _11099_);
  or (_11102_, _11101_, _11098_);
  or (_11103_, _11102_, _11097_);
  or (_11104_, _11103_, _11096_);
  nor (_11105_, _11104_, _11095_);
  and (_11106_, _05681_, \oc8051_golden_model_1.DPH [3]);
  and (_11107_, _05619_, \oc8051_golden_model_1.TCON [3]);
  and (_11108_, _05695_, \oc8051_golden_model_1.TMOD [3]);
  or (_11109_, _11108_, _11107_);
  nor (_11110_, _11109_, _11106_);
  and (_11111_, _11110_, _11105_);
  and (_11112_, _11111_, _11094_);
  and (_11113_, _11112_, _11079_);
  and (_11114_, _11113_, _11072_);
  nor (_11115_, _11114_, _05512_);
  or (_11116_, _11115_, _05516_);
  or (_11117_, _11116_, _11070_);
  nor (_11118_, _05267_, _02774_);
  nor (_11119_, _11118_, _03874_);
  and (_11120_, _11119_, _11117_);
  and (_11121_, _03874_, _05616_);
  or (_11122_, _11121_, _02585_);
  or (_11123_, _11122_, _11120_);
  and (_11124_, _02641_, _02585_);
  nor (_11125_, _11124_, _05225_);
  and (_11126_, _11125_, _11123_);
  and (_11127_, _04938_, _03087_);
  nor (_11128_, _11127_, _11007_);
  and (_11129_, _11128_, _05225_);
  or (_11130_, _11129_, _05223_);
  or (_11131_, _11130_, _11126_);
  nor (_11132_, _04938_, _02605_);
  and (_11133_, _04938_, _02605_);
  nor (_11134_, _11133_, _11132_);
  or (_11135_, _11134_, _05224_);
  and (_11136_, _11135_, _05222_);
  and (_11137_, _11136_, _11131_);
  or (_11138_, _11137_, _11008_);
  and (_11139_, _11138_, _05220_);
  and (_11140_, _11132_, _03880_);
  or (_11141_, _11140_, _02594_);
  or (_11142_, _11141_, _11139_);
  and (_11143_, _02641_, _02594_);
  nor (_11144_, _11143_, _05732_);
  and (_11145_, _11144_, _11142_);
  nor (_11146_, _11127_, _05737_);
  or (_11147_, _11146_, _05736_);
  or (_11148_, _11147_, _11145_);
  nand (_11149_, _11133_, _05736_);
  and (_11150_, _11149_, _05741_);
  and (_11151_, _11150_, _11148_);
  and (_11152_, _02620_, _02592_);
  or (_11153_, _06084_, _11152_);
  or (_11154_, _11153_, _11151_);
  not (_11155_, _03557_);
  and (_11156_, _11017_, _11155_);
  or (_11157_, _11156_, _06085_);
  and (_11158_, _11157_, _11154_);
  and (_11159_, _11017_, _03557_);
  or (_11160_, _11159_, _11158_);
  and (_11161_, _11160_, _05753_);
  or (_11162_, _11161_, _11006_);
  and (_11163_, _11162_, _06080_);
  nor (_11164_, _11014_, _06080_);
  or (_11165_, _11164_, _02988_);
  or (_11166_, _11165_, _11163_);
  nand (_11167_, _08902_, _02988_);
  and (_11168_, _11167_, _05218_);
  and (_11169_, _11168_, _11166_);
  and (_11170_, _02620_, _02572_);
  or (_11171_, _02780_, _11170_);
  or (_11172_, _11171_, _11169_);
  or (_11173_, _11057_, _02781_);
  and (_11174_, _11173_, _05216_);
  and (_11175_, _11174_, _11172_);
  or (_11176_, _11175_, _11003_);
  and (_11177_, _11176_, _06112_);
  or (_11178_, _07362_, _06116_);
  nor (_11179_, _06119_, _06112_);
  and (_11180_, _11179_, _11178_);
  or (_11181_, _11180_, _03914_);
  nor (_11182_, _11181_, _11177_);
  not (_11183_, _11182_);
  nor (_11184_, _05087_, _04939_);
  nor (_11185_, _11184_, _05088_);
  nor (_11186_, _11185_, _10792_);
  nor (_11187_, _11186_, _04520_);
  and (_11188_, _11187_, _11183_);
  or (_11189_, _11188_, _10421_);
  and (_11190_, _11189_, _11000_);
  nand (_11191_, _08859_, _02988_);
  or (_11192_, _09048_, _02988_);
  and (_11193_, _11192_, _11191_);
  and (_11194_, _11193_, _04513_);
  and (_11195_, _11194_, _10598_);
  or (_35646_, _11195_, _11190_);
  or (_11196_, _10405_, \oc8051_golden_model_1.IRAM[0] [4]);
  and (_11197_, _11196_, _10414_);
  nor (_11198_, _06119_, _06121_);
  nor (_11199_, _11198_, _07345_);
  or (_11200_, _11199_, _06112_);
  nor (_11201_, _05581_, _05189_);
  and (_11202_, _11201_, _05221_);
  nor (_11203_, _09507_, _09795_);
  or (_11204_, _11203_, _05270_);
  and (_11205_, _05434_, _05189_);
  nor (_11206_, _05434_, _05189_);
  nor (_11207_, _11206_, _11205_);
  nor (_11208_, _11207_, _03992_);
  or (_11209_, _06121_, _05311_);
  nor (_11210_, _05331_, _05143_);
  and (_11211_, _05331_, _05143_);
  or (_11212_, _11211_, _11210_);
  and (_11213_, _11212_, _05327_);
  and (_11214_, _09088_, _02804_);
  and (_11215_, _02546_, \oc8051_golden_model_1.ACC [4]);
  or (_11216_, _11215_, _11214_);
  and (_11217_, _11216_, _05325_);
  or (_11218_, _11217_, _03806_);
  or (_11219_, _11218_, _11213_);
  and (_11220_, _11219_, _03992_);
  and (_11221_, _11220_, _11209_);
  or (_11222_, _11221_, _11208_);
  and (_11223_, _11222_, _05310_);
  nand (_11224_, _09508_, _09795_);
  and (_11225_, _11224_, _03810_);
  or (_11226_, _11225_, _04239_);
  or (_11227_, _11226_, _11223_);
  nor (_11228_, _09088_, _02540_);
  nor (_11229_, _11228_, _03818_);
  and (_11230_, _11229_, _11227_);
  and (_11231_, _05200_, _03818_);
  or (_11232_, _11231_, _03827_);
  or (_11233_, _11232_, _11230_);
  and (_11234_, _11233_, _11204_);
  or (_11235_, _11234_, _02795_);
  nand (_11236_, _07593_, _02795_);
  and (_11237_, _11236_, _02793_);
  and (_11238_, _11237_, _11235_);
  not (_11239_, _09796_);
  and (_11240_, _11224_, _02792_);
  and (_11241_, _11240_, _11239_);
  or (_11242_, _11241_, _11238_);
  and (_11243_, _11242_, _02533_);
  or (_11244_, _09089_, _02533_);
  nand (_11245_, _11244_, _02922_);
  or (_11246_, _11245_, _11243_);
  nand (_11247_, _07593_, _02923_);
  and (_11248_, _11247_, _11246_);
  or (_11249_, _11248_, _03842_);
  and (_11250_, _06121_, _02743_);
  nand (_11251_, _07592_, _03842_);
  or (_11252_, _11251_, _11250_);
  and (_11253_, _11252_, _04289_);
  and (_11254_, _11253_, _11249_);
  nor (_11255_, _09530_, _09507_);
  and (_11256_, _09507_, \oc8051_golden_model_1.PSW [7]);
  nor (_11257_, _11256_, _11255_);
  nor (_11258_, _11257_, _04289_);
  or (_11259_, _11258_, _02518_);
  or (_11260_, _11259_, _11254_);
  and (_11261_, _09089_, _02518_);
  nor (_11262_, _11261_, _03862_);
  and (_11263_, _11262_, _11260_);
  and (_11264_, _05200_, _03862_);
  or (_11265_, _11264_, _03851_);
  or (_11266_, _11265_, _11263_);
  or (_11267_, _06121_, _03852_);
  and (_11268_, _11267_, _05512_);
  and (_11269_, _11268_, _11266_);
  nor (_11270_, _05517_, _05143_);
  not (_11271_, _11270_);
  and (_11272_, _05681_, \oc8051_golden_model_1.DPH [4]);
  and (_11273_, _05619_, \oc8051_golden_model_1.TCON [4]);
  and (_11274_, _05695_, \oc8051_golden_model_1.TMOD [4]);
  or (_11275_, _11274_, _11273_);
  nor (_11276_, _11275_, _11272_);
  and (_11277_, _05686_, \oc8051_golden_model_1.TH0 [4]);
  and (_11278_, _05656_, \oc8051_golden_model_1.TH1 [4]);
  and (_11279_, _05700_, \oc8051_golden_model_1.TL1 [4]);
  or (_11280_, _11279_, _11278_);
  nor (_11281_, _11280_, _11277_);
  and (_11282_, _11281_, _11276_);
  and (_11283_, _05659_, \oc8051_golden_model_1.IE [4]);
  and (_11284_, _05662_, \oc8051_golden_model_1.P3INREG [4]);
  and (_11285_, _05667_, \oc8051_golden_model_1.IP [4]);
  and (_11286_, _05631_, \oc8051_golden_model_1.PSW [4]);
  and (_11287_, _05635_, \oc8051_golden_model_1.ACC [4]);
  and (_11288_, _05626_, \oc8051_golden_model_1.B [4]);
  or (_11289_, _11288_, _11287_);
  or (_11290_, _11289_, _11286_);
  or (_11291_, _11290_, _11285_);
  or (_11292_, _11291_, _11284_);
  nor (_11293_, _11292_, _11283_);
  and (_11294_, _05698_, \oc8051_golden_model_1.TL0 [4]);
  and (_11295_, _05645_, \oc8051_golden_model_1.P1INREG [4]);
  and (_11296_, _05642_, \oc8051_golden_model_1.SCON [4]);
  and (_11297_, _05650_, \oc8051_golden_model_1.SBUF [4]);
  and (_11298_, _05665_, \oc8051_golden_model_1.P2INREG [4]);
  or (_11299_, _11298_, _11297_);
  or (_11300_, _11299_, _11296_);
  or (_11301_, _11300_, _11295_);
  nor (_11302_, _11301_, _11294_);
  and (_11303_, _05639_, \oc8051_golden_model_1.P0INREG [4]);
  and (_11304_, _05677_, \oc8051_golden_model_1.DPL [4]);
  nor (_11305_, _11304_, _11303_);
  and (_11306_, _05692_, \oc8051_golden_model_1.PCON [4]);
  and (_11307_, _05684_, \oc8051_golden_model_1.SP [4]);
  nor (_11308_, _11307_, _11306_);
  and (_11309_, _11308_, _11305_);
  and (_11310_, _11309_, _11302_);
  and (_11311_, _11310_, _11293_);
  and (_11312_, _11311_, _11282_);
  and (_11313_, _11312_, _11271_);
  nor (_11314_, _11313_, _05512_);
  or (_11315_, _11314_, _05516_);
  or (_11316_, _11315_, _11269_);
  and (_11317_, _05516_, _03620_);
  nor (_11318_, _11317_, _03874_);
  and (_11319_, _11318_, _11316_);
  and (_11320_, _05629_, _03874_);
  or (_11321_, _11320_, _02585_);
  or (_11322_, _11321_, _11319_);
  and (_11323_, _09089_, _02585_);
  nor (_11324_, _11323_, _05225_);
  and (_11325_, _11324_, _11322_);
  and (_11326_, _05581_, _05189_);
  nor (_11327_, _11326_, _11201_);
  and (_11328_, _11327_, _05225_);
  or (_11329_, _11328_, _05223_);
  or (_11330_, _11329_, _11325_);
  nor (_11331_, _05189_, _06814_);
  and (_11332_, _05189_, _06814_);
  nor (_11333_, _11332_, _11331_);
  or (_11334_, _11333_, _05224_);
  and (_11335_, _11334_, _05222_);
  and (_11336_, _11335_, _11330_);
  or (_11337_, _11336_, _11202_);
  and (_11338_, _11337_, _05220_);
  and (_11339_, _11331_, _03880_);
  or (_11340_, _11339_, _02594_);
  or (_11341_, _11340_, _11338_);
  and (_11342_, _09089_, _02594_);
  nor (_11343_, _11342_, _05732_);
  and (_11344_, _11343_, _11341_);
  nor (_11345_, _11326_, _05737_);
  or (_11346_, _11345_, _05736_);
  or (_11347_, _11346_, _11344_);
  nand (_11348_, _11332_, _05736_);
  and (_11349_, _11348_, _05741_);
  and (_11350_, _11349_, _11347_);
  nand (_11351_, _09088_, _02592_);
  nand (_11352_, _11351_, _06085_);
  or (_11353_, _11352_, _11350_);
  or (_11354_, _11212_, _06085_);
  and (_11355_, _11354_, _05753_);
  and (_11356_, _11355_, _11353_);
  and (_11357_, _05982_, _06072_);
  nor (_11358_, _05982_, _06072_);
  or (_11359_, _11358_, _11357_);
  and (_11360_, _11359_, _03898_);
  or (_11361_, _11360_, _11356_);
  and (_11362_, _11361_, _06080_);
  nor (_11363_, _11207_, _06080_);
  or (_11364_, _11363_, _02988_);
  or (_11365_, _11364_, _11362_);
  nand (_11366_, _08898_, _02988_);
  and (_11367_, _11366_, _05218_);
  and (_11368_, _11367_, _11365_);
  and (_11369_, _09088_, _02572_);
  or (_11370_, _11369_, _02780_);
  or (_11371_, _11370_, _11368_);
  or (_11372_, _11255_, _02781_);
  and (_11373_, _11372_, _05216_);
  and (_11374_, _11373_, _11371_);
  nor (_11375_, _05203_, _05200_);
  nor (_11376_, _11375_, _05204_);
  and (_11377_, _11376_, _06105_);
  or (_11378_, _11377_, _03912_);
  or (_11379_, _11378_, _11374_);
  and (_11380_, _11379_, _11200_);
  or (_11381_, _11380_, _03914_);
  nor (_11382_, _05190_, _05088_);
  nor (_11383_, _11382_, _05191_);
  or (_11384_, _11383_, _10792_);
  and (_11385_, _11384_, _04519_);
  and (_11386_, _11385_, _11381_);
  or (_11387_, _11386_, _10421_);
  and (_11388_, _11387_, _11197_);
  nand (_11389_, _08854_, _02988_);
  or (_11390_, _09043_, _02988_);
  and (_11391_, _11390_, _11389_);
  and (_11392_, _11391_, _04513_);
  and (_11393_, _11392_, _10598_);
  or (_35647_, _11393_, _11388_);
  or (_11394_, _10405_, \oc8051_golden_model_1.IRAM[0] [5]);
  and (_11395_, _11394_, _10414_);
  nor (_11396_, _11357_, _06027_);
  or (_11397_, _11396_, _06074_);
  and (_11398_, _11397_, _03898_);
  nor (_11399_, _11211_, _04839_);
  or (_11400_, _11399_, _05332_);
  and (_11401_, _11400_, _03557_);
  or (_11402_, _11400_, _06085_);
  nor (_11403_, _05612_, _04889_);
  and (_11404_, _11403_, _05221_);
  nor (_11405_, _09612_, _09845_);
  or (_11406_, _11405_, _05270_);
  nor (_11407_, _11205_, _04889_);
  nor (_11408_, _11407_, _05435_);
  nor (_11409_, _11408_, _03992_);
  or (_11410_, _06120_, _05311_);
  and (_11411_, _11400_, _05327_);
  and (_11412_, _02546_, \oc8051_golden_model_1.ACC [5]);
  and (_11413_, _09083_, _02804_);
  or (_11414_, _11413_, _11412_);
  and (_11415_, _11414_, _05325_);
  or (_11416_, _11415_, _03806_);
  or (_11417_, _11416_, _11411_);
  and (_11418_, _11417_, _03992_);
  and (_11419_, _11418_, _11410_);
  or (_11420_, _11419_, _11409_);
  and (_11421_, _11420_, _05310_);
  nand (_11422_, _09613_, _09845_);
  and (_11423_, _11422_, _03810_);
  or (_11424_, _11423_, _04239_);
  or (_11425_, _11424_, _11421_);
  nor (_11426_, _09083_, _02540_);
  nor (_11427_, _11426_, _03818_);
  and (_11428_, _11427_, _11425_);
  and (_11429_, _05199_, _03818_);
  or (_11430_, _11429_, _03827_);
  or (_11431_, _11430_, _11428_);
  and (_11432_, _11431_, _11406_);
  or (_11433_, _11432_, _02795_);
  nand (_11434_, _07572_, _02795_);
  and (_11435_, _11434_, _02793_);
  and (_11436_, _11435_, _11433_);
  not (_11437_, _09846_);
  and (_11438_, _11422_, _11437_);
  and (_11439_, _11438_, _02792_);
  or (_11440_, _11439_, _11436_);
  and (_11441_, _11440_, _02533_);
  or (_11442_, _09084_, _02533_);
  nand (_11443_, _11442_, _02922_);
  or (_11444_, _11443_, _11441_);
  nand (_11445_, _07572_, _02923_);
  and (_11446_, _11445_, _11444_);
  or (_11447_, _11446_, _03842_);
  and (_11448_, _06120_, _02743_);
  nand (_11449_, _07571_, _03842_);
  or (_11450_, _11449_, _11448_);
  and (_11451_, _11450_, _04289_);
  and (_11452_, _11451_, _11447_);
  nor (_11453_, _09636_, _09612_);
  and (_11454_, _09612_, \oc8051_golden_model_1.PSW [7]);
  nor (_11455_, _11454_, _11453_);
  nor (_11456_, _11455_, _04289_);
  or (_11457_, _11456_, _02518_);
  or (_11458_, _11457_, _11452_);
  and (_11459_, _09084_, _02518_);
  nor (_11460_, _11459_, _03862_);
  and (_11461_, _11460_, _11458_);
  and (_11462_, _05199_, _03862_);
  or (_11463_, _11462_, _03851_);
  or (_11464_, _11463_, _11461_);
  or (_11465_, _06120_, _03852_);
  and (_11466_, _11465_, _05512_);
  and (_11467_, _11466_, _11464_);
  nor (_11468_, _05517_, _04839_);
  not (_11469_, _11468_);
  and (_11470_, _05681_, \oc8051_golden_model_1.DPH [5]);
  and (_11471_, _05619_, \oc8051_golden_model_1.TCON [5]);
  and (_11472_, _05695_, \oc8051_golden_model_1.TMOD [5]);
  or (_11473_, _11472_, _11471_);
  nor (_11474_, _11473_, _11470_);
  and (_11475_, _05698_, \oc8051_golden_model_1.TL0 [5]);
  and (_11476_, _05700_, \oc8051_golden_model_1.TL1 [5]);
  and (_11477_, _05656_, \oc8051_golden_model_1.TH1 [5]);
  or (_11478_, _11477_, _11476_);
  nor (_11479_, _11478_, _11475_);
  and (_11480_, _11479_, _11474_);
  and (_11481_, _05659_, \oc8051_golden_model_1.IE [5]);
  and (_11482_, _05662_, \oc8051_golden_model_1.P3INREG [5]);
  and (_11483_, _05667_, \oc8051_golden_model_1.IP [5]);
  and (_11484_, _05631_, \oc8051_golden_model_1.PSW [5]);
  and (_11485_, _05626_, \oc8051_golden_model_1.B [5]);
  and (_11486_, _05635_, \oc8051_golden_model_1.ACC [5]);
  or (_11487_, _11486_, _11485_);
  or (_11488_, _11487_, _11484_);
  or (_11489_, _11488_, _11483_);
  or (_11490_, _11489_, _11482_);
  nor (_11491_, _11490_, _11481_);
  and (_11492_, _05686_, \oc8051_golden_model_1.TH0 [5]);
  and (_11493_, _05645_, \oc8051_golden_model_1.P1INREG [5]);
  and (_11494_, _05642_, \oc8051_golden_model_1.SCON [5]);
  and (_11495_, _05650_, \oc8051_golden_model_1.SBUF [5]);
  and (_11496_, _05665_, \oc8051_golden_model_1.P2INREG [5]);
  or (_11497_, _11496_, _11495_);
  or (_11498_, _11497_, _11494_);
  or (_11499_, _11498_, _11493_);
  nor (_11500_, _11499_, _11492_);
  and (_11501_, _05639_, \oc8051_golden_model_1.P0INREG [5]);
  and (_11502_, _05677_, \oc8051_golden_model_1.DPL [5]);
  nor (_11503_, _11502_, _11501_);
  and (_11504_, _05692_, \oc8051_golden_model_1.PCON [5]);
  and (_11505_, _05684_, \oc8051_golden_model_1.SP [5]);
  nor (_11506_, _11505_, _11504_);
  and (_11507_, _11506_, _11503_);
  and (_11508_, _11507_, _11500_);
  and (_11509_, _11508_, _11491_);
  and (_11510_, _11509_, _11480_);
  and (_11511_, _11510_, _11469_);
  nor (_11512_, _11511_, _05512_);
  or (_11513_, _11512_, _05516_);
  or (_11514_, _11513_, _11467_);
  and (_11515_, _05516_, _03179_);
  nor (_11516_, _11515_, _03874_);
  and (_11517_, _11516_, _11514_);
  and (_11518_, _05633_, _03874_);
  or (_11519_, _11518_, _02585_);
  or (_11520_, _11519_, _11517_);
  and (_11521_, _09084_, _02585_);
  nor (_11522_, _11521_, _05225_);
  and (_11523_, _11522_, _11520_);
  and (_11524_, _05612_, _04889_);
  nor (_11525_, _11524_, _11403_);
  and (_11526_, _11525_, _05225_);
  or (_11527_, _11526_, _05223_);
  or (_11528_, _11527_, _11523_);
  nor (_11529_, _04889_, _06808_);
  and (_11530_, _04889_, _06808_);
  nor (_11531_, _11530_, _11529_);
  or (_11532_, _11531_, _05224_);
  and (_11533_, _11532_, _05222_);
  and (_11534_, _11533_, _11528_);
  or (_11535_, _11534_, _11404_);
  and (_11536_, _11535_, _05220_);
  and (_11537_, _11529_, _03880_);
  or (_11538_, _11537_, _02594_);
  or (_11539_, _11538_, _11536_);
  and (_11540_, _09084_, _02594_);
  nor (_11541_, _11540_, _05732_);
  and (_11542_, _11541_, _11539_);
  nor (_11543_, _11524_, _05737_);
  or (_11544_, _11543_, _05736_);
  or (_11545_, _11544_, _11542_);
  nand (_11546_, _11530_, _05736_);
  and (_11547_, _11546_, _05741_);
  and (_11548_, _11547_, _11545_);
  and (_11549_, _09083_, _02592_);
  or (_11550_, _11549_, _06084_);
  or (_11551_, _11550_, _11548_);
  and (_11552_, _11551_, _11402_);
  or (_11553_, _11552_, _11401_);
  and (_11554_, _11553_, _05753_);
  or (_11555_, _11554_, _11398_);
  and (_11556_, _11555_, _06080_);
  nor (_11557_, _11408_, _06080_);
  or (_11558_, _11557_, _02988_);
  or (_11559_, _11558_, _11556_);
  nand (_11560_, _08893_, _02988_);
  and (_11561_, _11560_, _05218_);
  and (_11562_, _11561_, _11559_);
  and (_11563_, _09083_, _02572_);
  or (_11564_, _11563_, _02780_);
  or (_11565_, _11564_, _11562_);
  or (_11566_, _11453_, _02781_);
  and (_11567_, _11566_, _05216_);
  and (_11568_, _11567_, _11565_);
  nor (_11569_, _05204_, _05199_);
  nor (_11570_, _11569_, _05205_);
  and (_11571_, _11570_, _06105_);
  or (_11572_, _11571_, _11568_);
  and (_11573_, _11572_, _06112_);
  or (_11574_, _07345_, _06120_);
  nor (_11575_, _06123_, _06112_);
  and (_11576_, _11575_, _11574_);
  or (_11577_, _11576_, _03914_);
  or (_11578_, _11577_, _11573_);
  nor (_11579_, _05191_, _04890_);
  nor (_11580_, _11579_, _05192_);
  or (_11581_, _11580_, _10792_);
  and (_11582_, _11581_, _04519_);
  and (_11583_, _11582_, _11578_);
  or (_11584_, _11583_, _10421_);
  and (_11585_, _11584_, _11395_);
  nand (_11586_, _08849_, _02988_);
  or (_11587_, _09037_, _02988_);
  and (_11588_, _11587_, _11586_);
  and (_11589_, _11588_, _04513_);
  and (_11590_, _11589_, _10598_);
  or (_35648_, _11590_, _11585_);
  or (_11591_, _10405_, \oc8051_golden_model_1.IRAM[0] [6]);
  and (_11592_, _11591_, _10414_);
  nor (_11593_, _06123_, _05798_);
  nor (_11594_, _11593_, _06124_);
  or (_11595_, _11594_, _06112_);
  nor (_11596_, _06074_, _05799_);
  or (_11597_, _11596_, _06075_);
  and (_11598_, _11597_, _03898_);
  nor (_11599_, _04783_, _06762_);
  and (_11600_, _04783_, _06762_);
  nor (_11601_, _11600_, _11599_);
  and (_11602_, _11601_, _05223_);
  not (_11603_, _09821_);
  nand (_11604_, _09561_, _09820_);
  and (_11605_, _11604_, _11603_);
  and (_11606_, _11605_, _02792_);
  and (_11607_, _07242_, _03818_);
  or (_11608_, _11604_, _05310_);
  nor (_11609_, _05435_, _04783_);
  nor (_11610_, _11609_, _05436_);
  nor (_11611_, _11610_, _03992_);
  or (_11612_, _05798_, _05311_);
  nor (_11613_, _05332_, _04735_);
  or (_11614_, _11613_, _05333_);
  and (_11615_, _11614_, _05327_);
  and (_11616_, _09076_, _02804_);
  and (_11617_, _02546_, \oc8051_golden_model_1.ACC [6]);
  or (_11618_, _11617_, _11616_);
  and (_11619_, _11618_, _05325_);
  or (_11620_, _11619_, _03806_);
  or (_11621_, _11620_, _11615_);
  and (_11622_, _11621_, _03992_);
  and (_11623_, _11622_, _11612_);
  or (_11624_, _11623_, _11611_);
  or (_11625_, _11624_, _03810_);
  and (_11626_, _11625_, _11608_);
  or (_11627_, _11626_, _04239_);
  nor (_11628_, _09076_, _02540_);
  nor (_11629_, _11628_, _03818_);
  and (_11630_, _11629_, _11627_);
  or (_11631_, _11630_, _11607_);
  and (_11632_, _11631_, _05270_);
  nor (_11633_, _09560_, _09820_);
  and (_11634_, _11633_, _03827_);
  or (_11635_, _11634_, _02795_);
  or (_11636_, _11635_, _11632_);
  nand (_11637_, _07556_, _02795_);
  and (_11638_, _11637_, _02793_);
  and (_11639_, _11638_, _11636_);
  or (_11640_, _11639_, _11606_);
  and (_11641_, _11640_, _02533_);
  or (_11642_, _09077_, _02533_);
  nand (_11643_, _11642_, _02922_);
  or (_11644_, _11643_, _11641_);
  nand (_11645_, _07556_, _02923_);
  and (_11646_, _11645_, _11644_);
  or (_11647_, _11646_, _03842_);
  and (_11648_, _05798_, _02743_);
  nand (_11649_, _07555_, _03842_);
  or (_11650_, _11649_, _11648_);
  and (_11651_, _11650_, _04289_);
  and (_11652_, _11651_, _11647_);
  nor (_11653_, _09584_, _09560_);
  and (_11654_, _09560_, \oc8051_golden_model_1.PSW [7]);
  nor (_11655_, _11654_, _11653_);
  nor (_11656_, _11655_, _04289_);
  or (_11657_, _11656_, _02518_);
  or (_11658_, _11657_, _11652_);
  and (_11659_, _09077_, _02518_);
  nor (_11660_, _11659_, _03862_);
  and (_11661_, _11660_, _11658_);
  and (_11662_, _07242_, _03862_);
  or (_11663_, _11662_, _03851_);
  or (_11664_, _11663_, _11661_);
  or (_11665_, _05798_, _03852_);
  and (_11666_, _11665_, _05512_);
  and (_11667_, _11666_, _11664_);
  nor (_11668_, _05517_, _04735_);
  not (_11669_, _11668_);
  and (_11670_, _05692_, \oc8051_golden_model_1.PCON [6]);
  and (_11671_, _05619_, \oc8051_golden_model_1.TCON [6]);
  and (_11672_, _05695_, \oc8051_golden_model_1.TMOD [6]);
  or (_11673_, _11672_, _11671_);
  nor (_11674_, _11673_, _11670_);
  and (_11675_, _05698_, \oc8051_golden_model_1.TL0 [6]);
  and (_11676_, _05700_, \oc8051_golden_model_1.TL1 [6]);
  and (_11677_, _05656_, \oc8051_golden_model_1.TH1 [6]);
  or (_11678_, _11677_, _11676_);
  nor (_11679_, _11678_, _11675_);
  and (_11680_, _11679_, _11674_);
  and (_11681_, _05659_, \oc8051_golden_model_1.IE [6]);
  and (_11682_, _05662_, \oc8051_golden_model_1.P3INREG [6]);
  and (_11683_, _05667_, \oc8051_golden_model_1.IP [6]);
  and (_11684_, _05631_, \oc8051_golden_model_1.PSW [6]);
  and (_11685_, _05635_, \oc8051_golden_model_1.ACC [6]);
  and (_11686_, _05626_, \oc8051_golden_model_1.B [6]);
  or (_11687_, _11686_, _11685_);
  or (_11688_, _11687_, _11684_);
  or (_11689_, _11688_, _11683_);
  or (_11690_, _11689_, _11682_);
  nor (_11691_, _11690_, _11681_);
  and (_11692_, _05686_, \oc8051_golden_model_1.TH0 [6]);
  and (_11693_, _05642_, \oc8051_golden_model_1.SCON [6]);
  and (_11694_, _05645_, \oc8051_golden_model_1.P1INREG [6]);
  and (_11695_, _05650_, \oc8051_golden_model_1.SBUF [6]);
  and (_11696_, _05665_, \oc8051_golden_model_1.P2INREG [6]);
  or (_11697_, _11696_, _11695_);
  or (_11698_, _11697_, _11694_);
  or (_11699_, _11698_, _11693_);
  nor (_11700_, _11699_, _11692_);
  and (_11701_, _05639_, \oc8051_golden_model_1.P0INREG [6]);
  and (_11702_, _05677_, \oc8051_golden_model_1.DPL [6]);
  nor (_11703_, _11702_, _11701_);
  and (_11704_, _05681_, \oc8051_golden_model_1.DPH [6]);
  and (_11705_, _05684_, \oc8051_golden_model_1.SP [6]);
  nor (_11706_, _11705_, _11704_);
  and (_11707_, _11706_, _11703_);
  and (_11708_, _11707_, _11700_);
  and (_11709_, _11708_, _11691_);
  and (_11710_, _11709_, _11680_);
  and (_11711_, _11710_, _11669_);
  nor (_11712_, _11711_, _05512_);
  or (_11713_, _11712_, _05516_);
  or (_11714_, _11713_, _11667_);
  and (_11715_, _05516_, _02889_);
  nor (_11716_, _11715_, _03874_);
  and (_11717_, _11716_, _11714_);
  not (_11718_, _05549_);
  and (_11719_, _11718_, _03874_);
  or (_11720_, _11719_, _02585_);
  or (_11721_, _11720_, _11717_);
  nand (_11722_, _09077_, _02585_);
  and (_11723_, _11722_, _11721_);
  or (_11724_, _11723_, _05225_);
  not (_11725_, _05225_);
  and (_11726_, _05549_, _04783_);
  nor (_11727_, _05549_, _04783_);
  nor (_11728_, _11727_, _11726_);
  or (_11729_, _11728_, _11725_);
  and (_11730_, _11729_, _05224_);
  and (_11731_, _11730_, _11724_);
  or (_11732_, _11731_, _11602_);
  and (_11733_, _11732_, _05222_);
  and (_11734_, _11727_, _05221_);
  or (_11735_, _11734_, _11733_);
  and (_11736_, _11735_, _05220_);
  and (_11737_, _11599_, _03880_);
  or (_11738_, _11737_, _02594_);
  or (_11739_, _11738_, _11736_);
  and (_11740_, _09077_, _02594_);
  nor (_11741_, _11740_, _05732_);
  and (_11742_, _11741_, _11739_);
  nor (_11743_, _11726_, _05737_);
  or (_11744_, _11743_, _05736_);
  or (_11745_, _11744_, _11742_);
  nand (_11746_, _11600_, _05736_);
  and (_11747_, _11746_, _05741_);
  and (_11748_, _11747_, _11745_);
  nand (_11749_, _09076_, _02592_);
  nand (_11750_, _11749_, _06085_);
  or (_11751_, _11750_, _11748_);
  or (_11752_, _11614_, _06085_);
  and (_11753_, _11752_, _05753_);
  and (_11754_, _11753_, _11751_);
  or (_11755_, _11754_, _11598_);
  and (_11756_, _11755_, _06080_);
  nor (_11757_, _11610_, _06080_);
  or (_11758_, _11757_, _02988_);
  or (_11759_, _11758_, _11756_);
  nand (_11760_, _08886_, _02988_);
  and (_11761_, _11760_, _05218_);
  and (_11762_, _11761_, _11759_);
  and (_11763_, _09076_, _02572_);
  or (_11764_, _11763_, _02780_);
  or (_11765_, _11764_, _11762_);
  or (_11766_, _11653_, _02781_);
  and (_11767_, _11766_, _05216_);
  and (_11768_, _11767_, _11765_);
  nor (_11769_, _05205_, _04735_);
  and (_11770_, _05205_, _04735_);
  or (_11771_, _11770_, _11769_);
  and (_11772_, _11771_, _06105_);
  or (_11773_, _11772_, _03912_);
  or (_11774_, _11773_, _11768_);
  and (_11775_, _11774_, _11595_);
  or (_11776_, _11775_, _03914_);
  nor (_11777_, _05192_, _04784_);
  nor (_11778_, _11777_, _05193_);
  or (_11779_, _11778_, _10792_);
  and (_11780_, _11779_, _04519_);
  and (_11781_, _11780_, _11776_);
  or (_11782_, _11781_, _10421_);
  and (_11783_, _11782_, _11592_);
  nand (_11784_, _08842_, _02988_);
  or (_11785_, _09030_, _02988_);
  and (_11786_, _11785_, _11784_);
  and (_11787_, _11786_, _04513_);
  and (_11788_, _11787_, _10598_);
  or (_35649_, _11788_, _11783_);
  or (_11789_, _10405_, \oc8051_golden_model_1.IRAM[0] [7]);
  and (_11790_, _11789_, _10414_);
  nand (_11791_, _10405_, _06132_);
  and (_11792_, _11791_, _11790_);
  and (_11793_, _10598_, _06157_);
  or (_35650_, _11793_, _11792_);
  and (_11794_, _04521_, _04079_);
  and (_11795_, _11794_, _10419_);
  or (_11796_, _11795_, \oc8051_golden_model_1.IRAM[1] [0]);
  not (_11797_, _04231_);
  or (_11798_, _10412_, _11797_);
  or (_11799_, _11798_, _10408_);
  and (_11800_, _11799_, _11796_);
  not (_11801_, _11795_);
  or (_11802_, _11801_, _10592_);
  and (_11803_, _11802_, _11800_);
  and (_11804_, _04513_, _04231_);
  and (_11805_, _11804_, _10596_);
  and (_11806_, _11805_, _10602_);
  or (_35699_, _11806_, _11803_);
  or (_11807_, _11795_, \oc8051_golden_model_1.IRAM[1] [1]);
  and (_11808_, _11807_, _11799_);
  or (_11809_, _11801_, _10795_);
  and (_11810_, _11809_, _11808_);
  and (_11811_, _11805_, _10801_);
  or (_35700_, _11811_, _11810_);
  or (_11812_, _11795_, \oc8051_golden_model_1.IRAM[1] [2]);
  and (_11813_, _11812_, _11799_);
  or (_11814_, _11801_, _10991_);
  and (_11815_, _11814_, _11813_);
  and (_11816_, _11805_, _10997_);
  or (_35701_, _11816_, _11815_);
  or (_11817_, _11795_, \oc8051_golden_model_1.IRAM[1] [3]);
  and (_11818_, _11817_, _11799_);
  or (_11819_, _11801_, _11188_);
  and (_11820_, _11819_, _11818_);
  and (_11821_, _11805_, _11194_);
  or (_35702_, _11821_, _11820_);
  or (_11822_, _11795_, \oc8051_golden_model_1.IRAM[1] [4]);
  and (_11823_, _11822_, _11799_);
  or (_11824_, _11801_, _11386_);
  and (_11825_, _11824_, _11823_);
  and (_11826_, _11805_, _11392_);
  or (_35703_, _11826_, _11825_);
  or (_11827_, _11795_, \oc8051_golden_model_1.IRAM[1] [5]);
  and (_11828_, _11827_, _11799_);
  or (_11829_, _11801_, _11583_);
  and (_11830_, _11829_, _11828_);
  and (_11831_, _11805_, _11589_);
  or (_35704_, _11831_, _11830_);
  or (_11832_, _11795_, \oc8051_golden_model_1.IRAM[1] [6]);
  and (_11833_, _11832_, _11799_);
  or (_11834_, _11801_, _11781_);
  and (_11835_, _11834_, _11833_);
  and (_11836_, _11805_, _11787_);
  or (_35705_, _11836_, _11835_);
  or (_11837_, _11795_, \oc8051_golden_model_1.IRAM[1] [7]);
  and (_11838_, _11837_, _11799_);
  or (_11839_, _11801_, _06133_);
  and (_11840_, _11839_, _11838_);
  and (_11841_, _11805_, _06157_);
  or (_35706_, _11841_, _11840_);
  and (_11842_, _04175_, _03920_);
  and (_11843_, _11842_, _10401_);
  or (_11844_, _11843_, \oc8051_golden_model_1.IRAM[2] [0]);
  not (_11845_, _05340_);
  or (_11846_, _10412_, _11845_);
  or (_11847_, _11846_, _10408_);
  and (_11848_, _11847_, _11844_);
  and (_11849_, _10590_, _04173_);
  and (_11850_, _11849_, _10589_);
  not (_11851_, _11843_);
  or (_11852_, _11851_, _11850_);
  and (_11853_, _11852_, _11848_);
  and (_11854_, _05340_, _04513_);
  and (_11855_, _11854_, _10596_);
  and (_11856_, _11855_, _10602_);
  or (_35707_, _11856_, _11853_);
  or (_11857_, _11843_, \oc8051_golden_model_1.IRAM[2] [1]);
  and (_11858_, _11857_, _11847_);
  and (_11859_, _10793_, _04173_);
  and (_11860_, _11859_, _10791_);
  or (_11861_, _11851_, _11860_);
  and (_11862_, _11861_, _11858_);
  and (_11863_, _11855_, _10801_);
  or (_35708_, _11863_, _11862_);
  or (_11864_, _11843_, \oc8051_golden_model_1.IRAM[2] [2]);
  and (_11865_, _11864_, _11847_);
  and (_11866_, _10989_, _04173_);
  and (_11867_, _11866_, _10986_);
  or (_11868_, _11851_, _11867_);
  and (_11869_, _11868_, _11865_);
  and (_11870_, _11855_, _10997_);
  or (_35709_, _11870_, _11869_);
  or (_11871_, _11843_, \oc8051_golden_model_1.IRAM[2] [3]);
  and (_11872_, _11871_, _11847_);
  and (_11873_, _10416_, _03920_);
  nand (_11874_, _11873_, _10419_);
  or (_11875_, _11874_, _11188_);
  and (_11876_, _11875_, _11872_);
  and (_11877_, _11855_, _11194_);
  or (_35710_, _11877_, _11876_);
  or (_11878_, _11874_, _11386_);
  or (_11879_, _11843_, \oc8051_golden_model_1.IRAM[2] [4]);
  and (_11880_, _11879_, _11847_);
  and (_11881_, _11880_, _11878_);
  and (_11882_, _11855_, _11392_);
  or (_35711_, _11882_, _11881_);
  or (_11883_, _11843_, \oc8051_golden_model_1.IRAM[2] [5]);
  and (_11884_, _11883_, _11847_);
  and (_11885_, _11581_, _04173_);
  and (_11886_, _11885_, _11578_);
  or (_11887_, _11851_, _11886_);
  and (_11888_, _11887_, _11884_);
  and (_11889_, _11855_, _11589_);
  or (_35712_, _11889_, _11888_);
  or (_11890_, _11843_, \oc8051_golden_model_1.IRAM[2] [6]);
  and (_11891_, _11890_, _11847_);
  and (_11892_, _11779_, _04173_);
  and (_11893_, _11892_, _11776_);
  or (_11894_, _11851_, _11893_);
  and (_11895_, _11894_, _11891_);
  and (_11896_, _11855_, _11787_);
  or (_35713_, _11896_, _11895_);
  or (_11897_, _11843_, \oc8051_golden_model_1.IRAM[2] [7]);
  and (_11898_, _11897_, _11847_);
  nor (_11899_, _06132_, _04174_);
  or (_11900_, _11851_, _11899_);
  and (_11901_, _11900_, _11898_);
  and (_11902_, _11855_, _06157_);
  or (_35714_, _11902_, _11901_);
  and (_11903_, _10419_, _04523_);
  or (_11904_, _11903_, \oc8051_golden_model_1.IRAM[3] [0]);
  not (_11905_, _03924_);
  or (_11906_, _10412_, _11905_);
  or (_11907_, _11906_, _10408_);
  and (_11908_, _11907_, _11904_);
  not (_11909_, _11903_);
  or (_11910_, _11909_, _10592_);
  and (_11911_, _11910_, _11908_);
  and (_11912_, _04513_, _03924_);
  and (_11913_, _11912_, _10596_);
  and (_11914_, _11913_, _10602_);
  or (_35715_, _11914_, _11911_);
  or (_11915_, _11903_, \oc8051_golden_model_1.IRAM[3] [1]);
  and (_11916_, _11915_, _11907_);
  or (_11917_, _11909_, _10795_);
  and (_11918_, _11917_, _11916_);
  and (_11919_, _11913_, _10801_);
  or (_35716_, _11919_, _11918_);
  or (_11920_, _11903_, \oc8051_golden_model_1.IRAM[3] [2]);
  and (_11921_, _11920_, _11907_);
  or (_11922_, _11909_, _10991_);
  and (_11923_, _11922_, _11921_);
  and (_11924_, _11913_, _10997_);
  or (_35717_, _11924_, _11923_);
  or (_11925_, _11903_, \oc8051_golden_model_1.IRAM[3] [3]);
  and (_11926_, _11925_, _11907_);
  or (_11927_, _11909_, _11188_);
  and (_11928_, _11927_, _11926_);
  and (_11929_, _11913_, _11194_);
  or (_35718_, _11929_, _11928_);
  or (_11930_, _11909_, _11386_);
  or (_11931_, _11903_, \oc8051_golden_model_1.IRAM[3] [4]);
  and (_11932_, _11931_, _11907_);
  and (_11933_, _11932_, _11930_);
  and (_11934_, _11913_, _11392_);
  or (_35719_, _11934_, _11933_);
  or (_11935_, _11903_, \oc8051_golden_model_1.IRAM[3] [5]);
  and (_11936_, _11935_, _11907_);
  or (_11937_, _11909_, _11583_);
  and (_11938_, _11937_, _11936_);
  and (_11939_, _11913_, _11589_);
  or (_35720_, _11939_, _11938_);
  or (_11940_, _11903_, \oc8051_golden_model_1.IRAM[3] [6]);
  and (_11941_, _11940_, _11907_);
  or (_11942_, _11909_, _11781_);
  and (_11943_, _11942_, _11941_);
  and (_11944_, _11913_, _11787_);
  or (_35721_, _11944_, _11943_);
  or (_11945_, _11903_, \oc8051_golden_model_1.IRAM[3] [7]);
  and (_11946_, _11945_, _11907_);
  or (_11947_, _11909_, _06133_);
  and (_11948_, _11947_, _11946_);
  and (_11949_, _11913_, _06157_);
  or (_35722_, _11949_, _11948_);
  and (_11950_, _10418_, _04348_);
  and (_11951_, _11950_, _10417_);
  not (_11952_, _11951_);
  or (_11953_, _11952_, _10592_);
  not (_11954_, _04508_);
  and (_11955_, _10595_, _11954_);
  and (_11956_, _11955_, _03925_);
  nor (_11957_, _11951_, \oc8051_golden_model_1.IRAM[4] [0]);
  nor (_11958_, _11957_, _11956_);
  and (_11959_, _11958_, _11953_);
  and (_11960_, _11956_, _10602_);
  or (_35723_, _11960_, _11959_);
  or (_11961_, _11952_, _10795_);
  nor (_11962_, _11951_, \oc8051_golden_model_1.IRAM[4] [1]);
  nor (_11963_, _11962_, _11956_);
  and (_11964_, _11963_, _11961_);
  and (_11965_, _11956_, _10801_);
  or (_35724_, _11965_, _11964_);
  and (_11966_, _10410_, _11954_);
  nand (_11967_, _11966_, _03925_);
  and (_11968_, _04498_, _04348_);
  and (_11969_, _11968_, _10403_);
  or (_11970_, _11969_, \oc8051_golden_model_1.IRAM[4] [2]);
  and (_11971_, _11970_, _11967_);
  not (_11972_, _11969_);
  or (_11973_, _11972_, _11867_);
  and (_11974_, _11973_, _11971_);
  and (_11975_, _11956_, _10997_);
  or (_35725_, _11975_, _11974_);
  or (_11976_, _11952_, _11188_);
  nor (_11977_, _11951_, \oc8051_golden_model_1.IRAM[4] [3]);
  nor (_11978_, _11977_, _11956_);
  and (_11979_, _11978_, _11976_);
  and (_11980_, _11956_, _11194_);
  or (_35726_, _11980_, _11979_);
  or (_11981_, _11969_, \oc8051_golden_model_1.IRAM[4] [4]);
  and (_11982_, _11981_, _11967_);
  or (_11983_, _11952_, _11386_);
  and (_11984_, _11983_, _11982_);
  and (_11985_, _11956_, _11392_);
  or (_35727_, _11985_, _11984_);
  or (_11986_, _11969_, \oc8051_golden_model_1.IRAM[4] [5]);
  and (_11987_, _11986_, _11967_);
  or (_11988_, _11972_, _11886_);
  and (_11989_, _11988_, _11987_);
  and (_11990_, _11956_, _11589_);
  or (_35728_, _11990_, _11989_);
  or (_11991_, _11969_, \oc8051_golden_model_1.IRAM[4] [6]);
  and (_11992_, _11991_, _11967_);
  or (_11993_, _11972_, _11893_);
  and (_11994_, _11993_, _11992_);
  and (_11995_, _11956_, _11787_);
  or (_35729_, _11995_, _11994_);
  or (_11996_, _11969_, \oc8051_golden_model_1.IRAM[4] [7]);
  and (_11997_, _11996_, _11967_);
  or (_11998_, _11972_, _11899_);
  and (_11999_, _11998_, _11997_);
  and (_12000_, _11956_, _06157_);
  or (_35730_, _12000_, _11999_);
  and (_12001_, _11950_, _11794_);
  not (_12002_, _12001_);
  or (_12003_, _12002_, _10592_);
  and (_12004_, _11955_, _04231_);
  nor (_12005_, _12001_, \oc8051_golden_model_1.IRAM[5] [0]);
  nor (_12006_, _12005_, _12004_);
  and (_12007_, _12006_, _12003_);
  and (_12008_, _12004_, _10602_);
  or (_35731_, _12008_, _12007_);
  or (_12009_, _12002_, _10795_);
  nor (_12010_, _12001_, \oc8051_golden_model_1.IRAM[5] [1]);
  nor (_12011_, _12010_, _12004_);
  and (_12012_, _12011_, _12009_);
  and (_12013_, _12004_, _10801_);
  or (_35732_, _12013_, _12012_);
  nand (_12014_, _11966_, _04231_);
  or (_12015_, _12001_, \oc8051_golden_model_1.IRAM[5] [2]);
  and (_12016_, _12015_, _12014_);
  or (_12017_, _12002_, _10991_);
  and (_12018_, _12017_, _12016_);
  and (_12019_, _12004_, _10997_);
  or (_35733_, _12019_, _12018_);
  or (_12020_, _12002_, _11188_);
  nor (_12021_, _12001_, \oc8051_golden_model_1.IRAM[5] [3]);
  nor (_12022_, _12021_, _12004_);
  and (_12023_, _12022_, _12020_);
  and (_12024_, _12004_, _11194_);
  or (_35734_, _12024_, _12023_);
  or (_12025_, _12001_, \oc8051_golden_model_1.IRAM[5] [4]);
  and (_12026_, _12025_, _12014_);
  or (_12027_, _12002_, _11386_);
  and (_12028_, _12027_, _12026_);
  and (_12029_, _12004_, _11392_);
  or (_35735_, _12029_, _12028_);
  or (_12030_, _12001_, \oc8051_golden_model_1.IRAM[5] [5]);
  and (_12031_, _12030_, _12014_);
  or (_12032_, _12002_, _11583_);
  and (_12033_, _12032_, _12031_);
  and (_12034_, _12004_, _11589_);
  or (_35736_, _12034_, _12033_);
  or (_12035_, _12001_, \oc8051_golden_model_1.IRAM[5] [6]);
  and (_12036_, _12035_, _12014_);
  or (_12037_, _12002_, _11781_);
  and (_12038_, _12037_, _12036_);
  and (_12039_, _12004_, _11787_);
  or (_35737_, _12039_, _12038_);
  or (_12040_, _12001_, \oc8051_golden_model_1.IRAM[5] [7]);
  and (_12041_, _12040_, _12014_);
  or (_12042_, _12002_, _06133_);
  and (_12043_, _12042_, _12041_);
  and (_12044_, _12004_, _06157_);
  or (_35738_, _12044_, _12043_);
  and (_12045_, _11968_, _11842_);
  or (_12046_, _12045_, \oc8051_golden_model_1.IRAM[6] [0]);
  nand (_12047_, _11966_, _05340_);
  and (_12048_, _12047_, _12046_);
  not (_12049_, _12045_);
  or (_12050_, _12049_, _11850_);
  and (_12051_, _12050_, _12048_);
  and (_12052_, _11955_, _05340_);
  and (_12053_, _12052_, _10602_);
  or (_35739_, _12053_, _12051_);
  nor (_12054_, _12045_, _03947_);
  and (_12055_, _12045_, _11860_);
  or (_12056_, _12055_, _12054_);
  and (_12057_, _12056_, _12047_);
  and (_12058_, _12052_, _10801_);
  or (_35740_, _12058_, _12057_);
  or (_12059_, _12045_, \oc8051_golden_model_1.IRAM[6] [2]);
  and (_12060_, _12059_, _12047_);
  or (_12061_, _12049_, _11867_);
  and (_12062_, _12061_, _12060_);
  and (_12063_, _12052_, _10997_);
  or (_35741_, _12063_, _12062_);
  not (_12064_, _11188_);
  and (_12065_, _11950_, _11873_);
  nand (_12066_, _12065_, _12064_);
  nor (_12067_, _12065_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor (_12068_, _12067_, _12052_);
  and (_12069_, _12068_, _12066_);
  and (_12070_, _12052_, _11194_);
  or (_35742_, _12070_, _12069_);
  or (_12071_, _12045_, \oc8051_golden_model_1.IRAM[6] [4]);
  and (_12072_, _12071_, _12047_);
  and (_12073_, _11381_, _11384_);
  and (_12074_, _12073_, _04173_);
  or (_12075_, _12049_, _12074_);
  and (_12076_, _12075_, _12072_);
  and (_12077_, _12052_, _11392_);
  or (_35743_, _12077_, _12076_);
  or (_12078_, _12045_, \oc8051_golden_model_1.IRAM[6] [5]);
  and (_12079_, _12078_, _12047_);
  or (_12080_, _12049_, _11886_);
  and (_12081_, _12080_, _12079_);
  and (_12082_, _12052_, _11589_);
  or (_35744_, _12082_, _12081_);
  or (_12083_, _12045_, \oc8051_golden_model_1.IRAM[6] [6]);
  and (_12084_, _12083_, _12047_);
  or (_12085_, _12049_, _11893_);
  and (_12086_, _12085_, _12084_);
  and (_12087_, _12052_, _11787_);
  or (_35745_, _12087_, _12086_);
  or (_12088_, _12049_, _11899_);
  or (_12089_, _12045_, \oc8051_golden_model_1.IRAM[6] [7]);
  and (_12090_, _12089_, _12047_);
  and (_12091_, _12090_, _12088_);
  and (_12092_, _12052_, _06157_);
  or (_35746_, _12092_, _12091_);
  and (_12093_, _11968_, _04176_);
  not (_12094_, _12093_);
  or (_12095_, _12094_, _10592_);
  and (_12096_, _11966_, _03924_);
  not (_12097_, _12096_);
  or (_12098_, _12093_, \oc8051_golden_model_1.IRAM[7] [0]);
  and (_12099_, _12098_, _12097_);
  and (_12100_, _12099_, _12095_);
  and (_12101_, _12096_, _10602_);
  or (_35747_, _12101_, _12100_);
  or (_12102_, _12094_, _10795_);
  or (_12103_, _12093_, \oc8051_golden_model_1.IRAM[7] [1]);
  and (_12104_, _12103_, _12097_);
  and (_12105_, _12104_, _12102_);
  and (_12106_, _12096_, _10801_);
  or (_35748_, _12106_, _12105_);
  or (_12107_, _12094_, _10991_);
  or (_12108_, _12093_, \oc8051_golden_model_1.IRAM[7] [2]);
  and (_12109_, _12108_, _12097_);
  and (_12110_, _12109_, _12107_);
  and (_12111_, _12096_, _10997_);
  or (_35749_, _12111_, _12110_);
  or (_12112_, _12094_, _11188_);
  or (_12113_, _12093_, \oc8051_golden_model_1.IRAM[7] [3]);
  and (_12114_, _12113_, _12097_);
  and (_12115_, _12114_, _12112_);
  and (_12116_, _12096_, _11194_);
  or (_35750_, _12116_, _12115_);
  or (_12117_, _12094_, _11386_);
  or (_12118_, _12093_, \oc8051_golden_model_1.IRAM[7] [4]);
  and (_12119_, _12118_, _12097_);
  and (_12120_, _12119_, _12117_);
  and (_12121_, _12096_, _11392_);
  or (_35751_, _12121_, _12120_);
  or (_12122_, _12093_, \oc8051_golden_model_1.IRAM[7] [5]);
  and (_12123_, _12122_, _12097_);
  or (_12124_, _12094_, _11886_);
  and (_12125_, _12124_, _12123_);
  and (_12126_, _12096_, _11589_);
  or (_35752_, _12126_, _12125_);
  or (_12127_, _12093_, \oc8051_golden_model_1.IRAM[7] [6]);
  and (_12128_, _12127_, _12097_);
  or (_12129_, _12094_, _11893_);
  and (_12130_, _12129_, _12128_);
  and (_12131_, _12096_, _11787_);
  or (_35753_, _12131_, _12130_);
  or (_12132_, _12093_, \oc8051_golden_model_1.IRAM[7] [7]);
  and (_12133_, _12132_, _12097_);
  or (_12134_, _12094_, _11899_);
  and (_12135_, _12134_, _12133_);
  and (_12136_, _12096_, _06157_);
  or (_35754_, _12136_, _12135_);
  and (_12137_, _04525_, _04497_);
  and (_12138_, _12137_, _10417_);
  not (_12139_, _12138_);
  or (_12140_, _12139_, _10592_);
  not (_12141_, _04505_);
  and (_12142_, _04514_, _12141_);
  and (_12143_, _12142_, _03925_);
  not (_12144_, _12143_);
  or (_12145_, _12138_, \oc8051_golden_model_1.IRAM[8] [0]);
  and (_12146_, _12145_, _12144_);
  and (_12147_, _12146_, _12140_);
  and (_12148_, _12143_, _10602_);
  or (_35755_, _12148_, _12147_);
  or (_12149_, _12138_, \oc8051_golden_model_1.IRAM[8] [1]);
  and (_12150_, _12149_, _12144_);
  or (_12151_, _12139_, _10795_);
  and (_12152_, _12151_, _12150_);
  and (_12153_, _12143_, _10801_);
  or (_35756_, _12153_, _12152_);
  or (_12154_, _12138_, \oc8051_golden_model_1.IRAM[8] [2]);
  and (_12155_, _12154_, _12144_);
  or (_12156_, _12139_, _10991_);
  and (_12157_, _12156_, _12155_);
  and (_12158_, _12143_, _10997_);
  or (_35757_, _12158_, _12157_);
  or (_12159_, _12139_, _11188_);
  or (_12160_, _12138_, \oc8051_golden_model_1.IRAM[8] [3]);
  and (_12161_, _12160_, _12144_);
  and (_12162_, _12161_, _12159_);
  and (_12163_, _12143_, _11194_);
  or (_35758_, _12163_, _12162_);
  or (_12164_, _12138_, \oc8051_golden_model_1.IRAM[8] [4]);
  and (_12165_, _12164_, _12144_);
  or (_12166_, _12139_, _11386_);
  and (_12167_, _12166_, _12165_);
  and (_12168_, _12143_, _11392_);
  or (_35759_, _12168_, _12167_);
  or (_12169_, _12138_, \oc8051_golden_model_1.IRAM[8] [5]);
  and (_12170_, _12169_, _12144_);
  or (_12171_, _12139_, _11583_);
  and (_12172_, _12171_, _12170_);
  and (_12173_, _12143_, _11589_);
  or (_35760_, _12173_, _12172_);
  or (_12174_, _12138_, \oc8051_golden_model_1.IRAM[8] [6]);
  and (_12175_, _12174_, _12144_);
  or (_12176_, _12139_, _11781_);
  and (_12177_, _12176_, _12175_);
  and (_12178_, _12143_, _11787_);
  or (_35761_, _12178_, _12177_);
  or (_12179_, _12138_, \oc8051_golden_model_1.IRAM[8] [7]);
  or (_12180_, _12139_, _06133_);
  and (_12181_, _12180_, _12179_);
  and (_12182_, _12181_, _12144_);
  and (_12183_, _12143_, _06157_);
  or (_35762_, _12183_, _12182_);
  and (_12184_, _12137_, _11794_);
  not (_12185_, _12184_);
  or (_12186_, _12185_, _10592_);
  and (_12187_, _12142_, _04231_);
  nor (_12188_, _12184_, \oc8051_golden_model_1.IRAM[9] [0]);
  nor (_12189_, _12188_, _12187_);
  and (_12190_, _12189_, _12186_);
  and (_12191_, _12187_, _10602_);
  or (_35763_, _12191_, _12190_);
  nand (_12192_, _10411_, _04232_);
  or (_12193_, _12184_, \oc8051_golden_model_1.IRAM[9] [1]);
  and (_12194_, _12193_, _12192_);
  or (_12195_, _12185_, _10795_);
  and (_12196_, _12195_, _12194_);
  and (_12197_, _12187_, _10801_);
  or (_35764_, _12197_, _12196_);
  or (_12198_, _12184_, \oc8051_golden_model_1.IRAM[9] [2]);
  and (_12199_, _12198_, _12192_);
  or (_12200_, _12185_, _10991_);
  and (_12201_, _12200_, _12199_);
  and (_12202_, _12187_, _10997_);
  or (_35765_, _12202_, _12201_);
  or (_12203_, _12185_, _11188_);
  nor (_12204_, _12184_, \oc8051_golden_model_1.IRAM[9] [3]);
  nor (_12205_, _12204_, _12187_);
  and (_12206_, _12205_, _12203_);
  and (_12207_, _12187_, _11194_);
  or (_35766_, _12207_, _12206_);
  or (_12208_, _12184_, \oc8051_golden_model_1.IRAM[9] [4]);
  and (_12209_, _12208_, _12192_);
  or (_12210_, _12185_, _11386_);
  and (_12211_, _12210_, _12209_);
  and (_12212_, _12187_, _11392_);
  or (_35767_, _12212_, _12211_);
  or (_12213_, _12184_, \oc8051_golden_model_1.IRAM[9] [5]);
  and (_12214_, _12213_, _12192_);
  or (_12215_, _12185_, _11583_);
  and (_12216_, _12215_, _12214_);
  and (_12217_, _12187_, _11589_);
  or (_35768_, _12217_, _12216_);
  or (_12218_, _12184_, \oc8051_golden_model_1.IRAM[9] [6]);
  and (_12219_, _12218_, _12192_);
  or (_12220_, _12185_, _11781_);
  and (_12221_, _12220_, _12219_);
  and (_12222_, _12187_, _11787_);
  or (_35769_, _12222_, _12221_);
  or (_12223_, _12184_, \oc8051_golden_model_1.IRAM[9] [7]);
  and (_12224_, _12223_, _12192_);
  or (_12225_, _12185_, _06133_);
  and (_12226_, _12225_, _12224_);
  and (_12227_, _12187_, _06157_);
  or (_35770_, _12227_, _12226_);
  and (_12228_, _12137_, _11873_);
  not (_12229_, _12228_);
  or (_12230_, _12229_, _10592_);
  and (_12231_, _12142_, _05340_);
  not (_12232_, _12231_);
  or (_12233_, _12228_, \oc8051_golden_model_1.IRAM[10] [0]);
  and (_12234_, _12233_, _12232_);
  and (_12235_, _12234_, _12230_);
  and (_12236_, _12231_, _10602_);
  or (_35651_, _12236_, _12235_);
  or (_12237_, _12228_, \oc8051_golden_model_1.IRAM[10] [1]);
  and (_12238_, _12237_, _12232_);
  or (_12239_, _12229_, _10795_);
  and (_12240_, _12239_, _12238_);
  and (_12241_, _12231_, _10801_);
  or (_35652_, _12241_, _12240_);
  or (_12242_, _12228_, \oc8051_golden_model_1.IRAM[10] [2]);
  and (_12243_, _12242_, _12232_);
  or (_12244_, _12229_, _10991_);
  and (_12245_, _12244_, _12243_);
  and (_12246_, _12231_, _10997_);
  or (_35653_, _12246_, _12245_);
  or (_12247_, _12229_, _11188_);
  or (_12248_, _12228_, \oc8051_golden_model_1.IRAM[10] [3]);
  and (_12249_, _12248_, _12232_);
  and (_12250_, _12249_, _12247_);
  and (_12251_, _12231_, _11194_);
  or (_35654_, _12251_, _12250_);
  or (_12252_, _12228_, \oc8051_golden_model_1.IRAM[10] [4]);
  and (_12253_, _12252_, _12232_);
  or (_12254_, _12229_, _11386_);
  and (_12255_, _12254_, _12253_);
  and (_12256_, _12231_, _11392_);
  or (_35655_, _12256_, _12255_);
  or (_12257_, _12228_, \oc8051_golden_model_1.IRAM[10] [5]);
  and (_12258_, _12257_, _12232_);
  or (_12259_, _12229_, _11583_);
  and (_12260_, _12259_, _12258_);
  and (_12261_, _12231_, _11589_);
  or (_35656_, _12261_, _12260_);
  or (_12262_, _12228_, \oc8051_golden_model_1.IRAM[10] [6]);
  and (_12263_, _12262_, _12232_);
  or (_12264_, _12229_, _11781_);
  and (_12265_, _12264_, _12263_);
  and (_12266_, _12231_, _11787_);
  or (_35657_, _12266_, _12265_);
  or (_12267_, _12228_, \oc8051_golden_model_1.IRAM[10] [7]);
  and (_12268_, _12267_, _12232_);
  or (_12269_, _12229_, _06133_);
  and (_12270_, _12269_, _12268_);
  and (_12271_, _12231_, _06157_);
  or (_35658_, _12271_, _12270_);
  and (_12272_, _12137_, _04523_);
  not (_12273_, _12272_);
  or (_12274_, _12273_, _10592_);
  and (_12275_, _12142_, _03924_);
  not (_12276_, _12275_);
  or (_12277_, _12272_, \oc8051_golden_model_1.IRAM[11] [0]);
  and (_12278_, _12277_, _12276_);
  and (_12279_, _12278_, _12274_);
  and (_12280_, _12275_, _10602_);
  or (_35659_, _12280_, _12279_);
  or (_12281_, _12272_, \oc8051_golden_model_1.IRAM[11] [1]);
  and (_12282_, _12281_, _12276_);
  or (_12283_, _12273_, _10795_);
  and (_12284_, _12283_, _12282_);
  and (_12285_, _12275_, _10801_);
  or (_35660_, _12285_, _12284_);
  or (_12286_, _12272_, \oc8051_golden_model_1.IRAM[11] [2]);
  and (_12287_, _12286_, _12276_);
  or (_12288_, _12273_, _10991_);
  and (_12289_, _12288_, _12287_);
  and (_12290_, _12275_, _10997_);
  or (_35661_, _12290_, _12289_);
  or (_12291_, _12273_, _11188_);
  or (_12292_, _12272_, \oc8051_golden_model_1.IRAM[11] [3]);
  and (_12293_, _12292_, _12276_);
  and (_12294_, _12293_, _12291_);
  and (_12295_, _12275_, _11194_);
  or (_35662_, _12295_, _12294_);
  or (_12296_, _12272_, \oc8051_golden_model_1.IRAM[11] [4]);
  and (_12297_, _12296_, _12276_);
  or (_12298_, _12273_, _11386_);
  and (_12299_, _12298_, _12297_);
  and (_12300_, _12275_, _11392_);
  or (_35663_, _12300_, _12299_);
  or (_12301_, _12272_, \oc8051_golden_model_1.IRAM[11] [5]);
  and (_12302_, _12301_, _12276_);
  or (_12303_, _12273_, _11583_);
  and (_12304_, _12303_, _12302_);
  and (_12305_, _12275_, _11589_);
  or (_35664_, _12305_, _12304_);
  or (_12306_, _12272_, \oc8051_golden_model_1.IRAM[11] [6]);
  and (_12307_, _12306_, _12276_);
  or (_12308_, _12273_, _11781_);
  and (_12309_, _12308_, _12307_);
  and (_12310_, _12275_, _11787_);
  or (_35665_, _12310_, _12309_);
  nor (_12311_, _12272_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor (_12312_, _12273_, _06133_);
  or (_12313_, _12312_, _12311_);
  nand (_12314_, _12313_, _12276_);
  or (_12315_, _12276_, _06157_);
  and (_35666_, _12315_, _12314_);
  and (_12316_, _10403_, _04500_);
  not (_12317_, _12316_);
  or (_12318_, _12317_, _10592_);
  and (_12319_, _04515_, _03925_);
  not (_12320_, _12319_);
  or (_12321_, _12316_, \oc8051_golden_model_1.IRAM[12] [0]);
  and (_12322_, _12321_, _12320_);
  and (_12323_, _12322_, _12318_);
  and (_12324_, _12319_, _10602_);
  or (_35667_, _12324_, _12323_);
  or (_12325_, _12317_, _10795_);
  or (_12326_, _12316_, \oc8051_golden_model_1.IRAM[12] [1]);
  and (_12327_, _12326_, _12320_);
  and (_12328_, _12327_, _12325_);
  and (_12329_, _12319_, _10801_);
  or (_35668_, _12329_, _12328_);
  or (_12330_, _12316_, \oc8051_golden_model_1.IRAM[12] [2]);
  and (_12331_, _12330_, _12320_);
  or (_12332_, _12317_, _11867_);
  and (_12333_, _12332_, _12331_);
  and (_12334_, _12319_, _10997_);
  or (_35669_, _12334_, _12333_);
  or (_12335_, _12317_, _11188_);
  or (_12336_, _12316_, \oc8051_golden_model_1.IRAM[12] [3]);
  and (_12337_, _12336_, _12320_);
  and (_12338_, _12337_, _12335_);
  and (_12339_, _12319_, _11194_);
  or (_35670_, _12339_, _12338_);
  or (_12340_, _12317_, _11386_);
  or (_12341_, _12316_, \oc8051_golden_model_1.IRAM[12] [4]);
  and (_12342_, _12341_, _12320_);
  and (_12343_, _12342_, _12340_);
  and (_12344_, _12319_, _11392_);
  or (_35671_, _12344_, _12343_);
  or (_12345_, _12316_, \oc8051_golden_model_1.IRAM[12] [5]);
  and (_12346_, _12345_, _12320_);
  or (_12347_, _12317_, _11886_);
  and (_12348_, _12347_, _12346_);
  and (_12349_, _12319_, _11589_);
  or (_35672_, _12349_, _12348_);
  or (_12350_, _12316_, \oc8051_golden_model_1.IRAM[12] [6]);
  and (_12351_, _12350_, _12320_);
  or (_12352_, _12317_, _11893_);
  and (_12353_, _12352_, _12351_);
  and (_12354_, _12319_, _11787_);
  or (_35673_, _12354_, _12353_);
  or (_12355_, _12317_, _11899_);
  or (_12356_, _12316_, \oc8051_golden_model_1.IRAM[12] [7]);
  and (_12357_, _12356_, _12320_);
  and (_12358_, _12357_, _12355_);
  and (_12359_, _12319_, _06157_);
  or (_35674_, _12359_, _12358_);
  and (_12360_, _11794_, _04526_);
  not (_12361_, _12360_);
  or (_12362_, _12361_, _10592_);
  and (_12363_, _04515_, _04231_);
  not (_12364_, _12363_);
  or (_12365_, _12360_, \oc8051_golden_model_1.IRAM[13] [0]);
  and (_12366_, _12365_, _12364_);
  and (_12367_, _12366_, _12362_);
  and (_12368_, _12363_, _10602_);
  or (_35675_, _12368_, _12367_);
  or (_12369_, _12361_, _10795_);
  or (_12370_, _12360_, \oc8051_golden_model_1.IRAM[13] [1]);
  and (_12371_, _12370_, _12364_);
  and (_12372_, _12371_, _12369_);
  and (_12373_, _12363_, _10801_);
  or (_35676_, _12373_, _12372_);
  and (_12374_, _12363_, _10997_);
  and (_12375_, _10402_, _04079_);
  and (_12376_, _12375_, _04500_);
  or (_12377_, _12376_, \oc8051_golden_model_1.IRAM[13] [2]);
  and (_12378_, _12377_, _12364_);
  or (_12379_, _12361_, _10991_);
  and (_12380_, _12379_, _12378_);
  or (_35677_, _12380_, _12374_);
  or (_12381_, _12361_, _11188_);
  or (_12382_, _12360_, \oc8051_golden_model_1.IRAM[13] [3]);
  and (_12383_, _12382_, _12364_);
  and (_12384_, _12383_, _12381_);
  and (_12385_, _12363_, _11194_);
  or (_35678_, _12385_, _12384_);
  or (_12386_, _12376_, \oc8051_golden_model_1.IRAM[13] [4]);
  and (_12387_, _12386_, _12364_);
  or (_12388_, _12361_, _11386_);
  and (_12389_, _12388_, _12387_);
  and (_12390_, _12363_, _11392_);
  or (_35679_, _12390_, _12389_);
  or (_12391_, _12376_, \oc8051_golden_model_1.IRAM[13] [5]);
  and (_12392_, _12391_, _12364_);
  or (_12393_, _12361_, _11583_);
  and (_12394_, _12393_, _12392_);
  and (_12395_, _12363_, _11589_);
  or (_35680_, _12395_, _12394_);
  and (_12396_, _12363_, _11787_);
  or (_12397_, _12376_, \oc8051_golden_model_1.IRAM[13] [6]);
  and (_12398_, _12397_, _12364_);
  or (_12399_, _12361_, _11781_);
  and (_12400_, _12399_, _12398_);
  or (_35681_, _12400_, _12396_);
  or (_12401_, _12376_, \oc8051_golden_model_1.IRAM[13] [7]);
  and (_12402_, _12401_, _12364_);
  or (_12403_, _12361_, _06133_);
  and (_12404_, _12403_, _12402_);
  and (_12405_, _12363_, _06157_);
  or (_35682_, _12405_, _12404_);
  and (_12406_, _11873_, _04526_);
  not (_12407_, _12406_);
  or (_12408_, _12407_, _10592_);
  and (_12409_, _05340_, _04515_);
  not (_12410_, _12409_);
  or (_12411_, _12406_, \oc8051_golden_model_1.IRAM[14] [0]);
  and (_12412_, _12411_, _12410_);
  and (_12413_, _12412_, _12408_);
  and (_12414_, _12409_, _10602_);
  or (_35683_, _12414_, _12413_);
  or (_12415_, _12407_, _10795_);
  or (_12416_, _12406_, \oc8051_golden_model_1.IRAM[14] [1]);
  and (_12417_, _12416_, _12410_);
  and (_12418_, _12417_, _12415_);
  and (_12419_, _12409_, _10801_);
  or (_35684_, _12419_, _12418_);
  and (_12420_, _11842_, _04500_);
  or (_12421_, _12420_, \oc8051_golden_model_1.IRAM[14] [2]);
  and (_12422_, _12421_, _12410_);
  not (_12423_, _12420_);
  or (_12424_, _12423_, _11867_);
  and (_12425_, _12424_, _12422_);
  and (_12426_, _12409_, _10997_);
  or (_35685_, _12426_, _12425_);
  or (_12427_, _12407_, _11188_);
  or (_12428_, _12406_, \oc8051_golden_model_1.IRAM[14] [3]);
  and (_12429_, _12428_, _12410_);
  and (_12430_, _12429_, _12427_);
  and (_12431_, _12409_, _11194_);
  or (_35686_, _12431_, _12430_);
  or (_12432_, _12420_, \oc8051_golden_model_1.IRAM[14] [4]);
  and (_12433_, _12432_, _12410_);
  or (_12434_, _12407_, _11386_);
  and (_12435_, _12434_, _12433_);
  and (_12436_, _12409_, _11392_);
  or (_35687_, _12436_, _12435_);
  or (_12437_, _12420_, \oc8051_golden_model_1.IRAM[14] [5]);
  and (_12438_, _12437_, _12410_);
  or (_12439_, _12423_, _11886_);
  and (_12440_, _12439_, _12438_);
  and (_12441_, _12409_, _11589_);
  or (_35688_, _12441_, _12440_);
  or (_12442_, _12420_, \oc8051_golden_model_1.IRAM[14] [6]);
  and (_12443_, _12442_, _12410_);
  or (_12444_, _12423_, _11893_);
  and (_12445_, _12444_, _12443_);
  and (_12446_, _12409_, _11787_);
  or (_35689_, _12446_, _12445_);
  nor (_12447_, _12406_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor (_12448_, _12407_, _06133_);
  nor (_12449_, _12448_, _12447_);
  or (_12450_, _12449_, _12409_);
  or (_12451_, _12410_, _06157_);
  and (_35690_, _12451_, _12450_);
  or (_12452_, _10592_, _04528_);
  or (_12453_, _04527_, \oc8051_golden_model_1.IRAM[15] [0]);
  and (_12454_, _12453_, _04517_);
  and (_12455_, _12454_, _12452_);
  and (_12456_, _10602_, _04516_);
  or (_35691_, _12456_, _12455_);
  or (_12457_, _10795_, _04528_);
  or (_12458_, _04527_, \oc8051_golden_model_1.IRAM[15] [1]);
  and (_12459_, _12458_, _04517_);
  and (_12460_, _12459_, _12457_);
  and (_12461_, _10801_, _04516_);
  or (_35692_, _12461_, _12460_);
  or (_12462_, _04501_, \oc8051_golden_model_1.IRAM[15] [2]);
  and (_12463_, _12462_, _04517_);
  not (_12464_, _04501_);
  or (_12465_, _11867_, _12464_);
  and (_12466_, _12465_, _12463_);
  and (_12467_, _10997_, _04516_);
  or (_35693_, _12467_, _12466_);
  or (_12468_, _11188_, _04528_);
  or (_12469_, _04527_, \oc8051_golden_model_1.IRAM[15] [3]);
  and (_12470_, _12469_, _04517_);
  and (_12471_, _12470_, _12468_);
  and (_12472_, _11194_, _04516_);
  or (_35694_, _12472_, _12471_);
  or (_12473_, _04501_, \oc8051_golden_model_1.IRAM[15] [4]);
  and (_12474_, _12473_, _04517_);
  or (_12475_, _11386_, _04528_);
  and (_12476_, _12475_, _12474_);
  and (_12477_, _11392_, _04516_);
  or (_35695_, _12477_, _12476_);
  or (_12478_, _04501_, \oc8051_golden_model_1.IRAM[15] [5]);
  and (_12479_, _12478_, _04517_);
  or (_12480_, _11886_, _12464_);
  and (_12481_, _12480_, _12479_);
  and (_12482_, _11589_, _04516_);
  or (_35696_, _12482_, _12481_);
  or (_12483_, _04501_, \oc8051_golden_model_1.IRAM[15] [6]);
  and (_12484_, _12483_, _04517_);
  or (_12485_, _11893_, _12464_);
  and (_12486_, _12485_, _12484_);
  and (_12487_, _11787_, _04516_);
  or (_35697_, _12487_, _12486_);
  nor (_12488_, _34446_, _06743_);
  nor (_12489_, _04661_, _06743_);
  and (_12490_, _10546_, _04661_);
  or (_12491_, _12490_, _12489_);
  and (_12492_, _12491_, _03107_);
  and (_12493_, _04661_, _05647_);
  or (_12494_, _12493_, _12489_);
  or (_12495_, _12494_, _05261_);
  and (_12496_, _06114_, _04661_);
  or (_12497_, _12489_, _06726_);
  or (_12498_, _12497_, _12496_);
  and (_12499_, _04661_, _03805_);
  or (_12500_, _12499_, _12489_);
  or (_12501_, _12500_, _03860_);
  nor (_12502_, _05286_, _06743_);
  and (_12503_, _10441_, _05286_);
  or (_12504_, _12503_, _12502_);
  and (_12505_, _12504_, _02799_);
  nor (_12506_, _05036_, _06175_);
  or (_12507_, _12506_, _12489_);
  or (_12508_, _12507_, _06162_);
  and (_12509_, _04661_, \oc8051_golden_model_1.ACC [0]);
  or (_12510_, _12509_, _12489_);
  and (_12511_, _12510_, _02837_);
  nor (_12512_, _02837_, _06743_);
  or (_12513_, _12512_, _02932_);
  or (_12514_, _12513_, _12511_);
  and (_12515_, _12514_, _02939_);
  or (_12516_, _12515_, _02796_);
  and (_12517_, _12516_, _12508_);
  and (_12518_, _12500_, _02930_);
  or (_12519_, _12518_, _02928_);
  or (_12520_, _12519_, _12517_);
  or (_12521_, _12520_, _12505_);
  or (_12522_, _12509_, _02943_);
  and (_12523_, _12522_, _02927_);
  or (_12524_, _12523_, _12489_);
  and (_12525_, _12524_, _06189_);
  and (_12526_, _12525_, _12521_);
  and (_12527_, _12507_, _02790_);
  or (_12528_, _12527_, _06195_);
  or (_12529_, _12528_, _12526_);
  nor (_12530_, _06677_, _06675_);
  nor (_12531_, _12530_, _06678_);
  or (_12532_, _12531_, _06201_);
  and (_12533_, _12532_, _02966_);
  and (_12534_, _12533_, _12529_);
  nor (_12535_, _10473_, _06716_);
  or (_12536_, _12535_, _12502_);
  and (_12537_, _12536_, _02785_);
  or (_12538_, _12537_, _03861_);
  or (_12539_, _12538_, _12534_);
  and (_12540_, _12539_, _12501_);
  or (_12541_, _12540_, _03850_);
  and (_12542_, _12541_, _12498_);
  or (_12543_, _12542_, _02524_);
  nor (_12544_, _10530_, _06175_);
  or (_12545_, _12489_, _02970_);
  or (_12546_, _12545_, _12544_);
  and (_12547_, _12546_, _06737_);
  and (_12548_, _12547_, _12543_);
  nand (_12549_, _07086_, _02658_);
  nor (_12550_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nor (_12551_, _12550_, _06656_);
  or (_12552_, _07086_, _12551_);
  and (_12553_, _12552_, _06731_);
  and (_12554_, _12553_, _12549_);
  or (_12555_, _12554_, _02974_);
  or (_12556_, _12555_, _12548_);
  and (_12557_, _12556_, _12495_);
  or (_12558_, _12557_, _02977_);
  and (_12559_, _10427_, _04661_);
  or (_12560_, _12489_, _07092_);
  or (_12561_, _12560_, _12559_);
  and (_12562_, _12561_, _07104_);
  and (_12563_, _12562_, _12558_);
  or (_12564_, _12563_, _12492_);
  and (_12565_, _12564_, _03095_);
  nand (_12566_, _12494_, _02991_);
  nor (_12567_, _12566_, _12506_);
  or (_12568_, _12489_, _05036_);
  and (_12569_, _12510_, _03094_);
  and (_12570_, _12569_, _12568_);
  or (_12571_, _12570_, _02994_);
  or (_12572_, _12571_, _12567_);
  or (_12573_, _12572_, _12565_);
  nor (_12574_, _10425_, _06175_);
  or (_12575_, _12489_, _07120_);
  or (_12576_, _12575_, _12574_);
  and (_12577_, _12576_, _07118_);
  and (_12578_, _12577_, _12573_);
  nor (_12579_, _10423_, _06175_);
  or (_12580_, _12579_, _12489_);
  and (_12581_, _12580_, _03099_);
  or (_12582_, _12581_, _03133_);
  or (_12583_, _12582_, _12578_);
  or (_12584_, _12507_, _03138_);
  and (_12585_, _12584_, _03142_);
  and (_12586_, _12585_, _12583_);
  and (_12587_, _12489_, _02778_);
  or (_12588_, _12587_, _02852_);
  or (_12589_, _12588_, _12586_);
  or (_12590_, _12507_, _02853_);
  and (_12591_, _12590_, _34446_);
  and (_12592_, _12591_, _12589_);
  or (_12593_, _12592_, _12488_);
  and (_35615_[0], _12593_, _35583_);
  nor (_12594_, _34446_, _06738_);
  nand (_12595_, _04661_, _03660_);
  or (_12596_, _04661_, \oc8051_golden_model_1.B [1]);
  and (_12597_, _12596_, _02974_);
  and (_12598_, _12597_, _12595_);
  and (_12599_, _10622_, _04661_);
  not (_12600_, _12599_);
  and (_12601_, _12600_, _12596_);
  or (_12602_, _12601_, _06162_);
  nand (_12603_, _04661_, _02477_);
  and (_12604_, _12603_, _12596_);
  and (_12605_, _12604_, _02837_);
  nor (_12606_, _02837_, _06738_);
  or (_12607_, _12606_, _02932_);
  or (_12608_, _12607_, _12605_);
  and (_12609_, _12608_, _02939_);
  and (_12610_, _12609_, _12602_);
  nor (_12611_, _04661_, _06738_);
  nor (_12612_, _06175_, _03989_);
  or (_12613_, _12612_, _12611_);
  and (_12614_, _12613_, _02930_);
  nor (_12615_, _05286_, _06738_);
  and (_12616_, _10617_, _05286_);
  or (_12617_, _12616_, _12615_);
  and (_12618_, _12617_, _02799_);
  or (_12619_, _12618_, _12614_);
  or (_12620_, _12619_, _02928_);
  or (_12621_, _12620_, _12610_);
  or (_12622_, _12604_, _02943_);
  and (_12623_, _12622_, _12621_);
  or (_12624_, _12623_, _02796_);
  and (_12625_, _10620_, _05286_);
  or (_12626_, _12625_, _12615_);
  or (_12627_, _12626_, _02927_);
  and (_12628_, _12627_, _06189_);
  and (_12629_, _12628_, _12624_);
  and (_12630_, _12616_, _10616_);
  or (_12631_, _12630_, _12615_);
  and (_12632_, _12631_, _02790_);
  or (_12633_, _12632_, _06195_);
  or (_12634_, _12633_, _12629_);
  or (_12635_, _06622_, _06621_);
  nand (_12636_, _12635_, _06679_);
  or (_12637_, _12635_, _06679_);
  and (_12638_, _12637_, _12636_);
  or (_12639_, _12638_, _06201_);
  and (_12640_, _12639_, _02966_);
  and (_12641_, _12640_, _12634_);
  nor (_12642_, _10662_, _06716_);
  or (_12643_, _12642_, _12615_);
  and (_12644_, _12643_, _02785_);
  or (_12645_, _12644_, _03861_);
  or (_12646_, _12645_, _12641_);
  or (_12647_, _12613_, _03860_);
  and (_12648_, _12647_, _12646_);
  or (_12649_, _12648_, _03850_);
  and (_12650_, _06113_, _04661_);
  or (_12651_, _12611_, _06726_);
  or (_12652_, _12651_, _12650_);
  and (_12653_, _12652_, _02970_);
  and (_12654_, _12653_, _12649_);
  nand (_12655_, _10719_, _04661_);
  and (_12656_, _12596_, _02524_);
  and (_12657_, _12656_, _12655_);
  or (_12658_, _12657_, _06731_);
  or (_12659_, _12658_, _12654_);
  nor (_12660_, _07081_, _07080_);
  or (_12661_, _12660_, _07082_);
  nor (_12662_, _12661_, _07086_);
  and (_12663_, _07086_, _07033_);
  or (_12664_, _12663_, _12662_);
  or (_12665_, _12664_, _06737_);
  and (_12666_, _12665_, _05261_);
  and (_12667_, _12666_, _12659_);
  or (_12668_, _12667_, _12598_);
  and (_12669_, _12668_, _03882_);
  or (_12670_, _10613_, _06175_);
  and (_12671_, _12596_, _02991_);
  and (_12672_, _12671_, _12670_);
  or (_12673_, _10610_, _06175_);
  and (_12674_, _12596_, _03107_);
  and (_12675_, _12674_, _12673_);
  or (_12676_, _10614_, _06175_);
  and (_12677_, _12596_, _02977_);
  and (_12678_, _12677_, _12676_);
  or (_12679_, _12678_, _12675_);
  or (_12680_, _12679_, _12672_);
  or (_12681_, _12680_, _12669_);
  and (_12682_, _12681_, _06161_);
  or (_12683_, _12611_, _04988_);
  and (_12684_, _12604_, _03094_);
  and (_12685_, _12684_, _12683_);
  or (_12686_, _12685_, _12682_);
  and (_12687_, _12686_, _03100_);
  or (_12688_, _12595_, _04988_);
  and (_12689_, _12596_, _02994_);
  and (_12690_, _12689_, _12688_);
  or (_12691_, _12603_, _04988_);
  and (_12692_, _12596_, _03099_);
  and (_12693_, _12692_, _12691_);
  or (_12694_, _12693_, _03133_);
  or (_12695_, _12694_, _12690_);
  or (_12696_, _12695_, _12687_);
  or (_12697_, _12601_, _03138_);
  and (_12698_, _12697_, _03142_);
  and (_12699_, _12698_, _12696_);
  and (_12700_, _12626_, _02778_);
  or (_12701_, _12700_, _02852_);
  or (_12702_, _12701_, _12699_);
  or (_12703_, _12611_, _02853_);
  or (_12704_, _12703_, _12599_);
  and (_12705_, _12704_, _34446_);
  and (_12706_, _12705_, _12702_);
  or (_12707_, _12706_, _12594_);
  and (_35615_[1], _12707_, _35583_);
  nor (_12708_, _34446_, _06753_);
  nor (_12709_, _04661_, _06753_);
  and (_12710_, _10942_, _04661_);
  or (_12711_, _12710_, _12709_);
  and (_12712_, _12711_, _03107_);
  and (_12713_, _04661_, _05690_);
  or (_12714_, _12713_, _12709_);
  or (_12715_, _12714_, _05261_);
  nor (_12716_, _06175_, _04413_);
  or (_12717_, _12716_, _12709_);
  or (_12718_, _12717_, _03860_);
  nor (_12719_, _10824_, _06175_);
  or (_12720_, _12719_, _12709_);
  or (_12721_, _12720_, _06162_);
  and (_12722_, _04661_, \oc8051_golden_model_1.ACC [2]);
  or (_12723_, _12722_, _12709_);
  and (_12724_, _12723_, _02837_);
  nor (_12725_, _02837_, _06753_);
  or (_12726_, _12725_, _02932_);
  or (_12727_, _12726_, _12724_);
  and (_12728_, _12727_, _02939_);
  and (_12729_, _12728_, _12721_);
  and (_12730_, _12717_, _02930_);
  nor (_12731_, _05286_, _06753_);
  and (_12732_, _10815_, _05286_);
  or (_12733_, _12732_, _12731_);
  and (_12734_, _12733_, _02799_);
  or (_12735_, _12734_, _12730_);
  or (_12736_, _12735_, _02928_);
  or (_12737_, _12736_, _12729_);
  or (_12738_, _12723_, _02943_);
  and (_12739_, _12738_, _12737_);
  or (_12740_, _12739_, _02796_);
  and (_12741_, _10818_, _05286_);
  or (_12742_, _12741_, _12731_);
  or (_12743_, _12742_, _02927_);
  and (_12744_, _12743_, _06189_);
  and (_12745_, _12744_, _12740_);
  and (_12746_, _12732_, _10814_);
  or (_12747_, _12746_, _12731_);
  and (_12748_, _12747_, _02790_);
  or (_12749_, _12748_, _06195_);
  or (_12750_, _12749_, _12745_);
  nor (_12751_, _06681_, _06578_);
  nor (_12752_, _12751_, _06682_);
  or (_12753_, _12752_, _06201_);
  and (_12754_, _12753_, _02966_);
  and (_12755_, _12754_, _12750_);
  nor (_12756_, _10866_, _06716_);
  or (_12757_, _12756_, _12731_);
  and (_12758_, _12757_, _02785_);
  or (_12759_, _12758_, _03861_);
  or (_12760_, _12759_, _12755_);
  and (_12761_, _12760_, _12718_);
  or (_12762_, _12761_, _03850_);
  and (_12763_, _06117_, _04661_);
  or (_12764_, _12709_, _06726_);
  or (_12765_, _12764_, _12763_);
  and (_12766_, _12765_, _12762_);
  or (_12767_, _12766_, _02524_);
  nor (_12768_, _10922_, _06175_);
  or (_12769_, _12709_, _02970_);
  or (_12770_, _12769_, _12768_);
  and (_12771_, _12770_, _06737_);
  and (_12772_, _12771_, _12767_);
  nand (_12773_, _07086_, _07023_);
  nor (_12774_, _07082_, _07034_);
  not (_12775_, _12774_);
  and (_12776_, _12775_, _07026_);
  nor (_12777_, _12775_, _07026_);
  nor (_12778_, _12777_, _12776_);
  or (_12779_, _12778_, _07086_);
  and (_12780_, _12779_, _06731_);
  and (_12781_, _12780_, _12773_);
  or (_12782_, _12781_, _02974_);
  or (_12783_, _12782_, _12772_);
  and (_12784_, _12783_, _12715_);
  or (_12785_, _12784_, _02977_);
  and (_12786_, _10936_, _04661_);
  or (_12787_, _12709_, _07092_);
  or (_12788_, _12787_, _12786_);
  and (_12789_, _12788_, _07104_);
  and (_12790_, _12789_, _12785_);
  or (_12791_, _12790_, _12712_);
  and (_12792_, _12791_, _03095_);
  or (_12793_, _12709_, _05086_);
  and (_12794_, _12723_, _03094_);
  and (_12795_, _12714_, _02991_);
  or (_12796_, _12795_, _12794_);
  and (_12797_, _12796_, _12793_);
  or (_12798_, _12797_, _02994_);
  or (_12799_, _12798_, _12792_);
  nor (_12800_, _10935_, _06175_);
  or (_12801_, _12709_, _07120_);
  or (_12802_, _12801_, _12800_);
  and (_12803_, _12802_, _07118_);
  and (_12804_, _12803_, _12799_);
  nor (_12805_, _10941_, _06175_);
  or (_12806_, _12805_, _12709_);
  and (_12807_, _12806_, _03099_);
  or (_12808_, _12807_, _03133_);
  or (_12809_, _12808_, _12804_);
  or (_12810_, _12720_, _03138_);
  and (_12811_, _12810_, _03142_);
  and (_12812_, _12811_, _12809_);
  and (_12813_, _12742_, _02778_);
  or (_12814_, _12813_, _02852_);
  or (_12815_, _12814_, _12812_);
  and (_12816_, _10988_, _04661_);
  or (_12817_, _12709_, _02853_);
  or (_12818_, _12817_, _12816_);
  and (_12819_, _12818_, _34446_);
  and (_12820_, _12819_, _12815_);
  or (_12821_, _12820_, _12708_);
  and (_35615_[2], _12821_, _35583_);
  nor (_12822_, _34446_, _06754_);
  nor (_12823_, _04661_, _06754_);
  and (_12824_, _11134_, _04661_);
  or (_12825_, _12824_, _12823_);
  and (_12826_, _12825_, _03107_);
  and (_12827_, _04661_, _05616_);
  or (_12828_, _12827_, _12823_);
  or (_12829_, _12828_, _05261_);
  nor (_12830_, _06175_, _04226_);
  or (_12831_, _12830_, _12823_);
  or (_12832_, _12831_, _03860_);
  nor (_12833_, _11014_, _06175_);
  or (_12834_, _12833_, _12823_);
  or (_12835_, _12834_, _06162_);
  and (_12836_, _04661_, \oc8051_golden_model_1.ACC [3]);
  or (_12837_, _12836_, _12823_);
  and (_12838_, _12837_, _02837_);
  nor (_12839_, _02837_, _06754_);
  or (_12840_, _12839_, _02932_);
  or (_12841_, _12840_, _12838_);
  and (_12842_, _12841_, _02939_);
  and (_12843_, _12842_, _12835_);
  and (_12844_, _12831_, _02930_);
  nor (_12845_, _05286_, _06754_);
  and (_12846_, _11011_, _05286_);
  or (_12847_, _12846_, _12845_);
  and (_12848_, _12847_, _02799_);
  or (_12849_, _12848_, _12844_);
  or (_12850_, _12849_, _02928_);
  or (_12851_, _12850_, _12843_);
  or (_12852_, _12837_, _02943_);
  and (_12853_, _12852_, _12851_);
  or (_12854_, _12853_, _02796_);
  and (_12855_, _11009_, _05286_);
  or (_12856_, _12855_, _12845_);
  or (_12857_, _12856_, _02927_);
  and (_12858_, _12857_, _06189_);
  and (_12859_, _12858_, _12854_);
  and (_12860_, _12846_, _11040_);
  or (_12861_, _12860_, _12845_);
  and (_12862_, _12861_, _02790_);
  or (_12863_, _12862_, _06195_);
  or (_12864_, _12863_, _12859_);
  nor (_12865_, _06684_, _06520_);
  nor (_12866_, _12865_, _06685_);
  or (_12867_, _12866_, _06201_);
  and (_12868_, _12867_, _02966_);
  and (_12869_, _12868_, _12864_);
  nor (_12870_, _11058_, _06716_);
  or (_12871_, _12870_, _12845_);
  and (_12872_, _12871_, _02785_);
  or (_12873_, _12872_, _03861_);
  or (_12874_, _12873_, _12869_);
  and (_12875_, _12874_, _12832_);
  or (_12876_, _12875_, _03850_);
  and (_12877_, _06116_, _04661_);
  or (_12878_, _12823_, _06726_);
  or (_12879_, _12878_, _12877_);
  and (_12880_, _12879_, _12876_);
  or (_12881_, _12880_, _02524_);
  nor (_12882_, _11114_, _06175_);
  or (_12883_, _12823_, _02970_);
  or (_12884_, _12883_, _12882_);
  and (_12885_, _12884_, _06737_);
  and (_12886_, _12885_, _12881_);
  nand (_12887_, _07086_, _07014_);
  nor (_12888_, _12776_, _07025_);
  nor (_12889_, _12888_, _07017_);
  and (_12890_, _12888_, _07017_);
  or (_12891_, _12890_, _12889_);
  or (_12892_, _12891_, _07086_);
  and (_12893_, _12892_, _06731_);
  and (_12894_, _12893_, _12887_);
  or (_12895_, _12894_, _02974_);
  or (_12896_, _12895_, _12886_);
  and (_12897_, _12896_, _12829_);
  or (_12898_, _12897_, _02977_);
  and (_12899_, _11128_, _04661_);
  or (_12900_, _12823_, _07092_);
  or (_12901_, _12900_, _12899_);
  and (_12902_, _12901_, _07104_);
  and (_12903_, _12902_, _12898_);
  or (_12904_, _12903_, _12826_);
  and (_12905_, _12904_, _03095_);
  or (_12906_, _12823_, _04939_);
  and (_12907_, _12837_, _03094_);
  and (_12908_, _12828_, _02991_);
  or (_12909_, _12908_, _12907_);
  and (_12910_, _12909_, _12906_);
  or (_12911_, _12910_, _02994_);
  or (_12912_, _12911_, _12905_);
  nor (_12913_, _11127_, _06175_);
  or (_12914_, _12823_, _07120_);
  or (_12915_, _12914_, _12913_);
  and (_12916_, _12915_, _07118_);
  and (_12917_, _12916_, _12912_);
  nor (_12918_, _11133_, _06175_);
  or (_12919_, _12918_, _12823_);
  and (_12920_, _12919_, _03099_);
  or (_12921_, _12920_, _03133_);
  or (_12922_, _12921_, _12917_);
  or (_12923_, _12834_, _03138_);
  and (_12924_, _12923_, _03142_);
  and (_12925_, _12924_, _12922_);
  and (_12926_, _12856_, _02778_);
  or (_12927_, _12926_, _02852_);
  or (_12928_, _12927_, _12925_);
  and (_12929_, _11185_, _04661_);
  or (_12930_, _12823_, _02853_);
  or (_12931_, _12930_, _12929_);
  and (_12932_, _12931_, _34446_);
  and (_12933_, _12932_, _12928_);
  or (_12934_, _12933_, _12822_);
  and (_35615_[3], _12934_, _35583_);
  nor (_12935_, _34446_, _06755_);
  nor (_12936_, _04661_, _06755_);
  and (_12937_, _11333_, _04661_);
  or (_12938_, _12937_, _12936_);
  and (_12939_, _12938_, _03107_);
  and (_12940_, _05629_, _04661_);
  or (_12941_, _12940_, _12936_);
  or (_12942_, _12941_, _05261_);
  nor (_12943_, _11313_, _06175_);
  or (_12944_, _12943_, _12936_);
  and (_12945_, _12944_, _02524_);
  nor (_12946_, _05143_, _06175_);
  or (_12947_, _12946_, _12936_);
  or (_12948_, _12947_, _03860_);
  nor (_12949_, _11207_, _06175_);
  or (_12950_, _12949_, _12936_);
  or (_12951_, _12950_, _06162_);
  and (_12952_, _04661_, \oc8051_golden_model_1.ACC [4]);
  or (_12953_, _12952_, _12936_);
  and (_12954_, _12953_, _02837_);
  nor (_12955_, _02837_, _06755_);
  or (_12956_, _12955_, _02932_);
  or (_12957_, _12956_, _12954_);
  and (_12958_, _12957_, _02939_);
  and (_12959_, _12958_, _12951_);
  and (_12960_, _12947_, _02930_);
  nor (_12961_, _05286_, _06755_);
  and (_12962_, _11224_, _05286_);
  or (_12963_, _12962_, _12961_);
  and (_12964_, _12963_, _02799_);
  or (_12965_, _12964_, _12960_);
  or (_12966_, _12965_, _02928_);
  or (_12967_, _12966_, _12959_);
  or (_12968_, _12953_, _02943_);
  and (_12969_, _12968_, _12967_);
  or (_12970_, _12969_, _02796_);
  and (_12971_, _11203_, _05286_);
  or (_12972_, _12971_, _12961_);
  or (_12973_, _12972_, _02927_);
  and (_12974_, _12973_, _06189_);
  and (_12975_, _12974_, _12970_);
  or (_12976_, _12961_, _11239_);
  and (_12977_, _12976_, _02790_);
  and (_12978_, _12977_, _12963_);
  or (_12979_, _12978_, _06195_);
  or (_12980_, _12979_, _12975_);
  nor (_12981_, _06689_, _06687_);
  nor (_12982_, _12981_, _06690_);
  or (_12983_, _12982_, _06201_);
  and (_12984_, _12983_, _02966_);
  and (_12985_, _12984_, _12980_);
  nor (_12986_, _11257_, _06716_);
  or (_12987_, _12986_, _12961_);
  and (_12988_, _12987_, _02785_);
  or (_12989_, _12988_, _03861_);
  or (_12990_, _12989_, _12985_);
  and (_12991_, _12990_, _12948_);
  or (_12992_, _12991_, _03850_);
  and (_12993_, _06121_, _04661_);
  or (_12994_, _12936_, _06726_);
  or (_12995_, _12994_, _12993_);
  and (_12996_, _12995_, _02970_);
  and (_12997_, _12996_, _12992_);
  or (_12998_, _12997_, _12945_);
  and (_12999_, _12998_, _06737_);
  not (_13000_, _07086_);
  or (_13001_, _13000_, _07049_);
  nor (_13002_, _12888_, _07016_);
  or (_13003_, _13002_, _07015_);
  nand (_13004_, _13003_, _07052_);
  or (_13005_, _13003_, _07052_);
  and (_13006_, _13005_, _13004_);
  or (_13007_, _13006_, _07086_);
  and (_13008_, _13007_, _06731_);
  and (_13009_, _13008_, _13001_);
  or (_13010_, _13009_, _02974_);
  or (_13011_, _13010_, _12999_);
  and (_13012_, _13011_, _12942_);
  or (_13013_, _13012_, _02977_);
  and (_13014_, _11327_, _04661_);
  or (_13015_, _12936_, _07092_);
  or (_13016_, _13015_, _13014_);
  and (_13017_, _13016_, _07104_);
  and (_13018_, _13017_, _13013_);
  or (_13019_, _13018_, _12939_);
  and (_13020_, _13019_, _03095_);
  or (_13021_, _12936_, _05190_);
  and (_13022_, _12953_, _03094_);
  and (_13023_, _12941_, _02991_);
  or (_13024_, _13023_, _13022_);
  and (_13025_, _13024_, _13021_);
  or (_13026_, _13025_, _02994_);
  or (_13027_, _13026_, _13020_);
  nor (_13028_, _11326_, _06175_);
  or (_13029_, _12936_, _07120_);
  or (_13030_, _13029_, _13028_);
  and (_13031_, _13030_, _07118_);
  and (_13032_, _13031_, _13027_);
  nor (_13033_, _11332_, _06175_);
  or (_13034_, _13033_, _12936_);
  and (_13035_, _13034_, _03099_);
  or (_13036_, _13035_, _03133_);
  or (_13037_, _13036_, _13032_);
  or (_13038_, _12950_, _03138_);
  and (_13039_, _13038_, _03142_);
  and (_13040_, _13039_, _13037_);
  and (_13041_, _12972_, _02778_);
  or (_13042_, _13041_, _02852_);
  or (_13043_, _13042_, _13040_);
  and (_13044_, _11383_, _04661_);
  or (_13045_, _12936_, _02853_);
  or (_13046_, _13045_, _13044_);
  and (_13047_, _13046_, _34446_);
  and (_13048_, _13047_, _13043_);
  or (_13049_, _13048_, _12935_);
  and (_35615_[4], _13049_, _35583_);
  nor (_13050_, _34446_, _06756_);
  nor (_13051_, _04661_, _06756_);
  and (_13052_, _11531_, _04661_);
  or (_13053_, _13052_, _13051_);
  and (_13054_, _13053_, _03107_);
  and (_13055_, _05633_, _04661_);
  or (_13056_, _13055_, _13051_);
  or (_13057_, _13056_, _05261_);
  nor (_13058_, _11511_, _06175_);
  or (_13059_, _13058_, _13051_);
  and (_13060_, _13059_, _02524_);
  nor (_13061_, _11408_, _06175_);
  or (_13062_, _13061_, _13051_);
  or (_13063_, _13062_, _06162_);
  and (_13064_, _04661_, \oc8051_golden_model_1.ACC [5]);
  or (_13065_, _13064_, _13051_);
  and (_13066_, _13065_, _02837_);
  nor (_13067_, _02837_, _06756_);
  or (_13068_, _13067_, _02932_);
  or (_13069_, _13068_, _13066_);
  and (_13070_, _13069_, _02939_);
  and (_13071_, _13070_, _13063_);
  nor (_13072_, _04839_, _06175_);
  or (_13073_, _13072_, _13051_);
  and (_13074_, _13073_, _02930_);
  nor (_13075_, _05286_, _06756_);
  and (_13076_, _11422_, _05286_);
  or (_13077_, _13076_, _13075_);
  and (_13078_, _13077_, _02799_);
  or (_13079_, _13078_, _13074_);
  or (_13080_, _13079_, _02928_);
  or (_13081_, _13080_, _13071_);
  or (_13082_, _13065_, _02943_);
  and (_13083_, _13082_, _13081_);
  or (_13084_, _13083_, _02796_);
  and (_13085_, _11405_, _05286_);
  or (_13086_, _13085_, _13075_);
  or (_13087_, _13086_, _02927_);
  and (_13088_, _13087_, _06189_);
  and (_13089_, _13088_, _13084_);
  or (_13090_, _13075_, _11437_);
  and (_13091_, _13077_, _02790_);
  and (_13092_, _13091_, _13090_);
  or (_13093_, _13092_, _06195_);
  or (_13094_, _13093_, _13089_);
  nor (_13095_, _06692_, _06394_);
  nor (_13096_, _13095_, _06693_);
  or (_13097_, _13096_, _06201_);
  and (_13098_, _13097_, _02966_);
  and (_13099_, _13098_, _13094_);
  nor (_13100_, _11455_, _06716_);
  or (_13101_, _13100_, _13075_);
  and (_13102_, _13101_, _02785_);
  or (_13103_, _13102_, _03861_);
  or (_13104_, _13103_, _13099_);
  or (_13105_, _13073_, _03860_);
  and (_13106_, _13105_, _13104_);
  or (_13107_, _13106_, _03850_);
  and (_13108_, _06120_, _04661_);
  or (_13109_, _13051_, _06726_);
  or (_13110_, _13109_, _13108_);
  and (_13111_, _13110_, _02970_);
  and (_13112_, _13111_, _13107_);
  or (_13113_, _13112_, _13060_);
  and (_13114_, _13113_, _06737_);
  nand (_13115_, _07086_, _07059_);
  not (_13116_, _07051_);
  and (_13117_, _13004_, _13116_);
  nor (_13118_, _13117_, _07062_);
  and (_13119_, _13117_, _07062_);
  or (_13120_, _13119_, _13118_);
  or (_13121_, _13120_, _07086_);
  and (_13122_, _13121_, _06731_);
  and (_13123_, _13122_, _13115_);
  or (_13124_, _13123_, _02974_);
  or (_13125_, _13124_, _13114_);
  and (_13126_, _13125_, _13057_);
  or (_13127_, _13126_, _02977_);
  and (_13128_, _11525_, _04661_);
  or (_13129_, _13051_, _07092_);
  or (_13130_, _13129_, _13128_);
  and (_13131_, _13130_, _07104_);
  and (_13132_, _13131_, _13127_);
  or (_13133_, _13132_, _13054_);
  and (_13134_, _13133_, _03095_);
  or (_13135_, _13051_, _04890_);
  and (_13136_, _13065_, _03094_);
  and (_13137_, _13056_, _02991_);
  or (_13138_, _13137_, _13136_);
  and (_13139_, _13138_, _13135_);
  or (_13140_, _13139_, _02994_);
  or (_13141_, _13140_, _13134_);
  nor (_13142_, _11524_, _06175_);
  or (_13143_, _13051_, _07120_);
  or (_13144_, _13143_, _13142_);
  and (_13145_, _13144_, _07118_);
  and (_13146_, _13145_, _13141_);
  nor (_13147_, _11530_, _06175_);
  or (_13148_, _13147_, _13051_);
  and (_13149_, _13148_, _03099_);
  or (_13150_, _13149_, _03133_);
  or (_13151_, _13150_, _13146_);
  or (_13152_, _13062_, _03138_);
  and (_13153_, _13152_, _03142_);
  and (_13154_, _13153_, _13151_);
  and (_13155_, _13086_, _02778_);
  or (_13156_, _13155_, _02852_);
  or (_13157_, _13156_, _13154_);
  and (_13158_, _11580_, _04661_);
  or (_13159_, _13051_, _02853_);
  or (_13160_, _13159_, _13158_);
  and (_13161_, _13160_, _34446_);
  and (_13162_, _13161_, _13157_);
  or (_13163_, _13162_, _13050_);
  and (_35615_[5], _13163_, _35583_);
  nor (_13164_, _34446_, _06997_);
  nor (_13165_, _04661_, _06997_);
  and (_13166_, _11601_, _04661_);
  or (_13167_, _13166_, _13165_);
  and (_13168_, _13167_, _03107_);
  and (_13169_, _11718_, _04661_);
  or (_13170_, _13169_, _13165_);
  or (_13171_, _13170_, _05261_);
  nor (_13172_, _04735_, _06175_);
  or (_13173_, _13172_, _13165_);
  or (_13174_, _13173_, _03860_);
  nor (_13175_, _11610_, _06175_);
  or (_13176_, _13175_, _13165_);
  or (_13177_, _13176_, _06162_);
  and (_13178_, _04661_, \oc8051_golden_model_1.ACC [6]);
  or (_13179_, _13178_, _13165_);
  and (_13180_, _13179_, _02837_);
  nor (_13181_, _02837_, _06997_);
  or (_13182_, _13181_, _02932_);
  or (_13183_, _13182_, _13180_);
  and (_13184_, _13183_, _02939_);
  and (_13185_, _13184_, _13177_);
  and (_13186_, _13173_, _02930_);
  nor (_13187_, _05286_, _06997_);
  and (_13188_, _11604_, _05286_);
  or (_13189_, _13188_, _13187_);
  and (_13190_, _13189_, _02799_);
  or (_13191_, _13190_, _13186_);
  or (_13192_, _13191_, _02928_);
  or (_13193_, _13192_, _13185_);
  or (_13194_, _13179_, _02943_);
  and (_13195_, _13194_, _13193_);
  or (_13196_, _13195_, _02796_);
  and (_13197_, _11633_, _05286_);
  or (_13198_, _13197_, _13187_);
  or (_13199_, _13198_, _02927_);
  and (_13200_, _13199_, _06189_);
  and (_13201_, _13200_, _13196_);
  or (_13202_, _13187_, _11603_);
  and (_13203_, _13189_, _02790_);
  and (_13204_, _13203_, _13202_);
  or (_13205_, _13204_, _06195_);
  or (_13206_, _13205_, _13201_);
  nor (_13207_, _06708_, _06695_);
  nor (_13208_, _13207_, _06709_);
  or (_13209_, _13208_, _06201_);
  and (_13210_, _13209_, _02966_);
  and (_13211_, _13210_, _13206_);
  nor (_13212_, _11655_, _06716_);
  or (_13213_, _13212_, _13187_);
  and (_13214_, _13213_, _02785_);
  or (_13215_, _13214_, _03861_);
  or (_13216_, _13215_, _13211_);
  and (_13217_, _13216_, _13174_);
  or (_13218_, _13217_, _03850_);
  and (_13219_, _05798_, _04661_);
  or (_13220_, _13165_, _06726_);
  or (_13221_, _13220_, _13219_);
  and (_13222_, _13221_, _13218_);
  or (_13223_, _13222_, _02524_);
  nor (_13224_, _11711_, _06175_);
  or (_13225_, _13165_, _02970_);
  or (_13226_, _13225_, _13224_);
  and (_13227_, _13226_, _06737_);
  and (_13228_, _13227_, _13223_);
  nor (_13229_, _13117_, _07060_);
  or (_13230_, _13229_, _07061_);
  and (_13231_, _13230_, _07066_);
  nor (_13232_, _13230_, _07066_);
  or (_13233_, _13232_, _13231_);
  or (_13234_, _13233_, _07086_);
  or (_13235_, _13000_, _07003_);
  and (_13236_, _13235_, _06731_);
  and (_13237_, _13236_, _13234_);
  or (_13238_, _13237_, _02974_);
  or (_13239_, _13238_, _13228_);
  and (_13240_, _13239_, _13171_);
  or (_13241_, _13240_, _02977_);
  and (_13242_, _11728_, _04661_);
  or (_13243_, _13165_, _07092_);
  or (_13244_, _13243_, _13242_);
  and (_13245_, _13244_, _07104_);
  and (_13246_, _13245_, _13241_);
  or (_13247_, _13246_, _13168_);
  and (_13248_, _13247_, _03095_);
  or (_13249_, _13165_, _04784_);
  and (_13250_, _13179_, _03094_);
  and (_13251_, _13170_, _02991_);
  or (_13252_, _13251_, _13250_);
  and (_13253_, _13252_, _13249_);
  or (_13254_, _13253_, _02994_);
  or (_13255_, _13254_, _13248_);
  nor (_13256_, _11726_, _06175_);
  or (_13257_, _13165_, _07120_);
  or (_13258_, _13257_, _13256_);
  and (_13259_, _13258_, _07118_);
  and (_13260_, _13259_, _13255_);
  nor (_13261_, _11600_, _06175_);
  or (_13262_, _13261_, _13165_);
  and (_13263_, _13262_, _03099_);
  or (_13264_, _13263_, _03133_);
  or (_13265_, _13264_, _13260_);
  or (_13266_, _13176_, _03138_);
  and (_13267_, _13266_, _03142_);
  and (_13268_, _13267_, _13265_);
  and (_13269_, _13198_, _02778_);
  or (_13270_, _13269_, _02852_);
  or (_13271_, _13270_, _13268_);
  and (_13272_, _11778_, _04661_);
  or (_13273_, _13165_, _02853_);
  or (_13274_, _13273_, _13272_);
  and (_13275_, _13274_, _34446_);
  and (_13276_, _13275_, _13271_);
  or (_13277_, _13276_, _13164_);
  and (_35615_[6], _13277_, _35583_);
  nor (_13278_, _34446_, _02658_);
  and (_13279_, _08143_, \oc8051_golden_model_1.ACC [1]);
  nand (_13280_, _07143_, _05719_);
  nand (_13281_, _07684_, _02856_);
  and (_13282_, _13281_, _08074_);
  not (_13283_, _03541_);
  and (_13284_, _10346_, _02574_);
  not (_13285_, _07193_);
  and (_13286_, _03823_, _02658_);
  nor (_13287_, _13286_, _07218_);
  and (_13288_, _13287_, _13285_);
  nand (_13289_, _07946_, _07759_);
  nand (_13290_, _07899_, _08829_);
  nand (_13291_, _13286_, _07317_);
  or (_13292_, _07167_, _07876_);
  nor (_13293_, _04654_, _02658_);
  and (_13294_, _10427_, _04654_);
  nor (_13295_, _13294_, _13293_);
  nand (_13296_, _13295_, _02977_);
  nor (_13297_, _07808_, _02835_);
  and (_13298_, _04654_, _03805_);
  nor (_13299_, _13298_, _13293_);
  nand (_13300_, _13299_, _03861_);
  and (_13301_, _03495_, _02782_);
  nor (_13302_, _03680_, _02912_);
  nor (_13303_, _13302_, _02498_);
  nor (_13304_, _13303_, _03268_);
  or (_13305_, _07475_, _03805_);
  nor (_13306_, _05291_, _02658_);
  and (_13307_, _10441_, _05291_);
  nor (_13308_, _13307_, _13306_);
  nand (_13309_, _13308_, _02799_);
  and (_13310_, _13309_, _03693_);
  nor (_13311_, _07651_, _07406_);
  or (_13312_, _06114_, _07408_);
  or (_13313_, _07413_, _03805_);
  or (_13314_, _07415_, _02658_);
  nand (_13315_, _07415_, _02658_);
  and (_13316_, _13315_, _13314_);
  nand (_13317_, _13316_, _09158_);
  and (_13318_, _13317_, _13313_);
  and (_13319_, _13318_, _07406_);
  and (_13320_, _13319_, _13312_);
  or (_13321_, _13320_, _13311_);
  and (_13322_, _13321_, _07429_);
  and (_13323_, _07434_, \oc8051_golden_model_1.XRAM_DATA_IN [0]);
  or (_13324_, _13323_, _03806_);
  or (_13325_, _13324_, _13322_);
  or (_13326_, _06114_, _05311_);
  and (_13327_, _13326_, _06162_);
  and (_13328_, _13327_, _13325_);
  nor (_13329_, _05036_, _07325_);
  nor (_13330_, _13329_, _13293_);
  nor (_13331_, _13330_, _06162_);
  or (_13332_, _13331_, _02799_);
  or (_13333_, _13332_, _13328_);
  and (_13334_, _13333_, _13310_);
  nor (_13335_, _13299_, _03693_);
  or (_13336_, _13335_, _07476_);
  or (_13337_, _13336_, _13334_);
  and (_13338_, _13337_, _13305_);
  or (_13339_, _13338_, _03374_);
  or (_13340_, _06114_, _03375_);
  and (_13341_, _13340_, _02943_);
  and (_13342_, _13341_, _13339_);
  nor (_13343_, _07651_, _02943_);
  or (_13344_, _13343_, _07486_);
  or (_13345_, _13344_, _13342_);
  nand (_13346_, _07486_, _06814_);
  and (_13347_, _13346_, _13345_);
  or (_13348_, _13347_, _02796_);
  or (_13349_, _13293_, _02927_);
  and (_13350_, _13349_, _06189_);
  and (_13351_, _13350_, _13348_);
  nor (_13352_, _13330_, _06189_);
  or (_13353_, _13352_, _06195_);
  nor (_13354_, _13353_, _13351_);
  not (_13355_, _06656_);
  and (_13356_, _13355_, _06195_);
  or (_13357_, _13356_, _13354_);
  nand (_13358_, _13357_, _13304_);
  not (_13359_, _07524_);
  or (_13360_, _13359_, _13304_);
  and (_13361_, _13360_, _13358_);
  or (_13362_, _13361_, _13301_);
  nand (_13363_, _07524_, _13301_);
  and (_13364_, _13363_, _07330_);
  and (_13365_, _13364_, _13362_);
  nor (_13366_, _07381_, _02658_);
  nor (_13367_, _13366_, _07382_);
  nor (_13368_, _13367_, _07330_);
  or (_13369_, _13368_, _02898_);
  or (_13370_, _13369_, _13365_);
  nor (_13371_, _08006_, _02658_);
  nor (_13372_, _13371_, _10016_);
  nand (_13373_, _13372_, _02898_);
  and (_13374_, _13373_, _13370_);
  or (_13375_, _13374_, _07540_);
  nand (_13376_, _07759_, _07540_);
  and (_13377_, _13376_, _13375_);
  or (_13378_, _13377_, _07700_);
  nand (_13379_, _02835_, _07700_);
  and (_13380_, _13379_, _02966_);
  and (_13381_, _13380_, _13378_);
  nor (_13382_, _10473_, _07786_);
  nor (_13383_, _13382_, _13306_);
  nor (_13384_, _13383_, _02966_);
  or (_13385_, _13384_, _03861_);
  or (_13386_, _13385_, _13381_);
  and (_13387_, _13386_, _13300_);
  or (_13388_, _13387_, _03850_);
  and (_13389_, _06114_, _04654_);
  nor (_13390_, _13389_, _13293_);
  nand (_13391_, _13390_, _03850_);
  and (_13392_, _13391_, _02970_);
  and (_13393_, _13392_, _13388_);
  nor (_13394_, _10530_, _07325_);
  nor (_13395_, _13394_, _13293_);
  nor (_13396_, _13395_, _02970_);
  or (_13397_, _13396_, _06731_);
  or (_13398_, _13397_, _13393_);
  nand (_13399_, _07086_, _06731_);
  and (_13400_, _13399_, _13398_);
  and (_13401_, _13400_, _02552_);
  nor (_13402_, _02835_, _02552_);
  or (_13403_, _13402_, _02974_);
  or (_13404_, _13403_, _13401_);
  and (_13405_, _04654_, _05647_);
  nor (_13406_, _13405_, _13293_);
  nand (_13407_, _13406_, _02974_);
  and (_13408_, _13407_, _07808_);
  and (_13409_, _13408_, _13404_);
  or (_13410_, _13409_, _13297_);
  and (_13411_, _07822_, _07816_);
  and (_13412_, _13411_, _13410_);
  not (_13413_, _13411_);
  and (_13414_, _13413_, _13287_);
  or (_13415_, _13414_, _07829_);
  or (_13416_, _13415_, _13412_);
  and (_13417_, _10346_, _02581_);
  not (_13418_, _13417_);
  or (_13419_, _07828_, _13287_);
  and (_13420_, _13419_, _13418_);
  and (_13421_, _13420_, _13416_);
  and (_13422_, _05889_, _02658_);
  nor (_13423_, _13422_, _07167_);
  and (_13424_, _13417_, _13423_);
  or (_13425_, _13424_, _13421_);
  and (_13426_, _13425_, _03487_);
  and (_13427_, _13423_, _03486_);
  or (_13428_, _13427_, _03105_);
  or (_13429_, _13428_, _13426_);
  or (_13430_, _10546_, _03106_);
  and (_13431_, _13430_, _07846_);
  and (_13432_, _13431_, _13429_);
  and (_13433_, _07319_, _08830_);
  or (_13434_, _13433_, _02977_);
  or (_13435_, _13434_, _13432_);
  and (_13436_, _13435_, _13296_);
  or (_13437_, _13436_, _03107_);
  or (_13438_, _13293_, _07104_);
  and (_13439_, _13438_, _07868_);
  and (_13440_, _13439_, _13437_);
  or (_13441_, _07218_, _03499_);
  and (_13442_, _13441_, _09406_);
  or (_13443_, _13442_, _13440_);
  and (_13444_, _13443_, _13292_);
  or (_13445_, _13444_, _03092_);
  or (_13446_, _10545_, _03093_);
  and (_13447_, _13446_, _07886_);
  and (_13448_, _13447_, _13445_);
  and (_13449_, _07880_, _08117_);
  or (_13450_, _13449_, _13448_);
  and (_13451_, _13450_, _03881_);
  nor (_13452_, _13406_, _13329_);
  and (_13453_, _13452_, _02991_);
  or (_13454_, _13453_, _07317_);
  or (_13455_, _13454_, _13451_);
  and (_13456_, _13455_, _13291_);
  or (_13457_, _13456_, _07315_);
  nand (_13458_, _13422_, _07315_);
  and (_13459_, _13458_, _03098_);
  and (_13460_, _13459_, _13457_);
  nand (_13461_, _10423_, _07902_);
  and (_13462_, _13461_, _07901_);
  or (_13463_, _13462_, _13460_);
  and (_13464_, _13463_, _13290_);
  or (_13465_, _13464_, _02994_);
  nor (_13466_, _10425_, _07325_);
  nor (_13467_, _13466_, _13293_);
  nand (_13468_, _13467_, _02994_);
  and (_13469_, _13468_, _07241_);
  and (_13470_, _13469_, _13465_);
  nor (_13471_, _07241_, _07524_);
  or (_13472_, _13471_, _07236_);
  or (_13473_, _13472_, _13470_);
  nand (_13474_, _13367_, _07236_);
  and (_13475_, _13474_, _03104_);
  and (_13476_, _13475_, _13473_);
  nand (_13477_, _08029_, _13372_);
  and (_13478_, _13477_, _07948_);
  or (_13479_, _13478_, _13476_);
  and (_13480_, _13479_, _13289_);
  or (_13481_, _13480_, _08027_);
  nand (_13482_, _08027_, _07294_);
  and (_13483_, _13482_, _07193_);
  and (_13484_, _13483_, _13481_);
  nor (_13485_, _13484_, _13288_);
  nor (_13486_, _13485_, _13284_);
  and (_13487_, _13423_, _13284_);
  or (_13488_, _13487_, _13486_);
  and (_13489_, _13488_, _13283_);
  and (_13490_, _13423_, _03541_);
  or (_13491_, _13490_, _03124_);
  or (_13492_, _13491_, _13489_);
  and (_13493_, _13492_, _13282_);
  and (_13494_, _08073_, _08830_);
  or (_13495_, _13494_, _07143_);
  or (_13496_, _13495_, _13493_);
  and (_13497_, _13496_, _13280_);
  or (_13498_, _13497_, _03133_);
  nand (_13499_, _13330_, _03133_);
  and (_13500_, _13499_, _08139_);
  and (_13501_, _13500_, _13498_);
  and (_13502_, _08138_, _02658_);
  or (_13503_, _13502_, _13501_);
  and (_13504_, _13503_, _09716_);
  or (_13505_, _13504_, _13279_);
  and (_13506_, _13505_, _03142_);
  and (_13507_, _13293_, _02778_);
  or (_13508_, _13507_, _02852_);
  or (_13509_, _13508_, _13506_);
  nand (_13510_, _13330_, _02852_);
  and (_13511_, _13510_, _08161_);
  and (_13512_, _13511_, _13509_);
  nor (_13513_, _08167_, _02658_);
  nor (_13514_, _13513_, _09696_);
  or (_13515_, _13514_, _13512_);
  nand (_13516_, _08167_, _02477_);
  and (_13517_, _13516_, _34446_);
  and (_13518_, _13517_, _13515_);
  or (_13519_, _13518_, _13278_);
  and (_35614_[0], _13519_, _35583_);
  nor (_13520_, _34446_, _02477_);
  nand (_13521_, _07143_, _02658_);
  and (_13522_, _07927_, _07925_);
  nor (_13523_, _13522_, _07928_);
  or (_13524_, _13523_, _07917_);
  nand (_13525_, _07899_, _07760_);
  nand (_13526_, _07216_, _03242_);
  and (_13527_, _07869_, _07215_);
  nor (_13528_, _04654_, _02477_);
  and (_13529_, _10614_, _04654_);
  nor (_13530_, _13529_, _13528_);
  nand (_13531_, _13530_, _02977_);
  nor (_13532_, _07808_, _03742_);
  nor (_13533_, _07325_, _03989_);
  nor (_13534_, _13533_, _13528_);
  nand (_13535_, _13534_, _03861_);
  nor (_13536_, _07651_, _07764_);
  nor (_13537_, _13536_, _07763_);
  and (_13538_, _13537_, _07682_);
  nor (_13539_, _13537_, _07682_);
  or (_13540_, _13539_, _13538_);
  nand (_13541_, _13540_, _02898_);
  and (_13542_, _13541_, _07541_);
  nor (_13543_, _07638_, _07406_);
  or (_13544_, _06113_, _07408_);
  nor (_13545_, _07413_, _03989_);
  or (_13546_, _07415_, \oc8051_golden_model_1.ACC [1]);
  nand (_13547_, _07415_, \oc8051_golden_model_1.ACC [1]);
  and (_13548_, _13547_, _13546_);
  and (_13549_, _13548_, _07413_);
  or (_13550_, _13549_, _03343_);
  or (_13551_, _13550_, _13545_);
  and (_13552_, _13551_, _07406_);
  and (_13553_, _13552_, _13544_);
  or (_13554_, _13553_, _13543_);
  and (_13555_, _13554_, _07429_);
  and (_13556_, _07434_, \oc8051_golden_model_1.XRAM_DATA_IN [1]);
  or (_13557_, _13556_, _03806_);
  or (_13558_, _13557_, _13555_);
  or (_13559_, _06113_, _05311_);
  and (_13560_, _13559_, _06162_);
  and (_13561_, _13560_, _13558_);
  nor (_13562_, _04654_, \oc8051_golden_model_1.ACC [1]);
  and (_13563_, _10622_, _04654_);
  nor (_13564_, _13563_, _13562_);
  and (_13565_, _13564_, _02932_);
  or (_13566_, _13565_, _07402_);
  or (_13567_, _13566_, _13561_);
  nor (_13568_, _07441_, \oc8051_golden_model_1.PSW [6]);
  nor (_13569_, _13568_, \oc8051_golden_model_1.ACC [1]);
  and (_13570_, _13568_, \oc8051_golden_model_1.ACC [1]);
  nor (_13571_, _13570_, _13569_);
  nand (_13572_, _13571_, _07402_);
  and (_13573_, _13572_, _02939_);
  and (_13574_, _13573_, _13567_);
  nor (_13575_, _05291_, _02477_);
  and (_13576_, _10617_, _05291_);
  nor (_13577_, _13576_, _13575_);
  nor (_13578_, _13577_, _03186_);
  nor (_13579_, _13534_, _03693_);
  or (_13580_, _13579_, _07476_);
  or (_13581_, _13580_, _13578_);
  or (_13582_, _13581_, _13574_);
  nand (_13583_, _07476_, _03989_);
  and (_13584_, _13583_, _13582_);
  or (_13585_, _13584_, _03374_);
  or (_13586_, _06113_, _03375_);
  and (_13587_, _13586_, _02943_);
  and (_13588_, _13587_, _13585_);
  nor (_13589_, _07638_, _02943_);
  or (_13590_, _13589_, _07486_);
  or (_13591_, _13590_, _13588_);
  nand (_13592_, _07486_, _06808_);
  and (_13593_, _13592_, _13591_);
  or (_13594_, _13593_, _02796_);
  and (_13595_, _10620_, _05291_);
  nor (_13596_, _13595_, _13575_);
  nand (_13597_, _13596_, _02796_);
  and (_13598_, _13597_, _06189_);
  and (_13599_, _13598_, _13594_);
  and (_13600_, _13576_, _10616_);
  nor (_13601_, _13600_, _13575_);
  nor (_13602_, _13601_, _06189_);
  or (_13603_, _13602_, _06195_);
  or (_13604_, _13603_, _13599_);
  and (_13605_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  nor (_13606_, _13605_, _07029_);
  nor (_13607_, _13606_, _06657_);
  or (_13608_, _13607_, _06201_);
  and (_13609_, _13608_, _13604_);
  or (_13610_, _13609_, _07401_);
  not (_13611_, _07764_);
  and (_13612_, _13611_, _03805_);
  nor (_13613_, _13612_, _07763_);
  and (_13614_, _13613_, _07217_);
  nor (_13615_, _13613_, _07217_);
  or (_13616_, _13615_, _13614_);
  or (_13617_, _13616_, _07400_);
  and (_13618_, _13617_, _07330_);
  and (_13619_, _13618_, _13610_);
  and (_13620_, _13611_, _06114_);
  nor (_13621_, _13620_, _07763_);
  and (_13622_, _13621_, _07166_);
  nor (_13623_, _13621_, _07166_);
  or (_13624_, _13623_, _13622_);
  and (_13625_, _13624_, _07329_);
  or (_13626_, _13625_, _02898_);
  or (_13627_, _13626_, _13619_);
  and (_13628_, _13627_, _13542_);
  nor (_13629_, _07769_, _07541_);
  or (_13630_, _13629_, _07700_);
  or (_13631_, _13630_, _13628_);
  nand (_13632_, _03742_, _07700_);
  and (_13633_, _13632_, _02966_);
  and (_13634_, _13633_, _13631_);
  nor (_13635_, _10662_, _07786_);
  nor (_13636_, _13635_, _13575_);
  nor (_13637_, _13636_, _02966_);
  or (_13638_, _13637_, _03861_);
  or (_13639_, _13638_, _13634_);
  and (_13640_, _13639_, _13535_);
  or (_13641_, _13640_, _03850_);
  and (_13642_, _06113_, _04654_);
  nor (_13643_, _13642_, _13528_);
  nand (_13644_, _13643_, _03850_);
  and (_13645_, _13644_, _02970_);
  and (_13646_, _13645_, _13641_);
  nor (_13647_, _10719_, _07325_);
  nor (_13648_, _13647_, _13528_);
  nor (_13649_, _13648_, _02970_);
  or (_13650_, _13649_, _06731_);
  or (_13651_, _13650_, _13646_);
  or (_13652_, _06992_, _06737_);
  and (_13653_, _13652_, _13651_);
  and (_13654_, _13653_, _02552_);
  nor (_13655_, _03742_, _02552_);
  or (_13656_, _13655_, _02974_);
  or (_13657_, _13656_, _13654_);
  and (_13658_, _04654_, _03660_);
  nor (_13659_, _13658_, _13562_);
  or (_13660_, _13659_, _05261_);
  and (_13661_, _13660_, _07808_);
  and (_13662_, _13661_, _13657_);
  or (_13663_, _13662_, _13532_);
  and (_13664_, _13663_, _07816_);
  and (_13665_, _07817_, _07217_);
  nor (_13666_, _08819_, _08817_);
  not (_13667_, _13666_);
  or (_13668_, _13667_, _13665_);
  or (_13669_, _13668_, _13664_);
  or (_13670_, _13666_, _07217_);
  and (_13671_, _13670_, _07833_);
  and (_13672_, _13671_, _13669_);
  and (_13673_, _07166_, _07832_);
  or (_13674_, _13673_, _03105_);
  or (_13675_, _13674_, _13672_);
  or (_13676_, _10610_, _03106_);
  and (_13677_, _13676_, _07846_);
  and (_13678_, _13677_, _13675_);
  and (_13679_, _07319_, _07762_);
  or (_13680_, _13679_, _02977_);
  or (_13681_, _13680_, _13678_);
  and (_13682_, _13681_, _13531_);
  or (_13683_, _13682_, _03107_);
  or (_13684_, _13528_, _07104_);
  and (_13685_, _13684_, _07868_);
  and (_13686_, _13685_, _13683_);
  or (_13687_, _13686_, _13527_);
  and (_13688_, _13687_, _07876_);
  and (_13689_, _07164_, _03499_);
  or (_13690_, _13689_, _03092_);
  or (_13691_, _13690_, _13688_);
  or (_13692_, _10608_, _03093_);
  and (_13693_, _13692_, _07886_);
  and (_13694_, _13693_, _13691_);
  and (_13695_, _07880_, _07761_);
  or (_13696_, _13695_, _13694_);
  and (_13697_, _13696_, _03881_);
  and (_13698_, _10613_, _04654_);
  nor (_13699_, _13698_, _13528_);
  nor (_13700_, _13699_, _03881_);
  or (_13701_, _13700_, _03242_);
  or (_13702_, _13701_, _13697_);
  and (_13703_, _13702_, _13526_);
  and (_13704_, _04120_, _02588_);
  or (_13705_, _13704_, _13703_);
  nand (_13706_, _13704_, _07216_);
  and (_13707_, _13706_, _03525_);
  and (_13708_, _13707_, _13705_);
  nor (_13709_, _07216_, _03525_);
  or (_13710_, _13709_, _07315_);
  or (_13711_, _13710_, _13708_);
  nand (_13712_, _07165_, _07315_);
  and (_13713_, _13712_, _03098_);
  and (_13714_, _13713_, _13711_);
  nand (_13715_, _10609_, _07902_);
  and (_13716_, _13715_, _07901_);
  or (_13717_, _13716_, _13714_);
  and (_13718_, _13717_, _13525_);
  or (_13719_, _13718_, _02994_);
  nor (_13720_, _10612_, _07325_);
  or (_13721_, _13720_, _13528_);
  or (_13722_, _13721_, _07120_);
  and (_13723_, _13722_, _07241_);
  and (_13724_, _13723_, _13719_);
  and (_13725_, _07298_, _07293_);
  nor (_13726_, _13725_, _07299_);
  and (_13727_, _13726_, _07912_);
  or (_13728_, _13727_, _07236_);
  or (_13729_, _13728_, _13724_);
  and (_13730_, _13729_, _13524_);
  or (_13731_, _13730_, _03103_);
  and (_13732_, _08008_, _08004_);
  nor (_13733_, _13732_, _08009_);
  or (_13734_, _13733_, _03104_);
  and (_13735_, _13734_, _08029_);
  and (_13736_, _13735_, _13731_);
  and (_13737_, _08039_, _08037_);
  nor (_13738_, _13737_, _08040_);
  and (_13739_, _13738_, _07946_);
  or (_13740_, _13739_, _08027_);
  or (_13741_, _13740_, _13736_);
  nand (_13742_, _08027_, _02658_);
  and (_13743_, _13742_, _07193_);
  and (_13744_, _13743_, _13741_);
  nor (_13745_, _07218_, _07217_);
  nor (_13746_, _13745_, _07219_);
  and (_13747_, _13746_, _13285_);
  or (_13748_, _13747_, _07183_);
  or (_13749_, _13748_, _13744_);
  nor (_13750_, _07167_, _07166_);
  nor (_13751_, _13750_, _07168_);
  or (_13752_, _13751_, _08792_);
  and (_13753_, _13752_, _13749_);
  or (_13754_, _13753_, _02856_);
  and (_13755_, _08082_, _07682_);
  nor (_13756_, _13755_, _08083_);
  or (_13757_, _13756_, _02857_);
  and (_13758_, _13757_, _08074_);
  and (_13759_, _13758_, _13754_);
  nor (_13760_, _08117_, _07762_);
  nor (_13761_, _13760_, _08118_);
  and (_13762_, _13761_, _08073_);
  or (_13763_, _13762_, _07143_);
  or (_13764_, _13763_, _13759_);
  and (_13765_, _13764_, _13521_);
  or (_13766_, _13765_, _03133_);
  or (_13767_, _13564_, _03138_);
  and (_13768_, _13767_, _08139_);
  and (_13769_, _13768_, _13766_);
  nor (_13770_, _08168_, _08144_);
  not (_13771_, _13770_);
  and (_13772_, _13771_, _08138_);
  or (_13773_, _13772_, _08143_);
  or (_13774_, _13773_, _13769_);
  nand (_13775_, _08143_, _06908_);
  and (_13776_, _13775_, _03142_);
  and (_13777_, _13776_, _13774_);
  nor (_13778_, _13596_, _03142_);
  or (_13779_, _13778_, _02852_);
  or (_13780_, _13779_, _13777_);
  nor (_13781_, _13563_, _13528_);
  nand (_13782_, _13781_, _02852_);
  and (_13783_, _13782_, _08161_);
  and (_13784_, _13783_, _13780_);
  and (_13785_, _13770_, _08160_);
  or (_13786_, _13785_, _08167_);
  or (_13787_, _13786_, _13784_);
  nand (_13788_, _08167_, _06908_);
  and (_13789_, _13788_, _34446_);
  and (_13790_, _13789_, _13787_);
  or (_13791_, _13790_, _13520_);
  and (_35614_[1], _13791_, _35583_);
  nor (_13792_, _34446_, _06908_);
  nand (_13793_, _07143_, _02477_);
  and (_13794_, _07220_, _07214_);
  nor (_13795_, _13794_, _07221_);
  or (_13796_, _13795_, _07183_);
  and (_13797_, _13796_, _09455_);
  and (_13798_, _07929_, _07373_);
  nor (_13799_, _13798_, _07930_);
  or (_13800_, _13799_, _07917_);
  nand (_13801_, _07899_, _08114_);
  nand (_13802_, _07212_, _03242_);
  or (_13803_, _07160_, _07876_);
  nor (_13804_, _04654_, _06908_);
  and (_13805_, _10936_, _04654_);
  nor (_13806_, _13805_, _13804_);
  nand (_13807_, _13806_, _02977_);
  nor (_13808_, _07325_, _04413_);
  nor (_13809_, _13808_, _13804_);
  nand (_13810_, _13809_, _03861_);
  nand (_13811_, _07476_, _04413_);
  nor (_13812_, _07625_, _07406_);
  or (_13813_, _06117_, _07408_);
  nor (_13814_, _07413_, _04413_);
  nor (_13815_, _07415_, \oc8051_golden_model_1.ACC [2]);
  and (_13816_, _07415_, \oc8051_golden_model_1.ACC [2]);
  nor (_13817_, _13816_, _13815_);
  nand (_13818_, _13817_, _07413_);
  nand (_13819_, _13818_, _07408_);
  or (_13820_, _13819_, _13814_);
  and (_13821_, _13820_, _07406_);
  and (_13822_, _13821_, _13813_);
  or (_13823_, _13822_, _13812_);
  and (_13824_, _13823_, _07429_);
  and (_13825_, _07434_, \oc8051_golden_model_1.XRAM_DATA_IN [2]);
  or (_13826_, _13825_, _03806_);
  or (_13827_, _13826_, _13824_);
  or (_13828_, _06117_, _05311_);
  and (_13829_, _13828_, _06162_);
  and (_13830_, _13829_, _13827_);
  nor (_13831_, _10824_, _07325_);
  nor (_13832_, _13831_, _13804_);
  nor (_13833_, _13832_, _06162_);
  or (_13834_, _13833_, _07402_);
  or (_13835_, _13834_, _13830_);
  and (_13836_, _13568_, \oc8051_golden_model_1.ACC [2]);
  and (_13837_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.ACC [1]);
  nor (_13838_, _13837_, _07440_);
  nor (_13839_, _13838_, _13568_);
  nor (_13840_, _13839_, _13836_);
  nand (_13841_, _13840_, _07402_);
  and (_13842_, _13841_, _02939_);
  and (_13843_, _13842_, _13835_);
  nor (_13844_, _05291_, _06908_);
  and (_13845_, _10815_, _05291_);
  nor (_13846_, _13845_, _13844_);
  nor (_13847_, _13846_, _03186_);
  nor (_13848_, _13809_, _03693_);
  or (_13849_, _13848_, _07476_);
  or (_13850_, _13849_, _13847_);
  or (_13851_, _13850_, _13843_);
  and (_13852_, _13851_, _13811_);
  or (_13853_, _13852_, _03374_);
  or (_13854_, _06117_, _03375_);
  and (_13855_, _13854_, _02943_);
  and (_13856_, _13855_, _13853_);
  nor (_13857_, _07625_, _02943_);
  or (_13858_, _13857_, _07486_);
  or (_13859_, _13858_, _13856_);
  nand (_13860_, _07486_, _06762_);
  and (_13861_, _13860_, _13859_);
  or (_13862_, _13861_, _02796_);
  and (_13863_, _10818_, _05291_);
  nor (_13864_, _13863_, _13844_);
  nand (_13865_, _13864_, _02796_);
  and (_13866_, _13865_, _06189_);
  and (_13867_, _13866_, _13862_);
  and (_13868_, _13845_, _10814_);
  nor (_13869_, _13868_, _13844_);
  nor (_13870_, _13869_, _06189_);
  or (_13871_, _13870_, _06195_);
  or (_13872_, _13871_, _13867_);
  nor (_13873_, _06659_, _06657_);
  nor (_13874_, _13873_, _06660_);
  or (_13875_, _13874_, _06201_);
  and (_13876_, _13875_, _13872_);
  or (_13877_, _13876_, _07401_);
  and (_13878_, _03989_, \oc8051_golden_model_1.ACC [1]);
  and (_13879_, _03805_, _02658_);
  nor (_13880_, _13879_, _07217_);
  nor (_13881_, _13880_, _13878_);
  nor (_13882_, _13881_, _07213_);
  and (_13883_, _13881_, _07213_);
  nor (_13884_, _13883_, _13882_);
  nor (_13885_, _13287_, _07217_);
  not (_13886_, _13885_);
  or (_13887_, _13886_, _13884_);
  and (_13888_, _13887_, \oc8051_golden_model_1.PSW [7]);
  nor (_13889_, _13884_, \oc8051_golden_model_1.PSW [7]);
  or (_13890_, _13889_, _13888_);
  nand (_13891_, _13886_, _13884_);
  and (_13892_, _13891_, _13890_);
  nor (_13893_, _13892_, _07329_);
  or (_13894_, _13893_, _09285_);
  and (_13895_, _13894_, _13877_);
  and (_13896_, _05844_, \oc8051_golden_model_1.ACC [1]);
  and (_13897_, _06114_, _02658_);
  nor (_13898_, _13897_, _07166_);
  nor (_13899_, _13898_, _13896_);
  nor (_13900_, _13899_, _07162_);
  and (_13901_, _13899_, _07162_);
  nor (_13902_, _13901_, _13900_);
  nor (_13903_, _13423_, _07166_);
  not (_13904_, _13903_);
  or (_13905_, _13904_, _13902_);
  and (_13906_, _13905_, \oc8051_golden_model_1.PSW [7]);
  nor (_13907_, _13902_, \oc8051_golden_model_1.PSW [7]);
  or (_13908_, _13907_, _13906_);
  nand (_13909_, _13904_, _13902_);
  and (_13910_, _13909_, _13908_);
  nor (_13911_, _13910_, _07330_);
  or (_13912_, _13911_, _02898_);
  or (_13913_, _13912_, _13895_);
  nor (_13914_, _07656_, _07654_);
  nor (_13915_, _13914_, _07657_);
  and (_13916_, _07685_, \oc8051_golden_model_1.PSW [7]);
  not (_13917_, _13916_);
  nor (_13918_, _13917_, _13915_);
  and (_13919_, _13917_, _13915_);
  nor (_13920_, _13919_, _13918_);
  nand (_13921_, _13920_, _02898_);
  and (_13922_, _13921_, _07541_);
  and (_13923_, _13922_, _13913_);
  nor (_13924_, _02835_, \oc8051_golden_model_1.ACC [0]);
  nor (_13925_, _13924_, _07762_);
  nor (_13926_, _13925_, _09959_);
  nor (_13927_, _08115_, _13926_);
  and (_13928_, _08115_, _13926_);
  nor (_13929_, _13928_, _13927_);
  not (_13930_, _08831_);
  or (_13931_, _13930_, _13929_);
  and (_13932_, _13931_, \oc8051_golden_model_1.PSW [7]);
  nor (_13933_, _13929_, \oc8051_golden_model_1.PSW [7]);
  or (_13934_, _13933_, _13932_);
  nand (_13935_, _13930_, _13929_);
  and (_13936_, _13935_, _13934_);
  nor (_13937_, _13936_, _07541_);
  or (_13938_, _13937_, _07700_);
  or (_13939_, _13938_, _13923_);
  nand (_13940_, _03320_, _07700_);
  and (_13941_, _13940_, _02966_);
  and (_13942_, _13941_, _13939_);
  nor (_13943_, _10866_, _07786_);
  nor (_13944_, _13943_, _13844_);
  nor (_13945_, _13944_, _02966_);
  or (_13946_, _13945_, _03861_);
  or (_13947_, _13946_, _13942_);
  and (_13948_, _13947_, _13810_);
  or (_13949_, _13948_, _03850_);
  and (_13950_, _06117_, _04654_);
  nor (_13951_, _13950_, _13804_);
  nand (_13952_, _13951_, _03850_);
  and (_13953_, _13952_, _02970_);
  and (_13954_, _13953_, _13949_);
  nor (_13955_, _10922_, _07325_);
  nor (_13956_, _13955_, _13804_);
  nor (_13957_, _13956_, _02970_);
  or (_13958_, _13957_, _06731_);
  or (_13959_, _13958_, _13954_);
  or (_13960_, _06928_, _06737_);
  and (_13961_, _13960_, _13959_);
  and (_13962_, _13961_, _02552_);
  nor (_13963_, _03320_, _02552_);
  or (_13964_, _13963_, _02974_);
  or (_13965_, _13964_, _13962_);
  and (_13966_, _04654_, _05690_);
  nor (_13967_, _13966_, _13804_);
  nand (_13968_, _13967_, _02974_);
  and (_13969_, _13968_, _07808_);
  and (_13970_, _13969_, _13965_);
  nor (_13971_, _07808_, _03320_);
  or (_13972_, _13971_, _07817_);
  or (_13973_, _13972_, _13970_);
  nor (_13974_, _07827_, _03483_);
  nor (_13975_, _08817_, _07214_);
  or (_13976_, _13975_, _08818_);
  and (_13977_, _13976_, _13974_);
  and (_13978_, _13977_, _13973_);
  or (_13979_, _07827_, _07823_);
  and (_13980_, _13979_, _07213_);
  or (_13981_, _13980_, _03484_);
  or (_13982_, _13981_, _13978_);
  nand (_13983_, _07214_, _03484_);
  and (_13984_, _13983_, _07833_);
  and (_13985_, _13984_, _13982_);
  and (_13986_, _07162_, _07832_);
  or (_13987_, _13986_, _03105_);
  or (_13988_, _13987_, _13985_);
  or (_13989_, _10942_, _03106_);
  and (_13990_, _13989_, _07846_);
  and (_13991_, _13990_, _13988_);
  and (_13992_, _07319_, _08115_);
  or (_13993_, _13992_, _02977_);
  or (_13994_, _13993_, _13991_);
  and (_13995_, _13994_, _13807_);
  or (_13996_, _13995_, _03107_);
  or (_13997_, _13804_, _07104_);
  and (_13998_, _13997_, _07868_);
  and (_13999_, _13998_, _13996_);
  and (_14000_, _07869_, _07211_);
  or (_14001_, _14000_, _03499_);
  or (_14002_, _14001_, _13999_);
  and (_14003_, _14002_, _13803_);
  or (_14004_, _14003_, _03092_);
  or (_14005_, _10940_, _03093_);
  and (_14006_, _14005_, _07886_);
  and (_14007_, _14006_, _14004_);
  and (_14008_, _07880_, _08113_);
  or (_14009_, _14008_, _14007_);
  and (_14010_, _14009_, _03881_);
  or (_14011_, _13967_, _10941_);
  nor (_14012_, _14011_, _03881_);
  or (_14013_, _14012_, _03242_);
  or (_14014_, _14013_, _14010_);
  and (_14015_, _14014_, _13802_);
  or (_14016_, _14015_, _13704_);
  nand (_14017_, _13704_, _07212_);
  and (_14018_, _14017_, _03525_);
  and (_14019_, _14018_, _14016_);
  nor (_14020_, _07212_, _03525_);
  or (_14021_, _14020_, _07315_);
  or (_14022_, _14021_, _14019_);
  nand (_14023_, _07161_, _07315_);
  and (_14024_, _14023_, _03098_);
  and (_14025_, _14024_, _14022_);
  nand (_14026_, _10941_, _07902_);
  and (_14027_, _14026_, _07901_);
  or (_14028_, _14027_, _14025_);
  and (_14029_, _14028_, _13801_);
  or (_14030_, _14029_, _02994_);
  nor (_14031_, _10935_, _07325_);
  nor (_14032_, _14031_, _13804_);
  nand (_14033_, _14032_, _02994_);
  and (_14034_, _14033_, _07241_);
  and (_14035_, _14034_, _14030_);
  and (_14036_, _07300_, _07286_);
  nor (_14037_, _14036_, _07301_);
  and (_14038_, _14037_, _07912_);
  or (_14039_, _14038_, _07236_);
  or (_14040_, _14039_, _14035_);
  and (_14041_, _14040_, _13800_);
  or (_14042_, _14041_, _03103_);
  and (_14043_, _08010_, _07998_);
  nor (_14044_, _14043_, _08011_);
  or (_14045_, _14044_, _03104_);
  and (_14046_, _14045_, _08029_);
  and (_14047_, _14046_, _14042_);
  and (_14048_, _08041_, _07740_);
  nor (_14049_, _14048_, _08042_);
  and (_14050_, _14049_, _07946_);
  or (_14051_, _14050_, _08027_);
  or (_14052_, _14051_, _14047_);
  nand (_14053_, _08027_, _02477_);
  and (_14054_, _14053_, _07193_);
  and (_14055_, _14054_, _14052_);
  or (_14056_, _14055_, _13797_);
  and (_14057_, _07169_, _07163_);
  nor (_14058_, _14057_, _07170_);
  or (_14059_, _14058_, _08792_);
  and (_14060_, _14059_, _14056_);
  or (_14061_, _14060_, _02856_);
  and (_14062_, _08084_, _07656_);
  nor (_14063_, _14062_, _08085_);
  or (_14064_, _14063_, _02857_);
  and (_14065_, _14064_, _08074_);
  and (_14066_, _14065_, _14061_);
  and (_14067_, _08119_, _08116_);
  nor (_14068_, _14067_, _08120_);
  and (_14069_, _14068_, _08073_);
  or (_14070_, _14069_, _07143_);
  or (_14071_, _14070_, _14066_);
  and (_14072_, _14071_, _13793_);
  or (_14073_, _14072_, _03133_);
  nand (_14074_, _13832_, _03133_);
  and (_14075_, _14074_, _08139_);
  and (_14076_, _14075_, _14073_);
  and (_14077_, _07440_, _02658_);
  nor (_14078_, _08144_, _06908_);
  or (_14079_, _14078_, _14077_);
  and (_14080_, _14079_, _08138_);
  or (_14081_, _14080_, _08143_);
  or (_14082_, _14081_, _14076_);
  nand (_14083_, _08143_, _02605_);
  and (_14084_, _14083_, _03142_);
  and (_14085_, _14084_, _14082_);
  nor (_14086_, _13864_, _03142_);
  or (_14087_, _14086_, _02852_);
  or (_14088_, _14087_, _14085_);
  and (_14089_, _10988_, _04654_);
  nor (_14090_, _14089_, _13804_);
  nand (_14091_, _14090_, _02852_);
  and (_14092_, _14091_, _08161_);
  and (_14093_, _14092_, _14088_);
  and (_14094_, _08168_, \oc8051_golden_model_1.ACC [2]);
  nor (_14095_, _08168_, \oc8051_golden_model_1.ACC [2]);
  nor (_14096_, _14095_, _14094_);
  nor (_14097_, _14096_, _08167_);
  nor (_14098_, _14097_, _09696_);
  or (_14099_, _14098_, _14093_);
  nand (_14100_, _08167_, _02605_);
  and (_14101_, _14100_, _34446_);
  and (_14102_, _14101_, _14099_);
  or (_14103_, _14102_, _13792_);
  and (_35614_[2], _14103_, _35583_);
  nor (_14104_, _34446_, _02605_);
  nor (_14105_, _07210_, _07208_);
  nor (_14106_, _14105_, _07222_);
  and (_14107_, _14105_, _07222_);
  nor (_14108_, _14107_, _14106_);
  nand (_14109_, _14108_, _13285_);
  and (_14110_, _07302_, _07280_);
  nor (_14111_, _14110_, _07303_);
  or (_14112_, _14111_, _07241_);
  nor (_14113_, _04654_, _02605_);
  and (_14114_, _11128_, _04654_);
  nor (_14115_, _14114_, _14113_);
  nand (_14116_, _14115_, _02977_);
  not (_14117_, _03488_);
  and (_14118_, _07816_, _14117_);
  and (_14119_, _07807_, _02774_);
  nor (_14120_, _07325_, _04226_);
  nor (_14121_, _14120_, _14113_);
  nand (_14122_, _14121_, _03861_);
  nor (_14123_, _05291_, _02605_);
  and (_14124_, _11011_, _05291_);
  and (_14125_, _14124_, _11040_);
  nor (_14126_, _14125_, _14123_);
  nor (_14127_, _14126_, _06189_);
  nand (_14128_, _07476_, _04226_);
  nor (_14129_, _07611_, _07406_);
  or (_14130_, _06116_, _07408_);
  nor (_14131_, _07413_, _04226_);
  nor (_14132_, _07415_, \oc8051_golden_model_1.ACC [3]);
  and (_14133_, _07415_, \oc8051_golden_model_1.ACC [3]);
  nor (_14134_, _14133_, _14132_);
  nand (_14135_, _14134_, _07413_);
  nand (_14136_, _14135_, _07408_);
  or (_14137_, _14136_, _14131_);
  and (_14138_, _14137_, _07406_);
  and (_14139_, _14138_, _14130_);
  or (_14140_, _14139_, _14129_);
  and (_14141_, _14140_, _07429_);
  and (_14142_, _07434_, \oc8051_golden_model_1.XRAM_DATA_IN [3]);
  or (_14143_, _14142_, _03806_);
  or (_14144_, _14143_, _14141_);
  or (_14145_, _06116_, _05311_);
  and (_14146_, _14145_, _06162_);
  and (_14147_, _14146_, _14144_);
  nor (_14148_, _11014_, _07325_);
  nor (_14149_, _14148_, _14113_);
  nor (_14150_, _14149_, _06162_);
  or (_14151_, _14150_, _07402_);
  or (_14152_, _14151_, _14147_);
  not (_14153_, \oc8051_golden_model_1.PSW [6]);
  nor (_14154_, _07440_, _14153_);
  nor (_14155_, _14154_, \oc8051_golden_model_1.ACC [3]);
  nor (_14156_, _14155_, _07441_);
  or (_14157_, _14156_, _09879_);
  and (_14158_, _14157_, _02939_);
  and (_14159_, _14158_, _14152_);
  nor (_14160_, _14124_, _14123_);
  nor (_14161_, _14160_, _03186_);
  nor (_14162_, _14121_, _03693_);
  or (_14163_, _14162_, _07476_);
  or (_14164_, _14163_, _14161_);
  or (_14165_, _14164_, _14159_);
  and (_14166_, _14165_, _14128_);
  or (_14167_, _14166_, _03374_);
  or (_14168_, _06116_, _03375_);
  and (_14169_, _14168_, _02943_);
  and (_14170_, _14169_, _14167_);
  nor (_14171_, _07611_, _02943_);
  or (_14172_, _14171_, _07486_);
  or (_14173_, _14172_, _14170_);
  nand (_14174_, _07486_, _05719_);
  and (_14175_, _14174_, _14173_);
  or (_14176_, _14175_, _02796_);
  and (_14177_, _11009_, _05291_);
  nor (_14178_, _14177_, _14123_);
  nand (_14179_, _14178_, _02796_);
  and (_14180_, _14179_, _06189_);
  and (_14181_, _14180_, _14176_);
  or (_14182_, _14181_, _14127_);
  and (_14183_, _14182_, _06201_);
  nor (_14184_, _06662_, _06660_);
  nor (_14185_, _14184_, _06663_);
  nand (_14186_, _14185_, _06195_);
  nand (_14187_, _14186_, _07400_);
  or (_14188_, _14187_, _14183_);
  and (_14189_, _04413_, \oc8051_golden_model_1.ACC [2]);
  nor (_14190_, _13882_, _14189_);
  nor (_14191_, _14190_, _14105_);
  and (_14192_, _14190_, _14105_);
  nor (_14193_, _14192_, _14191_);
  and (_14194_, _14193_, \oc8051_golden_model_1.PSW [7]);
  nor (_14195_, _14193_, \oc8051_golden_model_1.PSW [7]);
  nor (_14196_, _14195_, _14194_);
  and (_14197_, _14196_, _13888_);
  nor (_14198_, _14196_, _13888_);
  or (_14199_, _14198_, _14197_);
  nand (_14200_, _14199_, _07401_);
  and (_14201_, _14200_, _14188_);
  or (_14202_, _14201_, _07329_);
  nor (_14203_, _07159_, _07158_);
  and (_14204_, _05980_, \oc8051_golden_model_1.ACC [2]);
  nor (_14205_, _13900_, _14204_);
  nor (_14206_, _14205_, _14203_);
  and (_14207_, _14205_, _14203_);
  nor (_14208_, _14207_, _14206_);
  and (_14209_, _14208_, \oc8051_golden_model_1.PSW [7]);
  nor (_14210_, _14208_, \oc8051_golden_model_1.PSW [7]);
  nor (_14211_, _14210_, _14209_);
  and (_14212_, _14211_, _13906_);
  nor (_14213_, _14211_, _13906_);
  or (_14214_, _14213_, _14212_);
  nand (_14215_, _14214_, _07329_);
  and (_14216_, _14215_, _02899_);
  and (_14217_, _14216_, _14202_);
  nor (_14218_, _07680_, _07658_);
  and (_14219_, _07680_, _07658_);
  or (_14220_, _14219_, _14218_);
  not (_14221_, _13918_);
  and (_14222_, _14221_, _14220_);
  nor (_14223_, _14222_, _07687_);
  nor (_14224_, _14223_, _02899_);
  or (_14225_, _14224_, _07540_);
  or (_14226_, _14225_, _14217_);
  and (_14227_, _03320_, \oc8051_golden_model_1.ACC [2]);
  nor (_14228_, _13927_, _14227_);
  nor (_14229_, _08832_, _14228_);
  and (_14230_, _08832_, _14228_);
  nor (_14231_, _14230_, _14229_);
  and (_14232_, _14231_, \oc8051_golden_model_1.PSW [7]);
  nor (_14233_, _14231_, \oc8051_golden_model_1.PSW [7]);
  nor (_14234_, _14233_, _14232_);
  and (_14235_, _14234_, _13932_);
  nor (_14236_, _14234_, _13932_);
  nor (_14237_, _14236_, _14235_);
  or (_14238_, _14237_, _07541_);
  and (_14239_, _14238_, _14226_);
  or (_14240_, _14239_, _07700_);
  or (_14241_, _02774_, _02499_);
  and (_14242_, _14241_, _02966_);
  and (_14243_, _14242_, _14240_);
  nor (_14244_, _11058_, _07786_);
  nor (_14245_, _14244_, _14123_);
  nor (_14246_, _14245_, _02966_);
  or (_14247_, _14246_, _03861_);
  or (_14248_, _14247_, _14243_);
  and (_14249_, _14248_, _14122_);
  or (_14250_, _14249_, _03850_);
  and (_14251_, _06116_, _04654_);
  nor (_14252_, _14251_, _14113_);
  nand (_14253_, _14252_, _03850_);
  and (_14254_, _14253_, _02970_);
  and (_14255_, _14254_, _14250_);
  nor (_14256_, _11114_, _07325_);
  nor (_14257_, _14256_, _14113_);
  nor (_14258_, _14257_, _02970_);
  or (_14259_, _14258_, _06731_);
  or (_14260_, _14259_, _14255_);
  or (_14261_, _06873_, _06737_);
  and (_14262_, _14261_, _14260_);
  and (_14263_, _14262_, _02552_);
  and (_14264_, _02774_, _02476_);
  or (_14265_, _14264_, _02974_);
  or (_14266_, _14265_, _14263_);
  and (_14267_, _04654_, _05616_);
  nor (_14268_, _14267_, _14113_);
  nand (_14269_, _14268_, _02974_);
  and (_14270_, _14269_, _07808_);
  and (_14271_, _14270_, _14266_);
  or (_14272_, _14271_, _14119_);
  and (_14273_, _14272_, _14118_);
  not (_14274_, _07821_);
  and (_14275_, _07828_, _14274_);
  not (_14276_, _14118_);
  nand (_14277_, _14276_, _14105_);
  nand (_14278_, _14277_, _14275_);
  or (_14279_, _14278_, _14273_);
  or (_14280_, _14275_, _14105_);
  and (_14281_, _14280_, _07833_);
  and (_14282_, _14281_, _14279_);
  and (_14283_, _14203_, _07832_);
  or (_14284_, _14283_, _03105_);
  or (_14285_, _14284_, _14282_);
  or (_14286_, _11134_, _03106_);
  and (_14287_, _14286_, _07846_);
  and (_14288_, _14287_, _14285_);
  and (_14289_, _07319_, _08832_);
  or (_14290_, _14289_, _02977_);
  or (_14291_, _14290_, _14288_);
  and (_14292_, _14291_, _14116_);
  or (_14293_, _14292_, _03107_);
  or (_14294_, _14113_, _07104_);
  and (_14295_, _14294_, _07868_);
  and (_14296_, _14295_, _14293_);
  and (_14297_, _07869_, _07208_);
  or (_14298_, _14297_, _03499_);
  or (_14299_, _14298_, _14296_);
  or (_14300_, _07158_, _07876_);
  and (_14301_, _14300_, _03093_);
  and (_14302_, _14301_, _14299_);
  or (_14303_, _11132_, _07880_);
  and (_14304_, _14303_, _07882_);
  or (_14305_, _14304_, _14302_);
  or (_14306_, _07886_, _08111_);
  and (_14307_, _14306_, _03881_);
  and (_14308_, _14307_, _14305_);
  not (_14309_, _02588_);
  nor (_14310_, _07238_, _14309_);
  or (_14311_, _14268_, _11133_);
  nor (_14312_, _14311_, _03881_);
  or (_14313_, _14312_, _14310_);
  or (_14314_, _14313_, _14308_);
  and (_14315_, _03857_, _02588_);
  and (_14316_, _14310_, _07210_);
  nor (_14317_, _14316_, _14315_);
  and (_14318_, _14317_, _14314_);
  not (_14319_, _07210_);
  and (_14320_, _14315_, _14319_);
  or (_14321_, _14320_, _07315_);
  or (_14322_, _14321_, _14318_);
  nand (_14323_, _07159_, _07315_);
  and (_14324_, _14323_, _03098_);
  and (_14325_, _14324_, _14322_);
  nand (_14326_, _11133_, _07902_);
  and (_14327_, _14326_, _07901_);
  or (_14328_, _14327_, _14325_);
  nand (_14329_, _07899_, _08112_);
  and (_14330_, _14329_, _07120_);
  and (_14331_, _14330_, _14328_);
  nor (_14332_, _11127_, _07325_);
  nor (_14333_, _14332_, _14113_);
  nor (_14334_, _14333_, _07120_);
  or (_14335_, _14334_, _07912_);
  or (_14336_, _14335_, _14331_);
  and (_14337_, _14336_, _14112_);
  or (_14338_, _14337_, _07236_);
  and (_14339_, _07931_, _07368_);
  nor (_14340_, _14339_, _07932_);
  or (_14341_, _14340_, _07917_);
  and (_14342_, _14341_, _03104_);
  and (_14343_, _14342_, _14338_);
  and (_14344_, _08012_, _07992_);
  nor (_14345_, _14344_, _08013_);
  and (_14346_, _14345_, _03103_);
  or (_14347_, _14346_, _07946_);
  or (_14348_, _14347_, _14343_);
  and (_14349_, _08043_, _07735_);
  nor (_14350_, _14349_, _08044_);
  or (_14351_, _14350_, _08029_);
  and (_14352_, _14351_, _08028_);
  and (_14353_, _14352_, _14348_);
  nand (_14354_, _08027_, \oc8051_golden_model_1.ACC [2]);
  nand (_14355_, _14354_, _07193_);
  or (_14356_, _14355_, _14353_);
  and (_14357_, _14356_, _14109_);
  or (_14358_, _14357_, _07183_);
  nor (_14359_, _14203_, _07171_);
  and (_14360_, _14203_, _07171_);
  nor (_14361_, _14360_, _14359_);
  nand (_14362_, _14361_, _07183_);
  and (_14363_, _14362_, _03125_);
  and (_14364_, _14363_, _14358_);
  nor (_14365_, _08086_, _07680_);
  and (_14366_, _08086_, _07680_);
  nor (_14367_, _14366_, _14365_);
  or (_14368_, _14367_, _02441_);
  and (_14369_, _14368_, _08772_);
  or (_14370_, _14369_, _14364_);
  nor (_14371_, _08121_, _08832_);
  and (_14372_, _08121_, _08832_);
  nor (_14373_, _14372_, _14371_);
  nand (_14374_, _14373_, _08073_);
  and (_14375_, _14374_, _09650_);
  and (_14376_, _14375_, _14370_);
  and (_14377_, _07143_, \oc8051_golden_model_1.ACC [2]);
  or (_14378_, _14377_, _03133_);
  or (_14379_, _14378_, _14376_);
  nand (_14380_, _14149_, _03133_);
  and (_14381_, _14380_, _08139_);
  and (_14382_, _14381_, _14379_);
  nor (_14383_, _14077_, _02605_);
  or (_14384_, _14383_, _08145_);
  and (_14385_, _14384_, _08138_);
  or (_14386_, _14385_, _08143_);
  or (_14387_, _14386_, _14382_);
  nand (_14388_, _08143_, _06814_);
  and (_14389_, _14388_, _03142_);
  and (_14390_, _14389_, _14387_);
  nor (_14391_, _14178_, _03142_);
  or (_14392_, _14391_, _02852_);
  or (_14393_, _14392_, _14390_);
  and (_14394_, _11185_, _04654_);
  nor (_14395_, _14394_, _14113_);
  nand (_14396_, _14395_, _02852_);
  and (_14397_, _14396_, _08161_);
  and (_14398_, _14397_, _14393_);
  or (_14399_, _14094_, \oc8051_golden_model_1.ACC [3]);
  and (_14400_, _14399_, _08169_);
  and (_14401_, _14400_, _08160_);
  or (_14402_, _14401_, _08167_);
  or (_14403_, _14402_, _14398_);
  nand (_14404_, _08167_, _06814_);
  and (_14405_, _14404_, _34446_);
  and (_14406_, _14405_, _14403_);
  or (_14407_, _14406_, _14104_);
  and (_35614_[3], _14407_, _35583_);
  nor (_14408_, _34446_, _06814_);
  nand (_14409_, _07899_, _08109_);
  and (_14410_, _03009_, _02588_);
  nand (_14411_, _14310_, _07205_);
  or (_14412_, _07155_, _07876_);
  nor (_14413_, _04654_, _06814_);
  and (_14414_, _11327_, _04654_);
  nor (_14415_, _14414_, _14413_);
  nand (_14416_, _14415_, _02977_);
  nor (_14417_, _05143_, _07325_);
  nor (_14418_, _14417_, _14413_);
  nand (_14419_, _14418_, _03861_);
  and (_14420_, _07688_, _07679_);
  nor (_14421_, _14420_, _07689_);
  nand (_14422_, _14421_, _02898_);
  and (_14423_, _14422_, _07541_);
  nand (_14424_, _07476_, _05143_);
  nor (_14425_, _11207_, _07325_);
  nor (_14426_, _14425_, _14413_);
  nand (_14427_, _14426_, _02932_);
  nor (_14428_, _07593_, _07406_);
  or (_14429_, _06121_, _07408_);
  nor (_14430_, _07413_, _05143_);
  or (_14431_, _07415_, \oc8051_golden_model_1.ACC [4]);
  nand (_14432_, _07415_, \oc8051_golden_model_1.ACC [4]);
  and (_14433_, _14432_, _14431_);
  and (_14434_, _14433_, _07413_);
  or (_14435_, _14434_, _03343_);
  or (_14436_, _14435_, _14430_);
  and (_14437_, _14436_, _07406_);
  and (_14438_, _14437_, _14429_);
  or (_14439_, _14438_, _14428_);
  and (_14440_, _14439_, _07429_);
  and (_14441_, _07434_, \oc8051_golden_model_1.XRAM_DATA_IN [4]);
  or (_14442_, _14441_, _02932_);
  or (_14443_, _14442_, _14440_);
  and (_14444_, _14443_, _14427_);
  or (_14445_, _14444_, _07402_);
  nor (_14446_, _07441_, \oc8051_golden_model_1.ACC [4]);
  nor (_14447_, _14446_, _07447_);
  not (_14448_, _14447_);
  nand (_14449_, _14448_, _07402_);
  and (_14450_, _14449_, _02939_);
  and (_14451_, _14450_, _14445_);
  nor (_14452_, _05291_, _06814_);
  and (_14453_, _11224_, _05291_);
  nor (_14454_, _14453_, _14452_);
  nor (_14455_, _14454_, _03186_);
  nor (_14456_, _14418_, _03693_);
  or (_14457_, _14456_, _07476_);
  or (_14458_, _14457_, _14455_);
  or (_14459_, _14458_, _14451_);
  and (_14460_, _14459_, _14424_);
  or (_14461_, _14460_, _03374_);
  or (_14462_, _06121_, _03375_);
  and (_14463_, _14462_, _02943_);
  and (_14464_, _14463_, _14461_);
  nor (_14465_, _07593_, _02943_);
  or (_14466_, _14465_, _07486_);
  or (_14467_, _14466_, _14464_);
  nand (_14468_, _07486_, _02658_);
  and (_14469_, _14468_, _14467_);
  or (_14470_, _14469_, _02796_);
  and (_14471_, _11203_, _05291_);
  nor (_14472_, _14471_, _14452_);
  nand (_14473_, _14472_, _02796_);
  and (_14474_, _14473_, _06189_);
  and (_14475_, _14474_, _14470_);
  and (_14476_, _14453_, _11239_);
  nor (_14477_, _14476_, _14452_);
  nor (_14478_, _14477_, _06189_);
  or (_14479_, _14478_, _06195_);
  or (_14480_, _14479_, _14475_);
  nor (_14481_, _06665_, _06663_);
  nor (_14482_, _14481_, _06666_);
  or (_14483_, _14482_, _06201_);
  and (_14484_, _14483_, _14480_);
  or (_14485_, _14484_, _07401_);
  or (_14486_, _14197_, _14194_);
  nor (_14487_, _04226_, \oc8051_golden_model_1.ACC [3]);
  nand (_14488_, _04226_, \oc8051_golden_model_1.ACC [3]);
  and (_14489_, _14190_, _14488_);
  or (_14490_, _14489_, _14487_);
  nor (_14491_, _14490_, _07206_);
  and (_14492_, _14490_, _07206_);
  nor (_14493_, _14492_, _14491_);
  and (_14494_, _14493_, \oc8051_golden_model_1.PSW [7]);
  nor (_14495_, _14493_, \oc8051_golden_model_1.PSW [7]);
  nor (_14496_, _14495_, _14494_);
  and (_14497_, _14496_, _14486_);
  nor (_14498_, _14496_, _14486_);
  nor (_14499_, _14498_, _14497_);
  or (_14500_, _14499_, _07400_);
  and (_14501_, _14500_, _14485_);
  or (_14502_, _14501_, _07329_);
  or (_14503_, _14212_, _14209_);
  and (_14504_, _06116_, _02605_);
  or (_14505_, _06116_, _02605_);
  and (_14506_, _14205_, _14505_);
  or (_14507_, _14506_, _14504_);
  nor (_14508_, _14507_, _07157_);
  and (_14509_, _14507_, _07157_);
  nor (_14510_, _14509_, _14508_);
  and (_14511_, _14510_, \oc8051_golden_model_1.PSW [7]);
  nor (_14512_, _14510_, \oc8051_golden_model_1.PSW [7]);
  nor (_14513_, _14512_, _14511_);
  and (_14514_, _14513_, _14503_);
  nor (_14515_, _14513_, _14503_);
  nor (_14516_, _14515_, _14514_);
  or (_14517_, _14516_, _07330_);
  and (_14518_, _14517_, _14502_);
  or (_14519_, _14518_, _02898_);
  and (_14520_, _14519_, _14423_);
  or (_14521_, _14235_, _14232_);
  or (_14522_, _14228_, _09965_);
  and (_14523_, _14522_, _09964_);
  nor (_14524_, _08110_, _14523_);
  and (_14525_, _08110_, _14523_);
  nor (_14526_, _14525_, _14524_);
  and (_14527_, _14526_, \oc8051_golden_model_1.PSW [7]);
  nor (_14528_, _14526_, \oc8051_golden_model_1.PSW [7]);
  nor (_14529_, _14528_, _14527_);
  and (_14530_, _14529_, _14521_);
  nor (_14531_, _14529_, _14521_);
  nor (_14532_, _14531_, _14530_);
  and (_14533_, _14532_, _07540_);
  or (_14534_, _14533_, _07700_);
  or (_14535_, _14534_, _14520_);
  nand (_14536_, _03620_, _07700_);
  and (_14537_, _14536_, _02966_);
  and (_14538_, _14537_, _14535_);
  nor (_14539_, _11257_, _07786_);
  nor (_14540_, _14539_, _14452_);
  nor (_14541_, _14540_, _02966_);
  or (_14542_, _14541_, _03861_);
  or (_14543_, _14542_, _14538_);
  and (_14544_, _14543_, _14419_);
  or (_14545_, _14544_, _03850_);
  and (_14546_, _06121_, _04654_);
  nor (_14547_, _14546_, _14413_);
  nand (_14548_, _14547_, _03850_);
  and (_14549_, _14548_, _02970_);
  and (_14550_, _14549_, _14545_);
  nor (_14551_, _11313_, _07325_);
  nor (_14552_, _14551_, _14413_);
  nor (_14553_, _14552_, _02970_);
  or (_14554_, _14553_, _06731_);
  or (_14555_, _14554_, _14550_);
  or (_14556_, _06823_, _06737_);
  and (_14557_, _14556_, _14555_);
  and (_14558_, _14557_, _02552_);
  nor (_14559_, _03620_, _02552_);
  or (_14560_, _14559_, _02974_);
  or (_14561_, _14560_, _14558_);
  and (_14562_, _05629_, _04654_);
  nor (_14563_, _14562_, _14413_);
  nand (_14564_, _14563_, _02974_);
  and (_14565_, _14564_, _07808_);
  and (_14566_, _14565_, _14561_);
  nor (_14567_, _07808_, _03620_);
  or (_14568_, _14567_, _07817_);
  or (_14569_, _14568_, _14566_);
  or (_14570_, _07816_, _07206_);
  and (_14571_, _14570_, _13666_);
  and (_14572_, _14571_, _14569_);
  and (_14573_, _13667_, _07206_);
  or (_14574_, _14573_, _07832_);
  or (_14575_, _14574_, _14572_);
  or (_14576_, _07157_, _03487_);
  nand (_14577_, _07832_, _02519_);
  or (_14578_, _14577_, _07157_);
  and (_14579_, _14578_, _14576_);
  and (_14580_, _14579_, _14575_);
  or (_14581_, _14580_, _03105_);
  or (_14582_, _11333_, _03106_);
  and (_14583_, _14582_, _07846_);
  and (_14584_, _14583_, _14581_);
  and (_14585_, _07319_, _08110_);
  or (_14586_, _14585_, _02977_);
  or (_14587_, _14586_, _14584_);
  and (_14588_, _14587_, _14416_);
  or (_14589_, _14588_, _03107_);
  or (_14590_, _14413_, _07104_);
  and (_14591_, _14590_, _07868_);
  and (_14592_, _14591_, _14589_);
  and (_14593_, _07869_, _07204_);
  or (_14594_, _14593_, _03499_);
  or (_14595_, _14594_, _14592_);
  and (_14596_, _14595_, _14412_);
  or (_14597_, _14596_, _03092_);
  or (_14598_, _11331_, _03093_);
  and (_14599_, _14598_, _07886_);
  and (_14600_, _14599_, _14597_);
  and (_14601_, _07880_, _08108_);
  or (_14602_, _14601_, _14600_);
  and (_14603_, _14602_, _03881_);
  or (_14604_, _14563_, _11332_);
  nor (_14605_, _14604_, _03881_);
  or (_14606_, _14605_, _14310_);
  or (_14607_, _14606_, _14603_);
  and (_14608_, _14607_, _14411_);
  or (_14609_, _14608_, _14410_);
  nand (_14610_, _14410_, _07205_);
  and (_14611_, _14610_, _03525_);
  and (_14612_, _14611_, _14609_);
  nor (_14613_, _07205_, _03525_);
  or (_14614_, _14613_, _07315_);
  or (_14615_, _14614_, _14612_);
  nand (_14616_, _07156_, _07315_);
  and (_14617_, _14616_, _03098_);
  and (_14618_, _14617_, _14615_);
  nand (_14619_, _11332_, _07902_);
  and (_14620_, _14619_, _07901_);
  or (_14621_, _14620_, _14618_);
  and (_14622_, _14621_, _14409_);
  or (_14623_, _14622_, _02994_);
  nor (_14624_, _11326_, _07325_);
  nor (_14625_, _14624_, _14413_);
  nand (_14626_, _14625_, _02994_);
  and (_14627_, _14626_, _07241_);
  and (_14628_, _14627_, _14623_);
  and (_14629_, _07304_, _07271_);
  nor (_14630_, _14629_, _07305_);
  and (_14631_, _14630_, _07912_);
  or (_14632_, _14631_, _07236_);
  or (_14633_, _14632_, _14628_);
  and (_14634_, _07933_, _07360_);
  nor (_14635_, _14634_, _07934_);
  or (_14636_, _14635_, _07917_);
  and (_14637_, _14636_, _03104_);
  and (_14638_, _14637_, _14633_);
  and (_14639_, _08014_, _07986_);
  nor (_14640_, _14639_, _08015_);
  or (_14641_, _14640_, _07946_);
  and (_14642_, _14641_, _07948_);
  or (_14643_, _14642_, _14638_);
  and (_14644_, _08045_, _07728_);
  nor (_14645_, _14644_, _08046_);
  or (_14646_, _14645_, _08029_);
  and (_14647_, _14646_, _14643_);
  or (_14648_, _14647_, _08027_);
  nand (_14649_, _08027_, _02605_);
  and (_14650_, _14649_, _08067_);
  and (_14651_, _14650_, _08062_);
  and (_14652_, _14651_, _14648_);
  and (_14653_, _07224_, _07207_);
  nor (_14654_, _14653_, _07225_);
  and (_14655_, _14654_, _13285_);
  or (_14656_, _14655_, _07183_);
  or (_14657_, _14656_, _14652_);
  nor (_14658_, _07173_, _07157_);
  nor (_14659_, _14658_, _07174_);
  or (_14660_, _14659_, _08792_);
  and (_14661_, _14660_, _02857_);
  and (_14662_, _14661_, _14657_);
  nor (_14663_, _08090_, _08078_);
  nor (_14664_, _14663_, _08091_);
  or (_14665_, _14664_, _02441_);
  and (_14666_, _14665_, _08772_);
  or (_14667_, _14666_, _14662_);
  nor (_14668_, _08123_, _08110_);
  nor (_14669_, _14668_, _08124_);
  or (_14670_, _14669_, _08074_);
  and (_14671_, _14670_, _09650_);
  and (_14672_, _14671_, _14667_);
  and (_14673_, _07143_, \oc8051_golden_model_1.ACC [3]);
  or (_14674_, _14673_, _03133_);
  or (_14675_, _14674_, _14672_);
  nand (_14676_, _14426_, _03133_);
  and (_14677_, _14676_, _08139_);
  and (_14678_, _14677_, _14675_);
  and (_14679_, _08145_, _06814_);
  nor (_14680_, _08145_, _06814_);
  nor (_14681_, _14680_, _14679_);
  not (_14682_, _14681_);
  and (_14683_, _14682_, _08138_);
  or (_14684_, _14683_, _08143_);
  or (_14685_, _14684_, _14678_);
  nand (_14686_, _08143_, _06808_);
  and (_14687_, _14686_, _03142_);
  and (_14688_, _14687_, _14685_);
  nor (_14689_, _14472_, _03142_);
  or (_14690_, _14689_, _02852_);
  or (_14691_, _14690_, _14688_);
  and (_14692_, _11383_, _04654_);
  nor (_14693_, _14692_, _14413_);
  nand (_14694_, _14693_, _02852_);
  and (_14695_, _14694_, _08161_);
  and (_14696_, _14695_, _14691_);
  and (_14697_, _08169_, _06814_);
  nor (_14698_, _14697_, _08170_);
  and (_14699_, _14698_, _08160_);
  or (_14700_, _14699_, _08167_);
  or (_14701_, _14700_, _14696_);
  nand (_14702_, _08167_, _06808_);
  and (_14703_, _14702_, _34446_);
  and (_14704_, _14703_, _14701_);
  or (_14705_, _14704_, _14408_);
  and (_35614_[4], _14705_, _35583_);
  nor (_14706_, _34446_, _06808_);
  nor (_14707_, _04654_, _06808_);
  nor (_14708_, _11524_, _07325_);
  nor (_14709_, _14708_, _14707_);
  nor (_14710_, _14709_, _07120_);
  nand (_14711_, _14310_, _07201_);
  and (_14712_, _11525_, _04654_);
  nor (_14713_, _14712_, _14707_);
  nand (_14714_, _14713_, _02977_);
  or (_14715_, _07153_, _07833_);
  nor (_14716_, _07808_, _03179_);
  nor (_14717_, _04839_, _07325_);
  nor (_14718_, _14717_, _14707_);
  nand (_14719_, _14718_, _03861_);
  and (_14720_, _03620_, \oc8051_golden_model_1.ACC [4]);
  nor (_14721_, _14524_, _14720_);
  nor (_14722_, _08834_, _14721_);
  and (_14723_, _08834_, _14721_);
  nor (_14724_, _14723_, _14722_);
  and (_14725_, _14724_, \oc8051_golden_model_1.PSW [7]);
  nor (_14726_, _14724_, \oc8051_golden_model_1.PSW [7]);
  nor (_14727_, _14726_, _14725_);
  nor (_14728_, _14530_, _14527_);
  not (_14729_, _14728_);
  and (_14730_, _14729_, _14727_);
  nor (_14731_, _14729_, _14727_);
  nor (_14732_, _14731_, _14730_);
  or (_14733_, _14732_, _07541_);
  and (_14734_, _06072_, \oc8051_golden_model_1.ACC [4]);
  nor (_14735_, _14508_, _14734_);
  nor (_14736_, _14735_, _07154_);
  and (_14737_, _14735_, _07154_);
  nor (_14738_, _14737_, _14736_);
  nor (_14739_, _14738_, _07294_);
  and (_14740_, _14738_, _07294_);
  nor (_14741_, _14740_, _14739_);
  nor (_14742_, _14514_, _14511_);
  not (_14743_, _14742_);
  and (_14744_, _14743_, _14741_);
  nor (_14745_, _14743_, _14741_);
  nor (_14746_, _14745_, _14744_);
  and (_14747_, _14746_, _07329_);
  nor (_14748_, _05291_, _06808_);
  and (_14749_, _11422_, _05291_);
  and (_14750_, _14749_, _11437_);
  nor (_14751_, _14750_, _14748_);
  nor (_14752_, _14751_, _06189_);
  nand (_14753_, _07476_, _04839_);
  nor (_14754_, _11408_, _07325_);
  nor (_14755_, _14754_, _14707_);
  nand (_14756_, _14755_, _02932_);
  nor (_14757_, _07572_, _07406_);
  or (_14758_, _06120_, _07408_);
  not (_14759_, _07413_);
  nand (_14760_, _14759_, _04839_);
  nor (_14761_, _07415_, \oc8051_golden_model_1.ACC [5]);
  and (_14762_, _07415_, \oc8051_golden_model_1.ACC [5]);
  or (_14763_, _14762_, _14761_);
  nand (_14764_, _14763_, _09158_);
  and (_14765_, _14764_, _14760_);
  and (_14766_, _14765_, _07406_);
  and (_14767_, _14766_, _14758_);
  or (_14768_, _14767_, _14757_);
  and (_14769_, _14768_, _07429_);
  not (_14770_, \oc8051_golden_model_1.XRAM_DATA_IN [5]);
  nor (_14771_, _07433_, _14770_);
  or (_14772_, _14771_, _02932_);
  or (_14773_, _14772_, _14769_);
  and (_14774_, _14773_, _14756_);
  or (_14775_, _14774_, _07402_);
  and (_14776_, _09890_, _07449_);
  nor (_14777_, _09890_, _07449_);
  nor (_14778_, _14777_, _14776_);
  nand (_14779_, _14778_, _07402_);
  and (_14780_, _14779_, _02939_);
  and (_14781_, _14780_, _14775_);
  nor (_14782_, _14749_, _14748_);
  nor (_14783_, _14782_, _03186_);
  nor (_14784_, _14718_, _03693_);
  or (_14785_, _14784_, _07476_);
  or (_14786_, _14785_, _14783_);
  or (_14787_, _14786_, _14781_);
  and (_14788_, _14787_, _14753_);
  or (_14789_, _14788_, _03374_);
  or (_14790_, _06120_, _03375_);
  and (_14791_, _14790_, _02943_);
  and (_14792_, _14791_, _14789_);
  nor (_14793_, _07572_, _02943_);
  or (_14794_, _14793_, _07486_);
  or (_14795_, _14794_, _14792_);
  nand (_14796_, _07486_, _02477_);
  and (_14797_, _14796_, _14795_);
  or (_14798_, _14797_, _02796_);
  and (_14799_, _11405_, _05291_);
  nor (_14800_, _14799_, _14748_);
  nand (_14801_, _14800_, _02796_);
  and (_14802_, _14801_, _06189_);
  and (_14803_, _14802_, _14798_);
  or (_14804_, _14803_, _14752_);
  and (_14805_, _14804_, _06201_);
  nor (_14806_, _06668_, _06666_);
  nor (_14807_, _14806_, _06669_);
  and (_14808_, _14807_, _06195_);
  or (_14809_, _14808_, _07401_);
  or (_14810_, _14809_, _14805_);
  and (_14811_, _05143_, \oc8051_golden_model_1.ACC [4]);
  nor (_14812_, _14491_, _14811_);
  nor (_14813_, _14812_, _07202_);
  and (_14814_, _14812_, _07202_);
  nor (_14815_, _14814_, _14813_);
  and (_14816_, _14815_, \oc8051_golden_model_1.PSW [7]);
  nor (_14817_, _14815_, \oc8051_golden_model_1.PSW [7]);
  nor (_14818_, _14817_, _14816_);
  nor (_14819_, _14497_, _14494_);
  not (_14820_, _14819_);
  and (_14821_, _14820_, _14818_);
  nor (_14822_, _14820_, _14818_);
  nor (_14823_, _14822_, _14821_);
  or (_14824_, _14823_, _07400_);
  and (_14825_, _14824_, _07330_);
  and (_14826_, _14825_, _14810_);
  or (_14827_, _14826_, _14747_);
  and (_14828_, _14827_, _02899_);
  and (_14829_, _07690_, _07677_);
  nor (_14830_, _14829_, _07691_);
  nor (_14831_, _14830_, _02899_);
  or (_14832_, _14831_, _07540_);
  or (_14833_, _14832_, _14828_);
  and (_14834_, _14833_, _14733_);
  or (_14835_, _14834_, _07700_);
  nand (_14836_, _03179_, _07700_);
  and (_14837_, _14836_, _02966_);
  and (_14838_, _14837_, _14835_);
  nor (_14839_, _11455_, _07786_);
  nor (_14840_, _14839_, _14748_);
  nor (_14841_, _14840_, _02966_);
  or (_14842_, _14841_, _03861_);
  or (_14843_, _14842_, _14838_);
  and (_14844_, _14843_, _14719_);
  or (_14845_, _14844_, _03850_);
  and (_14846_, _06120_, _04654_);
  nor (_14847_, _14846_, _14707_);
  nand (_14848_, _14847_, _03850_);
  and (_14849_, _14848_, _02970_);
  and (_14850_, _14849_, _14845_);
  nor (_14851_, _11511_, _07325_);
  nor (_14852_, _14851_, _14707_);
  nor (_14853_, _14852_, _02970_);
  or (_14854_, _14853_, _06731_);
  or (_14855_, _14854_, _14850_);
  or (_14856_, _06793_, _06737_);
  and (_14857_, _14856_, _14855_);
  and (_14858_, _14857_, _02552_);
  nor (_14859_, _03179_, _02552_);
  or (_14860_, _14859_, _02974_);
  or (_14861_, _14860_, _14858_);
  and (_14862_, _05633_, _04654_);
  nor (_14863_, _14862_, _14707_);
  nand (_14864_, _14863_, _02974_);
  and (_14865_, _14864_, _07808_);
  and (_14866_, _14865_, _14861_);
  or (_14867_, _14866_, _14716_);
  and (_14868_, _14867_, _14118_);
  and (_14869_, _14276_, _07202_);
  nor (_14870_, _14869_, _14868_);
  nor (_14871_, _14870_, _08816_);
  and (_14872_, _07202_, _08816_);
  or (_14873_, _14872_, _14871_);
  and (_14874_, _14873_, _08820_);
  and (_14875_, _08819_, _07202_);
  or (_14876_, _14875_, _07832_);
  or (_14877_, _14876_, _14874_);
  and (_14878_, _14877_, _14715_);
  or (_14879_, _14878_, _03105_);
  or (_14880_, _11531_, _03106_);
  and (_14881_, _14880_, _07846_);
  and (_14882_, _14881_, _14879_);
  and (_14883_, _07319_, _08834_);
  or (_14884_, _14883_, _02977_);
  or (_14885_, _14884_, _14882_);
  and (_14886_, _14885_, _14714_);
  or (_14887_, _14886_, _03107_);
  or (_14888_, _14707_, _07104_);
  and (_14889_, _14888_, _07868_);
  and (_14890_, _14889_, _14887_);
  and (_14891_, _07869_, _07200_);
  or (_14892_, _14891_, _03499_);
  or (_14893_, _14892_, _14890_);
  or (_14894_, _07151_, _07876_);
  and (_14895_, _14894_, _03093_);
  and (_14896_, _14895_, _14893_);
  or (_14897_, _11529_, _07880_);
  and (_14898_, _14897_, _07882_);
  or (_14899_, _14898_, _14896_);
  or (_14900_, _07886_, _08106_);
  and (_14901_, _14900_, _03881_);
  and (_14902_, _14901_, _14899_);
  or (_14903_, _14863_, _11530_);
  nor (_14904_, _14903_, _03881_);
  or (_14905_, _14904_, _14310_);
  or (_14906_, _14905_, _14902_);
  and (_14907_, _14906_, _14711_);
  or (_14908_, _14907_, _14410_);
  nand (_14909_, _14410_, _07201_);
  and (_14910_, _14909_, _03525_);
  and (_14911_, _14910_, _14908_);
  nor (_14912_, _07201_, _03525_);
  or (_14913_, _14912_, _07315_);
  or (_14914_, _14913_, _14911_);
  nand (_14915_, _07152_, _07315_);
  and (_14916_, _14915_, _03098_);
  and (_14917_, _14916_, _14914_);
  nand (_14918_, _11530_, _07902_);
  and (_14919_, _14918_, _07901_);
  or (_14920_, _14919_, _14917_);
  nand (_14921_, _07899_, _08107_);
  and (_14922_, _14921_, _07120_);
  and (_14923_, _14922_, _14920_);
  or (_14924_, _14923_, _14710_);
  and (_14925_, _14924_, _07241_);
  and (_14926_, _07306_, _07263_);
  nor (_14927_, _14926_, _07307_);
  and (_14928_, _14927_, _07912_);
  or (_14929_, _14928_, _07236_);
  or (_14930_, _14929_, _14925_);
  and (_14931_, _07935_, _07358_);
  nor (_14932_, _14931_, _07936_);
  or (_14933_, _14932_, _07917_);
  and (_14934_, _14933_, _03104_);
  and (_14935_, _14934_, _14930_);
  and (_14936_, _08016_, _07980_);
  nor (_14937_, _14936_, _08017_);
  or (_14938_, _14937_, _07946_);
  and (_14939_, _14938_, _07948_);
  or (_14940_, _14939_, _14935_);
  and (_14941_, _08047_, _07726_);
  nor (_14942_, _14941_, _08048_);
  or (_14943_, _14942_, _08029_);
  and (_14944_, _14943_, _08028_);
  and (_14945_, _14944_, _14940_);
  and (_14946_, _08027_, \oc8051_golden_model_1.ACC [4]);
  nor (_14947_, _14946_, _07183_);
  nand (_14948_, _14947_, _07193_);
  or (_14949_, _14948_, _14945_);
  and (_14950_, _07175_, _07154_);
  nor (_14951_, _14950_, _07176_);
  or (_14952_, _14951_, _08792_);
  and (_14953_, _07226_, _07203_);
  nor (_14954_, _14953_, _07227_);
  or (_14955_, _14954_, _07193_);
  and (_14956_, _14955_, _03125_);
  and (_14957_, _14956_, _14952_);
  and (_14958_, _14957_, _14949_);
  and (_14959_, _08092_, _07674_);
  nor (_14960_, _14959_, _08093_);
  or (_14961_, _14960_, _02441_);
  and (_14962_, _14961_, _08772_);
  or (_14963_, _14962_, _14958_);
  not (_14964_, _08834_);
  nor (_14965_, _08125_, _14964_);
  and (_14966_, _08125_, _14964_);
  nor (_14967_, _14966_, _14965_);
  or (_14968_, _14967_, _08074_);
  and (_14969_, _14968_, _09650_);
  and (_14970_, _14969_, _14963_);
  and (_14971_, _07143_, \oc8051_golden_model_1.ACC [4]);
  or (_14972_, _14971_, _03133_);
  or (_14973_, _14972_, _14970_);
  nand (_14974_, _14755_, _03133_);
  and (_14975_, _14974_, _08139_);
  and (_14976_, _14975_, _14973_);
  nor (_14977_, _14679_, _06808_);
  or (_14978_, _14977_, _08146_);
  and (_14979_, _14978_, _08138_);
  or (_14980_, _14979_, _08143_);
  or (_14981_, _14980_, _14976_);
  nand (_14982_, _08143_, _06762_);
  and (_14983_, _14982_, _03142_);
  and (_14984_, _14983_, _14981_);
  nor (_14985_, _14800_, _03142_);
  or (_14986_, _14985_, _02852_);
  or (_14987_, _14986_, _14984_);
  and (_14988_, _11580_, _04654_);
  nor (_14989_, _14988_, _14707_);
  nand (_14990_, _14989_, _02852_);
  and (_14991_, _14990_, _08161_);
  and (_14992_, _14991_, _14987_);
  nor (_14993_, _08170_, \oc8051_golden_model_1.ACC [5]);
  nor (_14994_, _14993_, _08171_);
  and (_14995_, _14994_, _08160_);
  or (_14996_, _14995_, _08167_);
  or (_14997_, _14996_, _14992_);
  nand (_14998_, _08167_, _06762_);
  and (_14999_, _14998_, _34446_);
  and (_15000_, _14999_, _14997_);
  or (_15001_, _15000_, _14706_);
  and (_35614_[5], _15001_, _35583_);
  nor (_15002_, _34446_, _06762_);
  nand (_15003_, _07143_, _06808_);
  and (_15004_, _08094_, _07559_);
  nor (_15005_, _15004_, _08095_);
  or (_15006_, _15005_, _02857_);
  and (_15007_, _15006_, _08074_);
  nand (_15008_, _07899_, _08104_);
  nand (_15009_, _07317_, _07198_);
  not (_15010_, _07197_);
  nand (_15011_, _15010_, _03496_);
  nor (_15012_, _04654_, _06762_);
  and (_15013_, _11728_, _04654_);
  nor (_15014_, _15013_, _15012_);
  nand (_15015_, _15014_, _02977_);
  and (_15016_, _13667_, _07199_);
  nor (_15017_, _04735_, _07325_);
  nor (_15018_, _15017_, _15012_);
  nand (_15019_, _15018_, _03861_);
  and (_15020_, _07692_, _07673_);
  nor (_15021_, _15020_, _07693_);
  nand (_15022_, _15021_, _02898_);
  and (_15023_, _15022_, _07541_);
  or (_15024_, _06120_, _06808_);
  and (_15025_, _06120_, _06808_);
  or (_15026_, _14735_, _15025_);
  and (_15027_, _15026_, _15024_);
  nor (_15028_, _15027_, _07150_);
  and (_15029_, _15027_, _07150_);
  nor (_15030_, _15029_, _15028_);
  nor (_15031_, _14744_, _14739_);
  and (_15032_, _15031_, \oc8051_golden_model_1.PSW [7]);
  nor (_15033_, _15032_, _15030_);
  and (_15034_, _15032_, _15030_);
  nor (_15035_, _15034_, _15033_);
  and (_15036_, _15035_, _07329_);
  nand (_15037_, _07476_, _04735_);
  nor (_15038_, _11610_, _07325_);
  nor (_15039_, _15038_, _15012_);
  nand (_15040_, _15039_, _02932_);
  nor (_15041_, _07556_, _07406_);
  or (_15042_, _05798_, _07408_);
  nor (_15043_, _07413_, _04735_);
  and (_15044_, _07415_, _06762_);
  nor (_15045_, _07415_, _06762_);
  or (_15046_, _15045_, _03343_);
  or (_15047_, _15046_, _15044_);
  and (_15048_, _15047_, _07413_);
  or (_15049_, _15048_, _15043_);
  and (_15050_, _15049_, _07406_);
  and (_15051_, _15050_, _15042_);
  or (_15052_, _15051_, _15041_);
  and (_15053_, _15052_, _07429_);
  and (_15054_, _07434_, \oc8051_golden_model_1.XRAM_DATA_IN [6]);
  or (_15055_, _15054_, _02932_);
  or (_15056_, _15055_, _15053_);
  and (_15057_, _15056_, _15040_);
  or (_15058_, _15057_, _07402_);
  not (_15059_, _07451_);
  nor (_15060_, _14777_, _15059_);
  and (_15061_, _09889_, _07452_);
  nor (_15062_, _15061_, _15060_);
  nand (_15063_, _15062_, _07402_);
  and (_15064_, _15063_, _02939_);
  and (_15065_, _15064_, _15058_);
  nor (_15066_, _05291_, _06762_);
  and (_15067_, _11604_, _05291_);
  nor (_15068_, _15067_, _15066_);
  nor (_15069_, _15068_, _03186_);
  nor (_15070_, _15018_, _03693_);
  or (_15071_, _15070_, _07476_);
  or (_15072_, _15071_, _15069_);
  or (_15073_, _15072_, _15065_);
  and (_15074_, _15073_, _15037_);
  or (_15075_, _15074_, _03374_);
  or (_15076_, _05798_, _03375_);
  and (_15077_, _15076_, _02943_);
  and (_15078_, _15077_, _15075_);
  nor (_15079_, _07556_, _02943_);
  or (_15080_, _15079_, _07486_);
  or (_15081_, _15080_, _15078_);
  nand (_15083_, _07486_, _06908_);
  and (_15084_, _15083_, _15081_);
  or (_15085_, _15084_, _02796_);
  and (_15086_, _11633_, _05291_);
  nor (_15087_, _15086_, _15066_);
  nand (_15088_, _15087_, _02796_);
  and (_15089_, _15088_, _06189_);
  and (_15090_, _15089_, _15085_);
  and (_15091_, _15067_, _11603_);
  nor (_15092_, _15091_, _15066_);
  nor (_15094_, _15092_, _06189_);
  or (_15095_, _15094_, _06195_);
  or (_15096_, _15095_, _15090_);
  nor (_15097_, _06671_, _06669_);
  nor (_15098_, _15097_, _06672_);
  or (_15099_, _15098_, _06201_);
  and (_15100_, _15099_, _15096_);
  or (_15101_, _15100_, _07401_);
  nand (_15102_, _04839_, \oc8051_golden_model_1.ACC [5]);
  nor (_15103_, _04839_, \oc8051_golden_model_1.ACC [5]);
  or (_15105_, _14812_, _15103_);
  and (_15106_, _15105_, _15102_);
  nor (_15107_, _15106_, _07199_);
  and (_15108_, _15106_, _07199_);
  nor (_15109_, _15108_, _15107_);
  nor (_15110_, _14821_, _14816_);
  and (_15111_, _15110_, \oc8051_golden_model_1.PSW [7]);
  nor (_15112_, _15111_, _15109_);
  and (_15113_, _15111_, _15109_);
  nor (_15114_, _15113_, _15112_);
  or (_15116_, _15114_, _07400_);
  and (_15117_, _15116_, _07330_);
  and (_15118_, _15117_, _15101_);
  or (_15119_, _15118_, _02898_);
  or (_15120_, _15119_, _15036_);
  and (_15121_, _15120_, _15023_);
  or (_15122_, _14721_, _09952_);
  and (_15123_, _15122_, _09951_);
  nor (_15124_, _15123_, _08105_);
  and (_15125_, _15123_, _08105_);
  nor (_15127_, _15125_, _15124_);
  nor (_15128_, _14730_, _14725_);
  and (_15129_, _15128_, \oc8051_golden_model_1.PSW [7]);
  nor (_15130_, _15129_, _15127_);
  and (_15131_, _15129_, _15127_);
  nor (_15132_, _15131_, _15130_);
  and (_15133_, _15132_, _07540_);
  or (_15134_, _15133_, _07700_);
  or (_15135_, _15134_, _15121_);
  nand (_15136_, _02889_, _07700_);
  and (_15138_, _15136_, _02966_);
  and (_15139_, _15138_, _15135_);
  nor (_15140_, _11655_, _07786_);
  nor (_15141_, _15140_, _15066_);
  nor (_15142_, _15141_, _02966_);
  or (_15143_, _15142_, _03861_);
  or (_15144_, _15143_, _15139_);
  and (_15145_, _15144_, _15019_);
  or (_15146_, _15145_, _03850_);
  and (_15147_, _05798_, _04654_);
  nor (_15149_, _15147_, _15012_);
  nand (_15150_, _15149_, _03850_);
  and (_15151_, _15150_, _02970_);
  and (_15152_, _15151_, _15146_);
  nor (_15153_, _11711_, _07325_);
  nor (_15154_, _15153_, _15012_);
  nor (_15155_, _15154_, _02970_);
  or (_15156_, _15155_, _06731_);
  or (_15157_, _15156_, _15152_);
  not (_15158_, _06763_);
  and (_15160_, _06767_, _15158_);
  or (_15161_, _15160_, _06737_);
  and (_15162_, _15161_, _15157_);
  and (_15163_, _15162_, _02552_);
  nor (_15164_, _02889_, _02552_);
  or (_15165_, _15164_, _02974_);
  or (_15166_, _15165_, _15163_);
  and (_15167_, _11718_, _04654_);
  nor (_15168_, _15167_, _15012_);
  nand (_15169_, _15168_, _02974_);
  and (_15171_, _15169_, _07808_);
  and (_15172_, _15171_, _15166_);
  nor (_15173_, _07808_, _02889_);
  or (_15174_, _15173_, _07817_);
  or (_15175_, _15174_, _15172_);
  or (_15176_, _07816_, _07199_);
  and (_15177_, _15176_, _13666_);
  and (_15178_, _15177_, _15175_);
  or (_15179_, _15178_, _15016_);
  and (_15180_, _15179_, _13418_);
  and (_15182_, _13417_, _07150_);
  or (_15183_, _15182_, _15180_);
  and (_15184_, _15183_, _03487_);
  and (_15185_, _07150_, _03486_);
  or (_15186_, _15185_, _03105_);
  or (_15187_, _15186_, _15184_);
  or (_15188_, _11601_, _03106_);
  and (_15189_, _15188_, _07846_);
  and (_15190_, _15189_, _15187_);
  and (_15191_, _07319_, _08105_);
  or (_15193_, _15191_, _02977_);
  or (_15194_, _15193_, _15190_);
  and (_15195_, _15194_, _15015_);
  or (_15196_, _15195_, _03107_);
  nand (_15197_, _03680_, _02593_);
  and (_15198_, _07865_, _15197_);
  or (_15199_, _15012_, _07104_);
  and (_15200_, _15199_, _15198_);
  and (_15201_, _15200_, _15196_);
  nor (_15202_, _15198_, _15010_);
  or (_15204_, _15202_, _15201_);
  or (_15205_, _15204_, _03496_);
  and (_15206_, _15205_, _15011_);
  or (_15207_, _15206_, _03499_);
  or (_15208_, _07148_, _07876_);
  and (_15209_, _15208_, _03093_);
  and (_15210_, _15209_, _15207_);
  or (_15211_, _11599_, _07880_);
  and (_15212_, _15211_, _07882_);
  or (_15213_, _15212_, _15210_);
  or (_15215_, _07886_, _08103_);
  and (_15216_, _15215_, _03881_);
  and (_15217_, _15216_, _15213_);
  or (_15218_, _15168_, _11600_);
  nor (_15219_, _15218_, _03881_);
  or (_15220_, _15219_, _07317_);
  or (_15221_, _15220_, _15217_);
  and (_15222_, _15221_, _15009_);
  or (_15223_, _15222_, _07315_);
  nand (_15224_, _07149_, _07315_);
  and (_15226_, _15224_, _03098_);
  and (_15227_, _15226_, _15223_);
  nand (_15228_, _11600_, _07902_);
  and (_15229_, _15228_, _07901_);
  or (_15230_, _15229_, _15227_);
  and (_15231_, _15230_, _15008_);
  or (_15232_, _15231_, _02994_);
  nor (_15233_, _11726_, _07325_);
  nor (_15234_, _15233_, _15012_);
  nand (_15235_, _15234_, _02994_);
  and (_15237_, _15235_, _07241_);
  and (_15238_, _15237_, _15232_);
  and (_15239_, _07308_, _07256_);
  nor (_15240_, _15239_, _07309_);
  and (_15241_, _15240_, _07912_);
  or (_15242_, _15241_, _07236_);
  or (_15243_, _15242_, _15238_);
  and (_15244_, _07937_, _07919_);
  nor (_15245_, _15244_, _07938_);
  or (_15246_, _15245_, _07917_);
  and (_15248_, _15246_, _15243_);
  or (_15249_, _15248_, _03103_);
  and (_15250_, _08018_, _07971_);
  nor (_15251_, _15250_, _08019_);
  or (_15252_, _15251_, _03104_);
  and (_15253_, _15252_, _08029_);
  and (_15254_, _15253_, _15249_);
  and (_15255_, _08049_, _08031_);
  nor (_15256_, _15255_, _08050_);
  and (_15257_, _15256_, _07946_);
  or (_15258_, _15257_, _08027_);
  or (_15259_, _15258_, _15254_);
  nand (_15260_, _08027_, _06808_);
  and (_15261_, _15260_, _08795_);
  and (_15262_, _15261_, _15259_);
  nor (_15263_, _07177_, _07150_);
  nor (_15264_, _15263_, _07178_);
  and (_15265_, _15264_, _07183_);
  nor (_15266_, _07228_, _07199_);
  nor (_15267_, _15266_, _07229_);
  and (_15269_, _15267_, _13285_);
  or (_15270_, _15269_, _03124_);
  or (_15271_, _15270_, _15265_);
  or (_15272_, _15271_, _15262_);
  and (_15273_, _15272_, _15007_);
  nor (_15274_, _08127_, _08105_);
  nor (_15275_, _15274_, _08128_);
  and (_15276_, _15275_, _08073_);
  or (_15277_, _15276_, _07143_);
  or (_15278_, _15277_, _15273_);
  and (_15280_, _15278_, _15003_);
  or (_15281_, _15280_, _03133_);
  nand (_15282_, _15039_, _03133_);
  and (_15283_, _15282_, _08139_);
  and (_15284_, _15283_, _15281_);
  nor (_15285_, _08146_, _06762_);
  or (_15286_, _15285_, _08147_);
  and (_15287_, _15286_, _08138_);
  or (_15288_, _15287_, _08143_);
  or (_15289_, _15288_, _15284_);
  nand (_15291_, _08143_, _05719_);
  and (_15292_, _15291_, _03142_);
  and (_15293_, _15292_, _15289_);
  nor (_15294_, _15087_, _03142_);
  or (_15295_, _15294_, _02852_);
  or (_15296_, _15295_, _15293_);
  and (_15297_, _11778_, _04654_);
  nor (_15298_, _15297_, _15012_);
  nand (_15299_, _15298_, _02852_);
  and (_15300_, _15299_, _08161_);
  and (_15302_, _15300_, _15296_);
  nor (_15303_, _08171_, \oc8051_golden_model_1.ACC [6]);
  nor (_15304_, _15303_, _08172_);
  nor (_15305_, _15304_, _08167_);
  nor (_15306_, _15305_, _09696_);
  or (_15307_, _15306_, _15302_);
  nand (_15308_, _08167_, _05719_);
  and (_15309_, _15308_, _34446_);
  and (_15310_, _15309_, _15307_);
  or (_15311_, _15310_, _15002_);
  and (_35614_[6], _15311_, _35583_);
  not (_15313_, \oc8051_golden_model_1.DPL [0]);
  nor (_15314_, _34446_, _15313_);
  nor (_15315_, _04670_, _15313_);
  and (_15316_, _04670_, _03805_);
  or (_15317_, _15316_, _15315_);
  or (_15318_, _15317_, _03860_);
  and (_15319_, _04670_, \oc8051_golden_model_1.ACC [0]);
  or (_15320_, _15319_, _15315_);
  or (_15321_, _15320_, _02943_);
  nor (_15323_, _05036_, _08190_);
  or (_15324_, _15323_, _15315_);
  or (_15325_, _15324_, _06162_);
  and (_15326_, _15320_, _02837_);
  nor (_15327_, _02837_, _15313_);
  or (_15328_, _15327_, _02932_);
  or (_15329_, _15328_, _15326_);
  and (_15330_, _15329_, _03693_);
  and (_15331_, _15330_, _15325_);
  and (_15332_, _15317_, _02930_);
  or (_15334_, _15332_, _02928_);
  or (_15335_, _15334_, _15331_);
  and (_15336_, _15335_, _15321_);
  or (_15337_, _15336_, _08209_);
  and (_15338_, _08209_, \oc8051_golden_model_1.DPL [0]);
  nor (_15339_, _15338_, _02975_);
  and (_15340_, _15339_, _15337_);
  nor (_15341_, _03471_, _08194_);
  or (_15342_, _15341_, _03861_);
  or (_15343_, _15342_, _15340_);
  and (_15345_, _15343_, _15318_);
  or (_15346_, _15345_, _03850_);
  and (_15347_, _06114_, _04670_);
  or (_15348_, _15315_, _06726_);
  or (_15349_, _15348_, _15347_);
  and (_15350_, _15349_, _15346_);
  or (_15351_, _15350_, _02524_);
  nor (_15352_, _10530_, _08190_);
  or (_15353_, _15315_, _02970_);
  or (_15354_, _15353_, _15352_);
  and (_15356_, _15354_, _05261_);
  and (_15357_, _15356_, _15351_);
  and (_15358_, _04670_, _05647_);
  or (_15359_, _15358_, _15315_);
  and (_15360_, _15359_, _02974_);
  or (_15361_, _15360_, _02977_);
  or (_15362_, _15361_, _15357_);
  and (_15363_, _10427_, _04670_);
  or (_15364_, _15363_, _15315_);
  or (_15365_, _15364_, _07092_);
  and (_15367_, _15365_, _15362_);
  or (_15368_, _15367_, _03107_);
  and (_15369_, _10546_, _04670_);
  or (_15370_, _15315_, _07104_);
  or (_15371_, _15370_, _15369_);
  and (_15372_, _15371_, _03881_);
  and (_15373_, _15372_, _15368_);
  nand (_15374_, _15359_, _02991_);
  nor (_15375_, _15374_, _15323_);
  or (_15376_, _15375_, _15373_);
  and (_15378_, _15376_, _06161_);
  or (_15379_, _15315_, _05036_);
  and (_15380_, _15320_, _03094_);
  and (_15381_, _15380_, _15379_);
  or (_15382_, _15381_, _02994_);
  or (_15383_, _15382_, _15378_);
  nor (_15384_, _10425_, _08190_);
  or (_15385_, _15315_, _07120_);
  or (_15386_, _15385_, _15384_);
  and (_15387_, _15386_, _07118_);
  and (_15389_, _15387_, _15383_);
  not (_15390_, _03330_);
  nor (_15391_, _10423_, _08190_);
  or (_15392_, _15391_, _15315_);
  and (_15393_, _15392_, _03099_);
  or (_15394_, _15393_, _15390_);
  or (_15395_, _15394_, _15389_);
  or (_15396_, _15324_, _03330_);
  and (_15397_, _15396_, _34446_);
  and (_15398_, _15397_, _15395_);
  or (_15400_, _15398_, _15314_);
  and (_35617_[0], _15400_, _35583_);
  not (_15401_, \oc8051_golden_model_1.DPL [1]);
  nor (_15402_, _34446_, _15401_);
  nand (_15403_, _04670_, _03660_);
  or (_15404_, _04670_, \oc8051_golden_model_1.DPL [1]);
  and (_15405_, _15404_, _02974_);
  and (_15406_, _15405_, _15403_);
  nand (_15407_, _10719_, _04670_);
  and (_15408_, _15404_, _02524_);
  and (_15410_, _15408_, _15407_);
  nor (_15411_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor (_15412_, _15411_, _08214_);
  and (_15413_, _15412_, _08209_);
  and (_15414_, _10622_, _04670_);
  not (_15415_, _15414_);
  and (_15416_, _15415_, _15404_);
  or (_15417_, _15416_, _06162_);
  nand (_15418_, _04670_, _02477_);
  and (_15419_, _15418_, _15404_);
  and (_15421_, _15419_, _02837_);
  nor (_15422_, _02837_, _15401_);
  or (_15423_, _15422_, _02932_);
  or (_15424_, _15423_, _15421_);
  and (_15425_, _15424_, _03693_);
  and (_15426_, _15425_, _15417_);
  nor (_15427_, _04670_, _15401_);
  nor (_15428_, _08190_, _03989_);
  or (_15429_, _15428_, _15427_);
  and (_15430_, _15429_, _02930_);
  or (_15432_, _15430_, _02928_);
  or (_15433_, _15432_, _15426_);
  or (_15434_, _15419_, _02943_);
  and (_15435_, _15434_, _08210_);
  and (_15436_, _15435_, _15433_);
  or (_15437_, _15436_, _15413_);
  and (_15438_, _15437_, _08194_);
  nor (_15439_, _03660_, _08194_);
  or (_15440_, _15439_, _03861_);
  or (_15441_, _15440_, _15438_);
  or (_15443_, _15429_, _03860_);
  and (_15444_, _15443_, _15441_);
  or (_15445_, _15444_, _03850_);
  and (_15446_, _06113_, _04670_);
  or (_15447_, _15427_, _06726_);
  or (_15448_, _15447_, _15446_);
  and (_15449_, _15448_, _02970_);
  and (_15450_, _15449_, _15445_);
  or (_15451_, _15450_, _15410_);
  and (_15452_, _15451_, _05261_);
  or (_15454_, _15452_, _15406_);
  and (_15455_, _15454_, _03882_);
  or (_15456_, _10613_, _08190_);
  and (_15457_, _15404_, _02991_);
  and (_15458_, _15457_, _15456_);
  or (_15459_, _10610_, _08190_);
  and (_15460_, _15404_, _03107_);
  and (_15461_, _15460_, _15459_);
  or (_15462_, _10614_, _08190_);
  and (_15463_, _15404_, _02977_);
  and (_15465_, _15463_, _15462_);
  or (_15466_, _15465_, _15461_);
  or (_15467_, _15466_, _15458_);
  or (_15468_, _15467_, _15455_);
  and (_15469_, _15468_, _06161_);
  or (_15470_, _15427_, _04988_);
  and (_15471_, _15419_, _03094_);
  and (_15472_, _15471_, _15470_);
  or (_15473_, _15472_, _15469_);
  and (_15474_, _15473_, _03100_);
  or (_15476_, _15403_, _04988_);
  and (_15477_, _15404_, _02994_);
  and (_15478_, _15477_, _15476_);
  or (_15479_, _15418_, _04988_);
  and (_15480_, _15404_, _03099_);
  and (_15481_, _15480_, _15479_);
  or (_15482_, _15481_, _03133_);
  or (_15483_, _15482_, _15478_);
  or (_15484_, _15483_, _15474_);
  or (_15485_, _15416_, _03138_);
  and (_15487_, _15485_, _15484_);
  or (_15488_, _15487_, _02852_);
  or (_15489_, _15427_, _02853_);
  or (_15490_, _15489_, _15414_);
  and (_15491_, _15490_, _34446_);
  and (_15492_, _15491_, _15488_);
  or (_15493_, _15492_, _15402_);
  and (_35617_[1], _15493_, _35583_);
  or (_15494_, _34446_, \oc8051_golden_model_1.DPL [2]);
  and (_15495_, _15494_, _35583_);
  not (_15497_, \oc8051_golden_model_1.DPL [2]);
  nor (_15498_, _04670_, _15497_);
  and (_15499_, _10942_, _04670_);
  or (_15500_, _15499_, _15498_);
  and (_15501_, _15500_, _03107_);
  nor (_15502_, _08190_, _04413_);
  or (_15503_, _15502_, _15498_);
  or (_15504_, _15503_, _03860_);
  or (_15505_, _15503_, _03693_);
  nor (_15506_, _10824_, _08190_);
  or (_15508_, _15506_, _15498_);
  and (_15509_, _15508_, _02932_);
  nor (_15510_, _02837_, _15497_);
  and (_15511_, _04670_, \oc8051_golden_model_1.ACC [2]);
  or (_15512_, _15511_, _15498_);
  and (_15513_, _15512_, _02837_);
  or (_15514_, _15513_, _15510_);
  and (_15515_, _15514_, _06162_);
  or (_15516_, _15515_, _02930_);
  or (_15517_, _15516_, _15509_);
  and (_15519_, _15517_, _15505_);
  or (_15520_, _15519_, _02928_);
  or (_15521_, _15512_, _02943_);
  and (_15522_, _15521_, _08210_);
  and (_15523_, _15522_, _15520_);
  nor (_15524_, _08214_, \oc8051_golden_model_1.DPL [2]);
  nor (_15525_, _15524_, _08215_);
  and (_15526_, _15525_, _08209_);
  or (_15527_, _15526_, _15523_);
  and (_15528_, _15527_, _08194_);
  nor (_15530_, _03223_, _08194_);
  or (_15531_, _15530_, _03861_);
  or (_15532_, _15531_, _15528_);
  and (_15533_, _15532_, _15504_);
  or (_15534_, _15533_, _03850_);
  and (_15535_, _06117_, _04670_);
  or (_15536_, _15498_, _06726_);
  or (_15537_, _15536_, _15535_);
  and (_15538_, _15537_, _02970_);
  and (_15539_, _15538_, _15534_);
  nor (_15541_, _10922_, _08190_);
  or (_15542_, _15541_, _15498_);
  and (_15543_, _15542_, _02524_);
  or (_15544_, _15543_, _02974_);
  or (_15545_, _15544_, _15539_);
  and (_15546_, _04670_, _05690_);
  or (_15547_, _15546_, _15498_);
  or (_15548_, _15547_, _05261_);
  and (_15549_, _15548_, _15545_);
  or (_15550_, _15549_, _02977_);
  and (_15552_, _10936_, _04670_);
  or (_15553_, _15498_, _07092_);
  or (_15554_, _15553_, _15552_);
  and (_15555_, _15554_, _07104_);
  and (_15556_, _15555_, _15550_);
  or (_15557_, _15556_, _15501_);
  and (_15558_, _15557_, _03095_);
  or (_15559_, _15498_, _05086_);
  and (_15560_, _15512_, _03094_);
  and (_15561_, _15547_, _02991_);
  or (_15563_, _15561_, _15560_);
  and (_15564_, _15563_, _15559_);
  or (_15565_, _15564_, _02994_);
  or (_15566_, _15565_, _15558_);
  nor (_15567_, _10935_, _08190_);
  or (_15568_, _15498_, _07120_);
  or (_15569_, _15568_, _15567_);
  and (_15570_, _15569_, _07118_);
  and (_15571_, _15570_, _15566_);
  nor (_15572_, _10941_, _08190_);
  or (_15574_, _15572_, _15498_);
  and (_15575_, _15574_, _03099_);
  or (_15576_, _15575_, _03133_);
  or (_15577_, _15576_, _15571_);
  or (_15578_, _15508_, _03138_);
  and (_15579_, _15578_, _02853_);
  and (_15580_, _15579_, _15577_);
  and (_15581_, _10988_, _04670_);
  or (_15582_, _15581_, _15498_);
  and (_15583_, _15582_, _02852_);
  or (_15585_, _15583_, _34450_);
  or (_15586_, _15585_, _15580_);
  and (_35617_[2], _15586_, _15495_);
  or (_15587_, _34446_, \oc8051_golden_model_1.DPL [3]);
  and (_15588_, _15587_, _35583_);
  and (_15589_, _08190_, \oc8051_golden_model_1.DPL [3]);
  and (_15590_, _11134_, _04670_);
  or (_15591_, _15590_, _15589_);
  and (_15592_, _15591_, _03107_);
  nor (_15593_, _08190_, _04226_);
  or (_15595_, _15593_, _15589_);
  or (_15596_, _15595_, _03860_);
  nor (_15597_, _08215_, \oc8051_golden_model_1.DPL [3]);
  nor (_15598_, _15597_, _08216_);
  and (_15599_, _15598_, _08209_);
  nor (_15600_, _11014_, _08190_);
  or (_15601_, _15600_, _15589_);
  or (_15602_, _15601_, _06162_);
  and (_15603_, _04670_, \oc8051_golden_model_1.ACC [3]);
  or (_15604_, _15603_, _15589_);
  and (_15606_, _15604_, _02837_);
  and (_15607_, _09167_, \oc8051_golden_model_1.DPL [3]);
  or (_15608_, _15607_, _02932_);
  or (_15609_, _15608_, _15606_);
  and (_15610_, _15609_, _03693_);
  and (_15611_, _15610_, _15602_);
  and (_15612_, _15595_, _02930_);
  or (_15613_, _15612_, _02928_);
  or (_15614_, _15613_, _15611_);
  or (_15615_, _15604_, _02943_);
  and (_15617_, _15615_, _08210_);
  and (_15618_, _15617_, _15614_);
  or (_15619_, _15618_, _15599_);
  and (_15620_, _15619_, _08194_);
  nor (_15621_, _03087_, _08194_);
  or (_15622_, _15621_, _03861_);
  or (_15623_, _15622_, _15620_);
  and (_15624_, _15623_, _15596_);
  or (_15625_, _15624_, _03850_);
  and (_15626_, _06116_, _04670_);
  or (_15628_, _15589_, _06726_);
  or (_15629_, _15628_, _15626_);
  and (_15630_, _15629_, _02970_);
  and (_15631_, _15630_, _15625_);
  nor (_15632_, _11114_, _08190_);
  or (_15633_, _15632_, _15589_);
  and (_15634_, _15633_, _02524_);
  or (_15635_, _15634_, _02974_);
  or (_15636_, _15635_, _15631_);
  and (_15637_, _04670_, _05616_);
  or (_15639_, _15637_, _15589_);
  or (_15640_, _15639_, _05261_);
  and (_15641_, _15640_, _15636_);
  or (_15642_, _15641_, _02977_);
  and (_15643_, _11128_, _04670_);
  or (_15644_, _15589_, _07092_);
  or (_15645_, _15644_, _15643_);
  and (_15646_, _15645_, _07104_);
  and (_15647_, _15646_, _15642_);
  or (_15648_, _15647_, _15592_);
  and (_15650_, _15648_, _03095_);
  or (_15651_, _15589_, _04939_);
  and (_15652_, _15604_, _03094_);
  and (_15653_, _15639_, _02991_);
  or (_15654_, _15653_, _15652_);
  and (_15655_, _15654_, _15651_);
  or (_15656_, _15655_, _02994_);
  or (_15657_, _15656_, _15650_);
  nor (_15658_, _11127_, _08190_);
  or (_15659_, _15589_, _07120_);
  or (_15661_, _15659_, _15658_);
  and (_15662_, _15661_, _07118_);
  and (_15663_, _15662_, _15657_);
  nor (_15664_, _11133_, _08190_);
  or (_15665_, _15664_, _15589_);
  and (_15666_, _15665_, _03099_);
  or (_15667_, _15666_, _03133_);
  or (_15668_, _15667_, _15663_);
  or (_15669_, _15601_, _03138_);
  and (_15670_, _15669_, _02853_);
  and (_15672_, _15670_, _15668_);
  and (_15673_, _11185_, _04670_);
  or (_15674_, _15673_, _15589_);
  and (_15675_, _15674_, _02852_);
  or (_15676_, _15675_, _34450_);
  or (_15677_, _15676_, _15672_);
  and (_35617_[3], _15677_, _15588_);
  or (_15678_, _34446_, \oc8051_golden_model_1.DPL [4]);
  and (_15679_, _15678_, _35583_);
  and (_15680_, _08190_, \oc8051_golden_model_1.DPL [4]);
  and (_15682_, _11333_, _04670_);
  or (_15683_, _15682_, _15680_);
  and (_15684_, _15683_, _03107_);
  nor (_15685_, _05143_, _08190_);
  or (_15686_, _15685_, _15680_);
  or (_15687_, _15686_, _03860_);
  nor (_15688_, _11207_, _08190_);
  or (_15689_, _15688_, _15680_);
  or (_15690_, _15689_, _06162_);
  and (_15691_, _04670_, \oc8051_golden_model_1.ACC [4]);
  or (_15693_, _15691_, _15680_);
  and (_15694_, _15693_, _02837_);
  and (_15695_, _09167_, \oc8051_golden_model_1.DPL [4]);
  or (_15696_, _15695_, _02932_);
  or (_15697_, _15696_, _15694_);
  and (_15698_, _15697_, _03693_);
  and (_15699_, _15698_, _15690_);
  and (_15700_, _15686_, _02930_);
  or (_15701_, _15700_, _02928_);
  or (_15702_, _15701_, _15699_);
  or (_15704_, _15693_, _02943_);
  and (_15705_, _15704_, _08210_);
  and (_15706_, _15705_, _15702_);
  nor (_15707_, _08216_, \oc8051_golden_model_1.DPL [4]);
  nor (_15708_, _15707_, _08217_);
  and (_15709_, _15708_, _08209_);
  or (_15710_, _15709_, _15706_);
  and (_15711_, _15710_, _08194_);
  nor (_15712_, _05581_, _08194_);
  or (_15713_, _15712_, _03861_);
  or (_15715_, _15713_, _15711_);
  and (_15716_, _15715_, _15687_);
  or (_15717_, _15716_, _03850_);
  and (_15718_, _06121_, _04670_);
  or (_15719_, _15680_, _06726_);
  or (_15720_, _15719_, _15718_);
  and (_15721_, _15720_, _02970_);
  and (_15722_, _15721_, _15717_);
  nor (_15723_, _11313_, _08190_);
  or (_15724_, _15723_, _15680_);
  and (_15726_, _15724_, _02524_);
  or (_15727_, _15726_, _02974_);
  or (_15728_, _15727_, _15722_);
  and (_15729_, _05629_, _04670_);
  or (_15730_, _15729_, _15680_);
  or (_15731_, _15730_, _05261_);
  and (_15732_, _15731_, _15728_);
  or (_15733_, _15732_, _02977_);
  and (_15734_, _11327_, _04670_);
  or (_15735_, _15680_, _07092_);
  or (_15737_, _15735_, _15734_);
  and (_15738_, _15737_, _07104_);
  and (_15739_, _15738_, _15733_);
  or (_15740_, _15739_, _15684_);
  and (_15741_, _15740_, _03095_);
  or (_15742_, _15680_, _05190_);
  and (_15743_, _15693_, _03094_);
  and (_15744_, _15730_, _02991_);
  or (_15745_, _15744_, _15743_);
  and (_15746_, _15745_, _15742_);
  or (_15748_, _15746_, _02994_);
  or (_15749_, _15748_, _15741_);
  nor (_15750_, _11326_, _08190_);
  or (_15751_, _15680_, _07120_);
  or (_15752_, _15751_, _15750_);
  and (_15753_, _15752_, _07118_);
  and (_15754_, _15753_, _15749_);
  nor (_15755_, _11332_, _08190_);
  or (_15756_, _15755_, _15680_);
  and (_15757_, _15756_, _03099_);
  or (_15759_, _15757_, _03133_);
  or (_15760_, _15759_, _15754_);
  or (_15761_, _15689_, _03138_);
  and (_15762_, _15761_, _02853_);
  and (_15763_, _15762_, _15760_);
  and (_15764_, _11383_, _04670_);
  or (_15765_, _15764_, _15680_);
  and (_15766_, _15765_, _02852_);
  or (_15767_, _15766_, _34450_);
  or (_15768_, _15767_, _15763_);
  and (_35617_[4], _15768_, _15679_);
  or (_15770_, _34446_, \oc8051_golden_model_1.DPL [5]);
  and (_15771_, _15770_, _35583_);
  and (_15772_, _08190_, \oc8051_golden_model_1.DPL [5]);
  and (_15773_, _11531_, _04670_);
  or (_15774_, _15773_, _15772_);
  and (_15775_, _15774_, _03107_);
  nor (_15776_, _04839_, _08190_);
  or (_15777_, _15776_, _15772_);
  or (_15778_, _15777_, _03860_);
  nor (_15780_, _11408_, _08190_);
  or (_15781_, _15780_, _15772_);
  or (_15782_, _15781_, _06162_);
  and (_15783_, _04670_, \oc8051_golden_model_1.ACC [5]);
  or (_15784_, _15783_, _15772_);
  and (_15785_, _15784_, _02837_);
  and (_15786_, _09167_, \oc8051_golden_model_1.DPL [5]);
  or (_15787_, _15786_, _02932_);
  or (_15788_, _15787_, _15785_);
  and (_15789_, _15788_, _03693_);
  and (_15791_, _15789_, _15782_);
  and (_15792_, _15777_, _02930_);
  or (_15793_, _15792_, _02928_);
  or (_15794_, _15793_, _15791_);
  or (_15795_, _15784_, _02943_);
  and (_15796_, _15795_, _08210_);
  and (_15797_, _15796_, _15794_);
  nor (_15798_, _08217_, \oc8051_golden_model_1.DPL [5]);
  nor (_15799_, _15798_, _08218_);
  and (_15800_, _15799_, _08209_);
  or (_15802_, _15800_, _15797_);
  and (_15803_, _15802_, _08194_);
  nor (_15804_, _05612_, _08194_);
  or (_15805_, _15804_, _03861_);
  or (_15806_, _15805_, _15803_);
  and (_15807_, _15806_, _15778_);
  or (_15808_, _15807_, _03850_);
  and (_15809_, _06120_, _04670_);
  or (_15810_, _15772_, _06726_);
  or (_15811_, _15810_, _15809_);
  and (_15813_, _15811_, _02970_);
  and (_15814_, _15813_, _15808_);
  nor (_15815_, _11511_, _08190_);
  or (_15816_, _15815_, _15772_);
  and (_15817_, _15816_, _02524_);
  or (_15818_, _15817_, _02974_);
  or (_15819_, _15818_, _15814_);
  and (_15820_, _05633_, _04670_);
  or (_15821_, _15820_, _15772_);
  or (_15822_, _15821_, _05261_);
  and (_15824_, _15822_, _15819_);
  or (_15825_, _15824_, _02977_);
  and (_15826_, _11525_, _04670_);
  or (_15827_, _15772_, _07092_);
  or (_15828_, _15827_, _15826_);
  and (_15829_, _15828_, _07104_);
  and (_15830_, _15829_, _15825_);
  or (_15831_, _15830_, _15775_);
  and (_15832_, _15831_, _03095_);
  or (_15833_, _15772_, _04890_);
  and (_15835_, _15784_, _03094_);
  and (_15836_, _15821_, _02991_);
  or (_15837_, _15836_, _15835_);
  and (_15838_, _15837_, _15833_);
  or (_15839_, _15838_, _02994_);
  or (_15840_, _15839_, _15832_);
  nor (_15841_, _11524_, _08190_);
  or (_15842_, _15772_, _07120_);
  or (_15843_, _15842_, _15841_);
  and (_15844_, _15843_, _07118_);
  and (_15846_, _15844_, _15840_);
  nor (_15847_, _11530_, _08190_);
  or (_15848_, _15847_, _15772_);
  and (_15849_, _15848_, _03099_);
  or (_15850_, _15849_, _03133_);
  or (_15851_, _15850_, _15846_);
  or (_15852_, _15781_, _03138_);
  and (_15853_, _15852_, _02853_);
  and (_15854_, _15853_, _15851_);
  and (_15855_, _11580_, _04670_);
  or (_15857_, _15855_, _15772_);
  and (_15858_, _15857_, _02852_);
  or (_15859_, _15858_, _34450_);
  or (_15860_, _15859_, _15854_);
  and (_35617_[5], _15860_, _15771_);
  or (_15861_, _34446_, \oc8051_golden_model_1.DPL [6]);
  and (_15862_, _15861_, _35583_);
  not (_15863_, \oc8051_golden_model_1.DPL [6]);
  nor (_15864_, _04670_, _15863_);
  and (_15865_, _11601_, _04670_);
  or (_15867_, _15865_, _15864_);
  and (_15868_, _15867_, _03107_);
  nor (_15869_, _04735_, _08190_);
  or (_15870_, _15869_, _15864_);
  or (_15871_, _15870_, _03860_);
  nor (_15872_, _11610_, _08190_);
  or (_15873_, _15872_, _15864_);
  or (_15874_, _15873_, _06162_);
  and (_15875_, _04670_, \oc8051_golden_model_1.ACC [6]);
  or (_15876_, _15875_, _15864_);
  and (_15878_, _15876_, _02837_);
  nor (_15879_, _02837_, _15863_);
  or (_15880_, _15879_, _02932_);
  or (_15881_, _15880_, _15878_);
  and (_15882_, _15881_, _03693_);
  and (_15883_, _15882_, _15874_);
  and (_15884_, _15870_, _02930_);
  or (_15885_, _15884_, _02928_);
  or (_15886_, _15885_, _15883_);
  or (_15887_, _15876_, _02943_);
  and (_15889_, _15887_, _08210_);
  and (_15890_, _15889_, _15886_);
  nor (_15891_, _08218_, \oc8051_golden_model_1.DPL [6]);
  nor (_15892_, _15891_, _08219_);
  and (_15893_, _15892_, _08209_);
  or (_15894_, _15893_, _15890_);
  and (_15895_, _15894_, _08194_);
  nor (_15896_, _05549_, _08194_);
  or (_15897_, _15896_, _03861_);
  or (_15898_, _15897_, _15895_);
  and (_15900_, _15898_, _15871_);
  or (_15901_, _15900_, _03850_);
  and (_15902_, _05798_, _04670_);
  or (_15903_, _15864_, _06726_);
  or (_15904_, _15903_, _15902_);
  and (_15905_, _15904_, _02970_);
  and (_15906_, _15905_, _15901_);
  nor (_15907_, _11711_, _08190_);
  or (_15908_, _15907_, _15864_);
  and (_15909_, _15908_, _02524_);
  or (_15911_, _15909_, _02974_);
  or (_15912_, _15911_, _15906_);
  and (_15913_, _11718_, _04670_);
  or (_15914_, _15913_, _15864_);
  or (_15915_, _15914_, _05261_);
  and (_15916_, _15915_, _15912_);
  or (_15917_, _15916_, _02977_);
  and (_15918_, _11728_, _04670_);
  or (_15919_, _15864_, _07092_);
  or (_15920_, _15919_, _15918_);
  and (_15922_, _15920_, _07104_);
  and (_15923_, _15922_, _15917_);
  or (_15924_, _15923_, _15868_);
  and (_15925_, _15924_, _03095_);
  or (_15926_, _15864_, _04784_);
  and (_15927_, _15876_, _03094_);
  and (_15928_, _15914_, _02991_);
  or (_15929_, _15928_, _15927_);
  and (_15930_, _15929_, _15926_);
  or (_15931_, _15930_, _02994_);
  or (_15933_, _15931_, _15925_);
  nor (_15934_, _11726_, _08190_);
  or (_15935_, _15864_, _07120_);
  or (_15936_, _15935_, _15934_);
  and (_15937_, _15936_, _07118_);
  and (_15938_, _15937_, _15933_);
  nor (_15939_, _11600_, _08190_);
  or (_15940_, _15939_, _15864_);
  and (_15941_, _15940_, _03099_);
  or (_15942_, _15941_, _03133_);
  or (_15944_, _15942_, _15938_);
  or (_15945_, _15873_, _03138_);
  and (_15946_, _15945_, _02853_);
  and (_15947_, _15946_, _15944_);
  and (_15948_, _11778_, _04670_);
  or (_15949_, _15948_, _15864_);
  and (_15950_, _15949_, _02852_);
  or (_15951_, _15950_, _34450_);
  or (_15952_, _15951_, _15947_);
  and (_35617_[6], _15952_, _15862_);
  nor (_15954_, _34446_, _09337_);
  nor (_15955_, _08221_, \oc8051_golden_model_1.DPH [0]);
  nor (_15956_, _15955_, _08306_);
  and (_15957_, _15956_, _08209_);
  nor (_15958_, _05183_, _09337_);
  nor (_15959_, _05036_, _08285_);
  or (_15960_, _15959_, _15958_);
  or (_15961_, _15960_, _06162_);
  and (_15962_, _05183_, \oc8051_golden_model_1.ACC [0]);
  or (_15963_, _15962_, _15958_);
  and (_15965_, _15963_, _02837_);
  nor (_15966_, _02837_, _09337_);
  or (_15967_, _15966_, _02932_);
  or (_15968_, _15967_, _15965_);
  and (_15969_, _15968_, _03693_);
  and (_15970_, _15969_, _15961_);
  and (_15971_, _04616_, _03805_);
  or (_15972_, _15971_, _15958_);
  and (_15973_, _15972_, _02930_);
  or (_15974_, _15973_, _02928_);
  or (_15976_, _15974_, _15970_);
  or (_15977_, _15963_, _02943_);
  and (_15978_, _15977_, _08210_);
  and (_15979_, _15978_, _15976_);
  or (_15980_, _15979_, _15957_);
  and (_15981_, _15980_, _08194_);
  nor (_15982_, _08194_, _02835_);
  or (_15983_, _15982_, _03861_);
  or (_15984_, _15983_, _15981_);
  or (_15985_, _15972_, _03860_);
  and (_15987_, _15985_, _15984_);
  or (_15988_, _15987_, _03850_);
  and (_15989_, _06114_, _05183_);
  or (_15990_, _15958_, _06726_);
  or (_15991_, _15990_, _15989_);
  and (_15992_, _15991_, _15988_);
  or (_15993_, _15992_, _02524_);
  nor (_15994_, _10530_, _08285_);
  or (_15995_, _15958_, _02970_);
  or (_15996_, _15995_, _15994_);
  and (_15998_, _15996_, _05261_);
  and (_15999_, _15998_, _15993_);
  and (_16000_, _05183_, _05647_);
  or (_16001_, _16000_, _15958_);
  and (_16002_, _16001_, _02974_);
  or (_16003_, _16002_, _02977_);
  or (_16004_, _16003_, _15999_);
  and (_16005_, _10427_, _05183_);
  or (_16006_, _16005_, _15958_);
  or (_16007_, _16006_, _07092_);
  and (_16009_, _16007_, _16004_);
  or (_16010_, _16009_, _03107_);
  and (_16011_, _10546_, _04616_);
  or (_16012_, _15958_, _07104_);
  or (_16013_, _16012_, _16011_);
  and (_16014_, _16013_, _03881_);
  and (_16015_, _16014_, _16010_);
  nand (_16016_, _16001_, _02991_);
  nor (_16017_, _16016_, _15959_);
  or (_16018_, _16017_, _16015_);
  and (_16020_, _16018_, _06161_);
  or (_16021_, _15958_, _05036_);
  and (_16022_, _15963_, _03094_);
  and (_16023_, _16022_, _16021_);
  or (_16024_, _16023_, _02994_);
  or (_16025_, _16024_, _16020_);
  nor (_16026_, _10425_, _08285_);
  or (_16027_, _15958_, _07120_);
  or (_16028_, _16027_, _16026_);
  and (_16029_, _16028_, _07118_);
  and (_16031_, _16029_, _16025_);
  nor (_16032_, _10423_, _08285_);
  or (_16033_, _16032_, _15958_);
  and (_16034_, _16033_, _03099_);
  or (_16035_, _16034_, _15390_);
  or (_16036_, _16035_, _16031_);
  or (_16037_, _15960_, _03330_);
  and (_16038_, _16037_, _34446_);
  and (_16039_, _16038_, _16036_);
  or (_16040_, _16039_, _15954_);
  and (_35616_[0], _16040_, _35583_);
  not (_16042_, \oc8051_golden_model_1.DPH [1]);
  nor (_16043_, _34446_, _16042_);
  nor (_16044_, _05183_, _16042_);
  or (_16045_, _16044_, _04988_);
  or (_16046_, _05183_, \oc8051_golden_model_1.DPH [1]);
  nand (_16047_, _04616_, _02477_);
  and (_16048_, _16047_, _16046_);
  and (_16049_, _16048_, _03094_);
  and (_16050_, _16049_, _16045_);
  and (_16052_, _16046_, _02974_);
  nand (_16053_, _04616_, _03660_);
  and (_16054_, _16053_, _16052_);
  nor (_16055_, _08306_, \oc8051_golden_model_1.DPH [1]);
  nor (_16056_, _16055_, _08307_);
  and (_16057_, _16056_, _08209_);
  nand (_16058_, _10622_, _04616_);
  and (_16059_, _16058_, _16046_);
  or (_16060_, _16059_, _06162_);
  and (_16061_, _16048_, _02837_);
  nor (_16063_, _02837_, _16042_);
  or (_16064_, _16063_, _02932_);
  or (_16065_, _16064_, _16061_);
  and (_16066_, _16065_, _03693_);
  and (_16067_, _16066_, _16060_);
  nor (_16068_, _08285_, _03989_);
  or (_16069_, _16068_, _16044_);
  and (_16070_, _16069_, _02930_);
  or (_16071_, _16070_, _02928_);
  or (_16072_, _16071_, _16067_);
  or (_16074_, _16048_, _02943_);
  and (_16075_, _16074_, _08210_);
  and (_16076_, _16075_, _16072_);
  or (_16077_, _16076_, _16057_);
  and (_16078_, _16077_, _08194_);
  nor (_16079_, _03742_, _08194_);
  or (_16080_, _16079_, _03861_);
  or (_16081_, _16080_, _16078_);
  or (_16082_, _16069_, _03860_);
  and (_16083_, _16082_, _16081_);
  or (_16085_, _16083_, _03850_);
  and (_16086_, _06113_, _05183_);
  or (_16087_, _16044_, _06726_);
  or (_16088_, _16087_, _16086_);
  and (_16089_, _16088_, _02970_);
  and (_16090_, _16089_, _16085_);
  and (_16091_, _16046_, _02524_);
  nand (_16092_, _10719_, _04616_);
  and (_16093_, _16092_, _16091_);
  or (_16094_, _16093_, _16090_);
  and (_16096_, _16094_, _05261_);
  or (_16097_, _16096_, _16054_);
  and (_16098_, _16097_, _03882_);
  or (_16099_, _10613_, _08285_);
  and (_16100_, _16046_, _02991_);
  and (_16101_, _16100_, _16099_);
  or (_16102_, _10610_, _08285_);
  and (_16103_, _16046_, _03107_);
  and (_16104_, _16103_, _16102_);
  or (_16105_, _10614_, _08285_);
  and (_16107_, _16046_, _02977_);
  and (_16108_, _16107_, _16105_);
  or (_16109_, _16108_, _16104_);
  or (_16110_, _16109_, _16101_);
  or (_16111_, _16110_, _16098_);
  and (_16112_, _16111_, _06161_);
  or (_16113_, _16112_, _16050_);
  and (_16114_, _16113_, _03100_);
  or (_16115_, _16047_, _04988_);
  and (_16116_, _16046_, _03099_);
  and (_16118_, _16116_, _16115_);
  or (_16119_, _16118_, _03133_);
  or (_16120_, _16053_, _04988_);
  and (_16121_, _16046_, _02994_);
  and (_16122_, _16121_, _16120_);
  or (_16123_, _16122_, _16119_);
  or (_16124_, _16123_, _16114_);
  or (_16125_, _16059_, _03138_);
  and (_16126_, _16125_, _16124_);
  or (_16127_, _16126_, _02852_);
  nor (_16129_, _16044_, _02853_);
  nand (_16130_, _16129_, _16058_);
  and (_16131_, _16130_, _34446_);
  and (_16132_, _16131_, _16127_);
  or (_16133_, _16132_, _16043_);
  and (_35616_[1], _16133_, _35583_);
  or (_16134_, _34446_, \oc8051_golden_model_1.DPH [2]);
  and (_16135_, _16134_, _35583_);
  not (_16136_, \oc8051_golden_model_1.DPH [2]);
  nor (_16137_, _05183_, _16136_);
  and (_16139_, _10942_, _04616_);
  or (_16140_, _16139_, _16137_);
  and (_16141_, _16140_, _03107_);
  nor (_16142_, _08285_, _04413_);
  or (_16143_, _16142_, _16137_);
  or (_16144_, _16143_, _03860_);
  nor (_16145_, _10824_, _08285_);
  or (_16146_, _16145_, _16137_);
  or (_16147_, _16146_, _06162_);
  and (_16148_, _05183_, \oc8051_golden_model_1.ACC [2]);
  or (_16150_, _16148_, _16137_);
  and (_16151_, _16150_, _02837_);
  nor (_16152_, _02837_, _16136_);
  or (_16153_, _16152_, _02932_);
  or (_16154_, _16153_, _16151_);
  and (_16155_, _16154_, _03693_);
  and (_16156_, _16155_, _16147_);
  and (_16157_, _16143_, _02930_);
  or (_16158_, _16157_, _02928_);
  or (_16159_, _16158_, _16156_);
  or (_16161_, _16150_, _02943_);
  and (_16162_, _16161_, _08210_);
  and (_16163_, _16162_, _16159_);
  or (_16164_, _08307_, \oc8051_golden_model_1.DPH [2]);
  nor (_16165_, _08308_, _08210_);
  and (_16166_, _16165_, _16164_);
  or (_16167_, _16166_, _16163_);
  and (_16168_, _16167_, _08194_);
  nor (_16169_, _03320_, _08194_);
  or (_16170_, _16169_, _03861_);
  or (_16172_, _16170_, _16168_);
  and (_16173_, _16172_, _16144_);
  or (_16174_, _16173_, _03850_);
  or (_16175_, _16137_, _06726_);
  and (_16176_, _06117_, _05183_);
  or (_16177_, _16176_, _16175_);
  and (_16178_, _16177_, _02970_);
  and (_16179_, _16178_, _16174_);
  not (_16180_, _05183_);
  nor (_16181_, _10922_, _16180_);
  or (_16183_, _16181_, _16137_);
  and (_16184_, _16183_, _02524_);
  or (_16185_, _16184_, _02974_);
  or (_16186_, _16185_, _16179_);
  and (_16187_, _05183_, _05690_);
  or (_16188_, _16187_, _16137_);
  or (_16189_, _16188_, _05261_);
  and (_16190_, _16189_, _16186_);
  or (_16191_, _16190_, _02977_);
  and (_16192_, _10936_, _04616_);
  or (_16194_, _16137_, _07092_);
  or (_16195_, _16194_, _16192_);
  and (_16196_, _16195_, _07104_);
  and (_16197_, _16196_, _16191_);
  or (_16198_, _16197_, _16141_);
  and (_16199_, _16198_, _03095_);
  or (_16200_, _16137_, _05086_);
  and (_16201_, _16150_, _03094_);
  and (_16202_, _16188_, _02991_);
  or (_16203_, _16202_, _16201_);
  and (_16205_, _16203_, _16200_);
  or (_16206_, _16205_, _02994_);
  or (_16207_, _16206_, _16199_);
  nor (_16208_, _10935_, _08285_);
  or (_16209_, _16137_, _07120_);
  or (_16210_, _16209_, _16208_);
  and (_16211_, _16210_, _07118_);
  and (_16212_, _16211_, _16207_);
  nor (_16213_, _10941_, _08285_);
  or (_16214_, _16213_, _16137_);
  and (_16216_, _16214_, _03099_);
  or (_16217_, _16216_, _03133_);
  or (_16218_, _16217_, _16212_);
  or (_16219_, _16146_, _03138_);
  and (_16220_, _16219_, _02853_);
  and (_16221_, _16220_, _16218_);
  and (_16222_, _10988_, _04616_);
  or (_16223_, _16222_, _16137_);
  and (_16224_, _16223_, _02852_);
  or (_16225_, _16224_, _34450_);
  or (_16227_, _16225_, _16221_);
  and (_35616_[2], _16227_, _16135_);
  or (_16228_, _34446_, \oc8051_golden_model_1.DPH [3]);
  and (_16229_, _16228_, _35583_);
  not (_16230_, \oc8051_golden_model_1.DPH [3]);
  nor (_16231_, _05183_, _16230_);
  and (_16232_, _11134_, _04616_);
  or (_16233_, _16232_, _16231_);
  and (_16234_, _16233_, _03107_);
  nor (_16235_, _08285_, _04226_);
  or (_16237_, _16235_, _16231_);
  or (_16238_, _16237_, _03860_);
  or (_16239_, _08308_, \oc8051_golden_model_1.DPH [3]);
  nand (_16240_, _16239_, _08209_);
  nor (_16241_, _16240_, _08309_);
  nor (_16242_, _11014_, _08285_);
  or (_16243_, _16242_, _16231_);
  or (_16244_, _16243_, _06162_);
  and (_16245_, _05183_, \oc8051_golden_model_1.ACC [3]);
  or (_16246_, _16245_, _16231_);
  and (_16248_, _16246_, _02837_);
  nor (_16249_, _02837_, _16230_);
  or (_16250_, _16249_, _02932_);
  or (_16251_, _16250_, _16248_);
  and (_16252_, _16251_, _03693_);
  and (_16253_, _16252_, _16244_);
  and (_16254_, _16237_, _02930_);
  or (_16255_, _16254_, _02928_);
  or (_16256_, _16255_, _16253_);
  or (_16257_, _16246_, _02943_);
  and (_16259_, _16257_, _08210_);
  and (_16260_, _16259_, _16256_);
  or (_16261_, _16260_, _16241_);
  and (_16262_, _16261_, _08194_);
  and (_16263_, _02975_, _02774_);
  or (_16264_, _16263_, _03861_);
  or (_16265_, _16264_, _16262_);
  and (_16266_, _16265_, _16238_);
  or (_16267_, _16266_, _03850_);
  or (_16268_, _16231_, _06726_);
  and (_16270_, _06116_, _05183_);
  or (_16271_, _16270_, _16268_);
  and (_16272_, _16271_, _02970_);
  and (_16273_, _16272_, _16267_);
  nor (_16274_, _11114_, _16180_);
  or (_16275_, _16274_, _16231_);
  and (_16276_, _16275_, _02524_);
  or (_16277_, _16276_, _02974_);
  or (_16278_, _16277_, _16273_);
  and (_16279_, _05183_, _05616_);
  or (_16281_, _16279_, _16231_);
  or (_16282_, _16281_, _05261_);
  and (_16283_, _16282_, _16278_);
  or (_16284_, _16283_, _02977_);
  and (_16285_, _11128_, _04616_);
  or (_16286_, _16231_, _07092_);
  or (_16287_, _16286_, _16285_);
  and (_16288_, _16287_, _07104_);
  and (_16289_, _16288_, _16284_);
  or (_16290_, _16289_, _16234_);
  and (_16292_, _16290_, _03095_);
  or (_16293_, _16231_, _04939_);
  and (_16294_, _16246_, _03094_);
  and (_16295_, _16281_, _02991_);
  or (_16296_, _16295_, _16294_);
  and (_16297_, _16296_, _16293_);
  or (_16298_, _16297_, _02994_);
  or (_16299_, _16298_, _16292_);
  nor (_16300_, _11127_, _08285_);
  or (_16301_, _16231_, _07120_);
  or (_16303_, _16301_, _16300_);
  and (_16304_, _16303_, _07118_);
  and (_16305_, _16304_, _16299_);
  nor (_16306_, _11133_, _08285_);
  or (_16307_, _16306_, _16231_);
  and (_16308_, _16307_, _03099_);
  or (_16309_, _16308_, _03133_);
  or (_16310_, _16309_, _16305_);
  or (_16311_, _16243_, _03138_);
  and (_16312_, _16311_, _02853_);
  and (_16314_, _16312_, _16310_);
  and (_16315_, _11185_, _04616_);
  or (_16316_, _16315_, _16231_);
  and (_16317_, _16316_, _02852_);
  or (_16318_, _16317_, _34450_);
  or (_16319_, _16318_, _16314_);
  and (_35616_[3], _16319_, _16229_);
  or (_16320_, _34446_, \oc8051_golden_model_1.DPH [4]);
  and (_16321_, _16320_, _35583_);
  not (_16322_, \oc8051_golden_model_1.DPH [4]);
  nor (_16324_, _05183_, _16322_);
  and (_16325_, _11333_, _04616_);
  or (_16326_, _16325_, _16324_);
  and (_16327_, _16326_, _03107_);
  nor (_16328_, _05143_, _08285_);
  or (_16329_, _16328_, _16324_);
  or (_16330_, _16329_, _03860_);
  nor (_16331_, _11207_, _08285_);
  or (_16332_, _16331_, _16324_);
  or (_16333_, _16332_, _06162_);
  and (_16335_, _05183_, \oc8051_golden_model_1.ACC [4]);
  or (_16336_, _16335_, _16324_);
  and (_16337_, _16336_, _02837_);
  nor (_16338_, _02837_, _16322_);
  or (_16339_, _16338_, _02932_);
  or (_16340_, _16339_, _16337_);
  and (_16341_, _16340_, _03693_);
  and (_16342_, _16341_, _16333_);
  and (_16343_, _16329_, _02930_);
  or (_16344_, _16343_, _02928_);
  or (_16346_, _16344_, _16342_);
  or (_16347_, _16336_, _02943_);
  and (_16348_, _16347_, _08210_);
  and (_16349_, _16348_, _16346_);
  or (_16350_, _08309_, \oc8051_golden_model_1.DPH [4]);
  nor (_16351_, _08310_, _08210_);
  and (_16352_, _16351_, _16350_);
  or (_16353_, _16352_, _16349_);
  and (_16354_, _16353_, _08194_);
  nor (_16355_, _03620_, _08194_);
  or (_16357_, _16355_, _03861_);
  or (_16358_, _16357_, _16354_);
  and (_16359_, _16358_, _16330_);
  or (_16360_, _16359_, _03850_);
  or (_16361_, _16324_, _06726_);
  and (_16362_, _06121_, _05183_);
  or (_16363_, _16362_, _16361_);
  and (_16364_, _16363_, _02970_);
  and (_16365_, _16364_, _16360_);
  nor (_16366_, _11313_, _16180_);
  or (_16368_, _16366_, _16324_);
  and (_16369_, _16368_, _02524_);
  or (_16370_, _16369_, _02974_);
  or (_16371_, _16370_, _16365_);
  and (_16372_, _05629_, _05183_);
  or (_16373_, _16372_, _16324_);
  or (_16374_, _16373_, _05261_);
  and (_16375_, _16374_, _16371_);
  or (_16376_, _16375_, _02977_);
  and (_16377_, _11327_, _04616_);
  or (_16378_, _16324_, _07092_);
  or (_16379_, _16378_, _16377_);
  and (_16380_, _16379_, _07104_);
  and (_16381_, _16380_, _16376_);
  or (_16382_, _16381_, _16327_);
  and (_16383_, _16382_, _03095_);
  or (_16384_, _16324_, _05190_);
  and (_16385_, _16336_, _03094_);
  and (_16386_, _16373_, _02991_);
  or (_16387_, _16386_, _16385_);
  and (_16390_, _16387_, _16384_);
  or (_16391_, _16390_, _02994_);
  or (_16392_, _16391_, _16383_);
  nor (_16393_, _11326_, _08285_);
  or (_16394_, _16324_, _07120_);
  or (_16395_, _16394_, _16393_);
  and (_16396_, _16395_, _07118_);
  and (_16397_, _16396_, _16392_);
  nor (_16398_, _11332_, _08285_);
  or (_16399_, _16398_, _16324_);
  and (_16401_, _16399_, _03099_);
  or (_16402_, _16401_, _03133_);
  or (_16403_, _16402_, _16397_);
  or (_16404_, _16332_, _03138_);
  and (_16405_, _16404_, _02853_);
  and (_16406_, _16405_, _16403_);
  and (_16407_, _11383_, _04616_);
  or (_16408_, _16407_, _16324_);
  and (_16409_, _16408_, _02852_);
  or (_16410_, _16409_, _34450_);
  or (_16412_, _16410_, _16406_);
  and (_35616_[4], _16412_, _16321_);
  or (_16413_, _34446_, \oc8051_golden_model_1.DPH [5]);
  and (_16414_, _16413_, _35583_);
  and (_16415_, _16180_, \oc8051_golden_model_1.DPH [5]);
  and (_16416_, _11531_, _04616_);
  or (_16417_, _16416_, _16415_);
  and (_16418_, _16417_, _03107_);
  nor (_16419_, _04839_, _08285_);
  or (_16420_, _16419_, _16415_);
  or (_16422_, _16420_, _03860_);
  nor (_16423_, _11408_, _08285_);
  or (_16424_, _16423_, _16415_);
  or (_16425_, _16424_, _06162_);
  and (_16426_, _05183_, \oc8051_golden_model_1.ACC [5]);
  or (_16427_, _16426_, _16415_);
  and (_16428_, _16427_, _02837_);
  and (_16429_, _09167_, \oc8051_golden_model_1.DPH [5]);
  or (_16430_, _16429_, _02932_);
  or (_16431_, _16430_, _16428_);
  and (_16433_, _16431_, _03693_);
  and (_16434_, _16433_, _16425_);
  and (_16435_, _16420_, _02930_);
  or (_16436_, _16435_, _02928_);
  or (_16437_, _16436_, _16434_);
  or (_16438_, _16427_, _02943_);
  and (_16439_, _16438_, _08210_);
  and (_16440_, _16439_, _16437_);
  or (_16441_, _08310_, \oc8051_golden_model_1.DPH [5]);
  nor (_16442_, _08311_, _08210_);
  and (_16444_, _16442_, _16441_);
  or (_16445_, _16444_, _16440_);
  and (_16446_, _16445_, _08194_);
  nor (_16447_, _03179_, _08194_);
  or (_16448_, _16447_, _03861_);
  or (_16449_, _16448_, _16446_);
  and (_16450_, _16449_, _16422_);
  or (_16451_, _16450_, _03850_);
  or (_16452_, _16415_, _06726_);
  and (_16453_, _06120_, _05183_);
  or (_16455_, _16453_, _16452_);
  and (_16456_, _16455_, _02970_);
  and (_16457_, _16456_, _16451_);
  nor (_16458_, _11511_, _16180_);
  or (_16459_, _16458_, _16415_);
  and (_16460_, _16459_, _02524_);
  or (_16461_, _16460_, _02974_);
  or (_16462_, _16461_, _16457_);
  and (_16463_, _05633_, _05183_);
  or (_16464_, _16463_, _16415_);
  or (_16466_, _16464_, _05261_);
  and (_16467_, _16466_, _16462_);
  or (_16468_, _16467_, _02977_);
  and (_16469_, _11525_, _04616_);
  or (_16470_, _16415_, _07092_);
  or (_16471_, _16470_, _16469_);
  and (_16472_, _16471_, _07104_);
  and (_16473_, _16472_, _16468_);
  or (_16474_, _16473_, _16418_);
  and (_16475_, _16474_, _03095_);
  or (_16477_, _16415_, _04890_);
  and (_16478_, _16427_, _03094_);
  and (_16479_, _16464_, _02991_);
  or (_16480_, _16479_, _16478_);
  and (_16481_, _16480_, _16477_);
  or (_16482_, _16481_, _02994_);
  or (_16483_, _16482_, _16475_);
  nor (_16484_, _11524_, _08285_);
  or (_16485_, _16415_, _07120_);
  or (_16486_, _16485_, _16484_);
  and (_16488_, _16486_, _07118_);
  and (_16489_, _16488_, _16483_);
  nor (_16490_, _11530_, _08285_);
  or (_16491_, _16490_, _16415_);
  and (_16492_, _16491_, _03099_);
  or (_16493_, _16492_, _03133_);
  or (_16494_, _16493_, _16489_);
  or (_16495_, _16424_, _03138_);
  and (_16496_, _16495_, _02853_);
  and (_16497_, _16496_, _16494_);
  and (_16499_, _11580_, _04616_);
  or (_16500_, _16499_, _16415_);
  and (_16501_, _16500_, _02852_);
  or (_16502_, _16501_, _34450_);
  or (_16503_, _16502_, _16497_);
  and (_35616_[5], _16503_, _16414_);
  or (_16504_, _34446_, \oc8051_golden_model_1.DPH [6]);
  and (_16505_, _16504_, _35583_);
  not (_16506_, \oc8051_golden_model_1.DPH [6]);
  nor (_16507_, _05183_, _16506_);
  and (_16509_, _11601_, _04616_);
  or (_16510_, _16509_, _16507_);
  and (_16511_, _16510_, _03107_);
  nor (_16512_, _04735_, _08285_);
  or (_16513_, _16512_, _16507_);
  or (_16514_, _16513_, _03860_);
  nor (_16515_, _11610_, _08285_);
  or (_16516_, _16515_, _16507_);
  or (_16517_, _16516_, _06162_);
  and (_16518_, _05183_, \oc8051_golden_model_1.ACC [6]);
  or (_16520_, _16518_, _16507_);
  and (_16521_, _16520_, _02837_);
  nor (_16522_, _02837_, _16506_);
  or (_16523_, _16522_, _02932_);
  or (_16524_, _16523_, _16521_);
  and (_16525_, _16524_, _03693_);
  and (_16526_, _16525_, _16517_);
  and (_16527_, _16513_, _02930_);
  or (_16528_, _16527_, _02928_);
  or (_16529_, _16528_, _16526_);
  or (_16531_, _16520_, _02943_);
  and (_16532_, _16531_, _08210_);
  and (_16533_, _16532_, _16529_);
  or (_16534_, _08311_, \oc8051_golden_model_1.DPH [6]);
  nor (_16535_, _08312_, _08210_);
  and (_16536_, _16535_, _16534_);
  or (_16537_, _16536_, _16533_);
  and (_16538_, _16537_, _08194_);
  nor (_16539_, _08194_, _02889_);
  or (_16540_, _16539_, _03861_);
  or (_16542_, _16540_, _16538_);
  and (_16543_, _16542_, _16514_);
  or (_16544_, _16543_, _03850_);
  or (_16545_, _16507_, _06726_);
  and (_16546_, _05798_, _05183_);
  or (_16547_, _16546_, _16545_);
  and (_16548_, _16547_, _02970_);
  and (_16549_, _16548_, _16544_);
  nor (_16550_, _11711_, _16180_);
  or (_16551_, _16550_, _16507_);
  and (_16553_, _16551_, _02524_);
  or (_16554_, _16553_, _02974_);
  or (_16555_, _16554_, _16549_);
  and (_16556_, _11718_, _05183_);
  or (_16557_, _16556_, _16507_);
  or (_16558_, _16557_, _05261_);
  and (_16559_, _16558_, _16555_);
  or (_16560_, _16559_, _02977_);
  and (_16561_, _11728_, _04616_);
  or (_16562_, _16507_, _07092_);
  or (_16564_, _16562_, _16561_);
  and (_16565_, _16564_, _07104_);
  and (_16566_, _16565_, _16560_);
  or (_16567_, _16566_, _16511_);
  and (_16568_, _16567_, _03095_);
  or (_16569_, _16507_, _04784_);
  and (_16570_, _16520_, _03094_);
  and (_16571_, _16557_, _02991_);
  or (_16572_, _16571_, _16570_);
  and (_16573_, _16572_, _16569_);
  or (_16575_, _16573_, _02994_);
  or (_16576_, _16575_, _16568_);
  nor (_16577_, _11726_, _08285_);
  or (_16578_, _16507_, _07120_);
  or (_16579_, _16578_, _16577_);
  and (_16580_, _16579_, _07118_);
  and (_16581_, _16580_, _16576_);
  nor (_16582_, _11600_, _08285_);
  or (_16583_, _16582_, _16507_);
  and (_16584_, _16583_, _03099_);
  or (_16586_, _16584_, _03133_);
  or (_16587_, _16586_, _16581_);
  or (_16588_, _16516_, _03138_);
  and (_16589_, _16588_, _02853_);
  and (_16590_, _16589_, _16587_);
  and (_16591_, _11778_, _04616_);
  or (_16592_, _16591_, _16507_);
  and (_16593_, _16592_, _02852_);
  or (_16594_, _16593_, _34450_);
  or (_16595_, _16594_, _16590_);
  and (_35616_[6], _16595_, _16505_);
  and (_35618_[0], \oc8051_golden_model_1.IE [0], _35583_);
  and (_35618_[1], \oc8051_golden_model_1.IE [1], _35583_);
  and (_35618_[2], \oc8051_golden_model_1.IE [2], _35583_);
  and (_35618_[3], \oc8051_golden_model_1.IE [3], _35583_);
  and (_35618_[4], \oc8051_golden_model_1.IE [4], _35583_);
  and (_35618_[5], \oc8051_golden_model_1.IE [5], _35583_);
  and (_35618_[6], \oc8051_golden_model_1.IE [6], _35583_);
  and (_35619_[0], \oc8051_golden_model_1.IP [0], _35583_);
  and (_35619_[1], \oc8051_golden_model_1.IP [1], _35583_);
  and (_35619_[2], \oc8051_golden_model_1.IP [2], _35583_);
  and (_35619_[3], \oc8051_golden_model_1.IP [3], _35583_);
  and (_35619_[4], \oc8051_golden_model_1.IP [4], _35583_);
  and (_35619_[5], \oc8051_golden_model_1.IP [5], _35583_);
  and (_35619_[6], \oc8051_golden_model_1.IP [6], _35583_);
  not (_16598_, \oc8051_golden_model_1.P0 [0]);
  nor (_16599_, _34446_, _16598_);
  or (_16600_, _16599_, rst);
  nor (_16601_, _04673_, _16598_);
  and (_16602_, _10546_, _04673_);
  or (_16604_, _16602_, _16601_);
  and (_16605_, _16604_, _03107_);
  and (_16606_, _04673_, _03805_);
  or (_16607_, _16606_, _16601_);
  or (_16608_, _16607_, _03860_);
  nor (_16609_, _05036_, _08395_);
  or (_16610_, _16609_, _16601_);
  or (_16611_, _16610_, _06162_);
  and (_16612_, _04673_, \oc8051_golden_model_1.ACC [0]);
  or (_16613_, _16612_, _16601_);
  and (_16615_, _16613_, _02837_);
  nor (_16616_, _02837_, _16598_);
  or (_16617_, _16616_, _02932_);
  or (_16618_, _16617_, _16615_);
  and (_16619_, _16618_, _02939_);
  and (_16620_, _16619_, _16611_);
  and (_16621_, _16607_, _02930_);
  or (_16622_, _16621_, _16620_);
  nor (_16623_, _04613_, _16598_);
  and (_16624_, _10441_, _04613_);
  or (_16626_, _16624_, _16623_);
  and (_16627_, _16626_, _02799_);
  or (_16628_, _16627_, _02928_);
  or (_16629_, _16628_, _16622_);
  or (_16630_, _16613_, _02943_);
  and (_16631_, _16630_, _16629_);
  or (_16632_, _16631_, _02796_);
  or (_16633_, _16601_, _02927_);
  and (_16634_, _16633_, _06189_);
  and (_16635_, _16634_, _16632_);
  and (_16637_, _16610_, _02790_);
  or (_16638_, _16637_, _16635_);
  and (_16639_, _16638_, _02966_);
  or (_16640_, _10472_, _10429_);
  and (_16641_, _16640_, _04613_);
  or (_16642_, _16641_, _16623_);
  and (_16643_, _16642_, _02785_);
  or (_16644_, _16643_, _03861_);
  or (_16645_, _16644_, _16639_);
  and (_16646_, _16645_, _16608_);
  or (_16648_, _16646_, _03850_);
  and (_16649_, _06114_, _04673_);
  or (_16650_, _16601_, _06726_);
  or (_16651_, _16650_, _16649_);
  and (_16652_, _16651_, _02970_);
  and (_16653_, _16652_, _16648_);
  nor (_16654_, _10530_, _08395_);
  or (_16655_, _16654_, _16601_);
  and (_16656_, _16655_, _02524_);
  or (_16657_, _16656_, _02974_);
  or (_16659_, _16657_, _16653_);
  and (_16660_, _04673_, _05647_);
  or (_16661_, _16660_, _16601_);
  or (_16662_, _16661_, _05261_);
  and (_16663_, _16662_, _16659_);
  or (_16664_, _16663_, _02977_);
  and (_16665_, _10427_, _04673_);
  or (_16666_, _16601_, _07092_);
  or (_16667_, _16666_, _16665_);
  and (_16668_, _16667_, _07104_);
  and (_16670_, _16668_, _16664_);
  or (_16671_, _16670_, _16605_);
  and (_16672_, _16671_, _03095_);
  nand (_16673_, _16661_, _02991_);
  nor (_16674_, _16673_, _16609_);
  or (_16675_, _16601_, _05036_);
  and (_16676_, _16613_, _03094_);
  and (_16677_, _16676_, _16675_);
  or (_16678_, _16677_, _02994_);
  or (_16679_, _16678_, _16674_);
  or (_16681_, _16679_, _16672_);
  nor (_16682_, _10425_, _08395_);
  or (_16683_, _16601_, _07120_);
  or (_16684_, _16683_, _16682_);
  and (_16685_, _16684_, _07118_);
  and (_16686_, _16685_, _16681_);
  nor (_16687_, _10423_, _08395_);
  or (_16688_, _16687_, _16601_);
  and (_16689_, _16688_, _03099_);
  or (_16690_, _16689_, _03133_);
  or (_16692_, _16690_, _16686_);
  or (_16693_, _16610_, _03138_);
  and (_16694_, _16693_, _03142_);
  and (_16695_, _16694_, _16692_);
  and (_16696_, _16601_, _02778_);
  or (_16697_, _16696_, _02852_);
  or (_16698_, _16697_, _16695_);
  or (_16699_, _16610_, _02853_);
  and (_16700_, _16699_, _34446_);
  and (_16701_, _16700_, _16698_);
  or (_35621_[0], _16701_, _16600_);
  not (_16703_, \oc8051_golden_model_1.P0 [1]);
  nor (_16704_, _34446_, _16703_);
  or (_16705_, _16704_, rst);
  nand (_16706_, _04673_, _03660_);
  or (_16707_, _04673_, \oc8051_golden_model_1.P0 [1]);
  and (_16708_, _16707_, _02974_);
  and (_16709_, _16708_, _16706_);
  or (_16710_, _10661_, _10620_);
  and (_16711_, _16710_, _04613_);
  nor (_16713_, _04613_, _16703_);
  or (_16714_, _16713_, _02966_);
  or (_16715_, _16714_, _16711_);
  and (_16716_, _10622_, _04673_);
  not (_16717_, _16716_);
  and (_16718_, _16717_, _16707_);
  or (_16719_, _16718_, _06162_);
  nand (_16720_, _04673_, _02477_);
  and (_16721_, _16720_, _16707_);
  and (_16722_, _16721_, _02837_);
  nor (_16724_, _02837_, _16703_);
  or (_16725_, _16724_, _02932_);
  or (_16726_, _16725_, _16722_);
  and (_16727_, _16726_, _02939_);
  and (_16728_, _16727_, _16719_);
  nor (_16729_, _04673_, _16703_);
  nor (_16730_, _08395_, _03989_);
  or (_16731_, _16730_, _16729_);
  and (_16732_, _16731_, _02930_);
  and (_16733_, _10617_, _04613_);
  or (_16735_, _16733_, _16713_);
  and (_16736_, _16735_, _02799_);
  or (_16737_, _16736_, _16732_);
  or (_16738_, _16737_, _02928_);
  or (_16739_, _16738_, _16728_);
  or (_16740_, _16721_, _02943_);
  and (_16741_, _16740_, _16739_);
  or (_16742_, _16741_, _02796_);
  and (_16743_, _10620_, _04613_);
  or (_16744_, _16743_, _16713_);
  or (_16746_, _16744_, _02927_);
  and (_16747_, _16746_, _06189_);
  and (_16748_, _16747_, _16742_);
  and (_16749_, _16733_, _10616_);
  or (_16750_, _16749_, _16713_);
  and (_16751_, _16750_, _02790_);
  or (_16752_, _16751_, _02785_);
  or (_16753_, _16752_, _16748_);
  and (_16754_, _16753_, _16715_);
  or (_16755_, _16754_, _03861_);
  or (_16757_, _16731_, _03860_);
  and (_16758_, _16757_, _16755_);
  or (_16759_, _16758_, _03850_);
  and (_16760_, _06113_, _04673_);
  or (_16761_, _16729_, _06726_);
  or (_16762_, _16761_, _16760_);
  and (_16763_, _16762_, _02970_);
  and (_16764_, _16763_, _16759_);
  nor (_16765_, _10719_, _08395_);
  or (_16766_, _16765_, _16729_);
  and (_16768_, _16766_, _02524_);
  or (_16769_, _16768_, _16764_);
  and (_16770_, _16769_, _05261_);
  or (_16771_, _16770_, _16709_);
  and (_16772_, _16771_, _03882_);
  or (_16773_, _10613_, _08395_);
  and (_16774_, _16707_, _02991_);
  and (_16775_, _16774_, _16773_);
  or (_16776_, _10610_, _08395_);
  and (_16777_, _16707_, _03107_);
  and (_16779_, _16777_, _16776_);
  or (_16780_, _10614_, _08395_);
  and (_16781_, _16707_, _02977_);
  and (_16782_, _16781_, _16780_);
  or (_16783_, _16782_, _16779_);
  or (_16784_, _16783_, _16775_);
  or (_16785_, _16784_, _16772_);
  and (_16786_, _16785_, _06161_);
  or (_16787_, _16729_, _04988_);
  and (_16788_, _16721_, _03094_);
  and (_16790_, _16788_, _16787_);
  or (_16791_, _16790_, _16786_);
  and (_16792_, _16791_, _03100_);
  or (_16793_, _16706_, _04988_);
  and (_16794_, _16707_, _02994_);
  and (_16795_, _16794_, _16793_);
  or (_16796_, _16720_, _04988_);
  and (_16797_, _16707_, _03099_);
  and (_16798_, _16797_, _16796_);
  or (_16799_, _16798_, _03133_);
  or (_16801_, _16799_, _16795_);
  or (_16802_, _16801_, _16792_);
  or (_16803_, _16718_, _03138_);
  and (_16804_, _16803_, _03142_);
  and (_16805_, _16804_, _16802_);
  and (_16806_, _16744_, _02778_);
  or (_16807_, _16806_, _02852_);
  or (_16808_, _16807_, _16805_);
  or (_16809_, _16729_, _02853_);
  or (_16810_, _16809_, _16716_);
  and (_16812_, _16810_, _34446_);
  and (_16813_, _16812_, _16808_);
  or (_35621_[1], _16813_, _16705_);
  not (_16814_, \oc8051_golden_model_1.P0 [2]);
  nor (_16815_, _34446_, _16814_);
  or (_16816_, _16815_, rst);
  nor (_16817_, _04673_, _16814_);
  and (_16818_, _10942_, _04673_);
  or (_16819_, _16818_, _16817_);
  and (_16820_, _16819_, _03107_);
  nor (_16822_, _08395_, _04413_);
  or (_16823_, _16822_, _16817_);
  or (_16824_, _16823_, _03860_);
  nor (_16825_, _10824_, _08395_);
  or (_16826_, _16825_, _16817_);
  or (_16827_, _16826_, _06162_);
  and (_16828_, _04673_, \oc8051_golden_model_1.ACC [2]);
  or (_16829_, _16828_, _16817_);
  and (_16830_, _16829_, _02837_);
  nor (_16831_, _02837_, _16814_);
  or (_16833_, _16831_, _02932_);
  or (_16834_, _16833_, _16830_);
  and (_16835_, _16834_, _02939_);
  and (_16836_, _16835_, _16827_);
  and (_16837_, _16823_, _02930_);
  nor (_16838_, _04613_, _16814_);
  and (_16839_, _10815_, _04613_);
  or (_16840_, _16839_, _16838_);
  and (_16841_, _16840_, _02799_);
  or (_16842_, _16841_, _16837_);
  or (_16844_, _16842_, _02928_);
  or (_16845_, _16844_, _16836_);
  or (_16846_, _16829_, _02943_);
  and (_16847_, _16846_, _16845_);
  or (_16848_, _16847_, _02796_);
  and (_16849_, _10818_, _04613_);
  or (_16850_, _16849_, _16838_);
  or (_16851_, _16850_, _02927_);
  and (_16852_, _16851_, _06189_);
  and (_16853_, _16852_, _16848_);
  and (_16855_, _16839_, _10814_);
  or (_16856_, _16855_, _16838_);
  and (_16857_, _16856_, _02790_);
  or (_16858_, _16857_, _16853_);
  and (_16859_, _16858_, _02966_);
  or (_16860_, _10865_, _10818_);
  and (_16861_, _16860_, _04613_);
  or (_16862_, _16838_, _16861_);
  and (_16863_, _16862_, _02785_);
  or (_16864_, _16863_, _03861_);
  or (_16866_, _16864_, _16859_);
  and (_16867_, _16866_, _16824_);
  or (_16868_, _16867_, _03850_);
  and (_16869_, _06117_, _04673_);
  or (_16870_, _16817_, _06726_);
  or (_16871_, _16870_, _16869_);
  and (_16872_, _16871_, _02970_);
  and (_16873_, _16872_, _16868_);
  nor (_16874_, _10922_, _08395_);
  or (_16875_, _16874_, _16817_);
  and (_16877_, _16875_, _02524_);
  or (_16878_, _16877_, _02974_);
  or (_16879_, _16878_, _16873_);
  and (_16880_, _04673_, _05690_);
  or (_16881_, _16880_, _16817_);
  or (_16882_, _16881_, _05261_);
  and (_16883_, _16882_, _16879_);
  or (_16884_, _16883_, _02977_);
  and (_16885_, _10936_, _04673_);
  or (_16886_, _16817_, _07092_);
  or (_16888_, _16886_, _16885_);
  and (_16889_, _16888_, _07104_);
  and (_16890_, _16889_, _16884_);
  or (_16891_, _16890_, _16820_);
  and (_16892_, _16891_, _03095_);
  or (_16893_, _16817_, _05086_);
  and (_16894_, _16829_, _03094_);
  and (_16895_, _16881_, _02991_);
  or (_16896_, _16895_, _16894_);
  and (_16897_, _16896_, _16893_);
  or (_16899_, _16897_, _02994_);
  or (_16900_, _16899_, _16892_);
  nor (_16901_, _10935_, _08395_);
  or (_16902_, _16817_, _07120_);
  or (_16903_, _16902_, _16901_);
  and (_16904_, _16903_, _07118_);
  and (_16905_, _16904_, _16900_);
  nor (_16906_, _10941_, _08395_);
  or (_16907_, _16906_, _16817_);
  and (_16908_, _16907_, _03099_);
  or (_16910_, _16908_, _03133_);
  or (_16911_, _16910_, _16905_);
  or (_16912_, _16826_, _03138_);
  and (_16913_, _16912_, _03142_);
  and (_16914_, _16913_, _16911_);
  and (_16915_, _16850_, _02778_);
  or (_16916_, _16915_, _02852_);
  or (_16917_, _16916_, _16914_);
  and (_16918_, _10988_, _04673_);
  or (_16919_, _16817_, _02853_);
  or (_16921_, _16919_, _16918_);
  and (_16922_, _16921_, _34446_);
  and (_16923_, _16922_, _16917_);
  or (_35621_[2], _16923_, _16816_);
  not (_16924_, \oc8051_golden_model_1.P0 [3]);
  nor (_16925_, _34446_, _16924_);
  or (_16926_, _16925_, rst);
  nor (_16927_, _04673_, _16924_);
  and (_16928_, _11134_, _04673_);
  or (_16929_, _16928_, _16927_);
  and (_16931_, _16929_, _03107_);
  nor (_16932_, _08395_, _04226_);
  or (_16933_, _16932_, _16927_);
  or (_16934_, _16933_, _03860_);
  or (_16935_, _11009_, _11056_);
  and (_16936_, _16935_, _04613_);
  nor (_16937_, _04613_, _16924_);
  or (_16938_, _16937_, _02966_);
  or (_16939_, _16938_, _16936_);
  nor (_16940_, _11014_, _08395_);
  or (_16942_, _16940_, _16927_);
  or (_16943_, _16942_, _06162_);
  and (_16944_, _04673_, \oc8051_golden_model_1.ACC [3]);
  or (_16945_, _16944_, _16927_);
  and (_16946_, _16945_, _02837_);
  nor (_16947_, _02837_, _16924_);
  or (_16948_, _16947_, _02932_);
  or (_16949_, _16948_, _16946_);
  and (_16950_, _16949_, _02939_);
  and (_16951_, _16950_, _16943_);
  and (_16953_, _16933_, _02930_);
  and (_16954_, _11011_, _04613_);
  or (_16955_, _16954_, _16937_);
  and (_16956_, _16955_, _02799_);
  or (_16957_, _16956_, _16953_);
  or (_16958_, _16957_, _02928_);
  or (_16959_, _16958_, _16951_);
  or (_16960_, _16945_, _02943_);
  and (_16961_, _16960_, _16959_);
  or (_16962_, _16961_, _02796_);
  and (_16964_, _11009_, _04613_);
  or (_16965_, _16964_, _16937_);
  or (_16966_, _16965_, _02927_);
  and (_16967_, _16966_, _06189_);
  and (_16968_, _16967_, _16962_);
  or (_16969_, _16937_, _11040_);
  and (_16970_, _16955_, _02790_);
  and (_16971_, _16970_, _16969_);
  or (_16972_, _16971_, _02785_);
  or (_16973_, _16972_, _16968_);
  and (_16975_, _16973_, _16939_);
  or (_16976_, _16975_, _03861_);
  and (_16977_, _16976_, _16934_);
  or (_16978_, _16977_, _03850_);
  and (_16979_, _06116_, _04673_);
  or (_16980_, _16927_, _06726_);
  or (_16981_, _16980_, _16979_);
  and (_16982_, _16981_, _02970_);
  and (_16983_, _16982_, _16978_);
  nor (_16984_, _11114_, _08395_);
  or (_16986_, _16984_, _16927_);
  and (_16987_, _16986_, _02524_);
  or (_16988_, _16987_, _02974_);
  or (_16989_, _16988_, _16983_);
  and (_16990_, _04673_, _05616_);
  or (_16991_, _16990_, _16927_);
  or (_16992_, _16991_, _05261_);
  and (_16993_, _16992_, _16989_);
  or (_16994_, _16993_, _02977_);
  and (_16995_, _11128_, _04673_);
  or (_16997_, _16927_, _07092_);
  or (_16998_, _16997_, _16995_);
  and (_16999_, _16998_, _07104_);
  and (_17000_, _16999_, _16994_);
  or (_17001_, _17000_, _16931_);
  and (_17002_, _17001_, _03095_);
  or (_17003_, _16927_, _04939_);
  and (_17004_, _16945_, _03094_);
  and (_17005_, _16991_, _02991_);
  or (_17006_, _17005_, _17004_);
  and (_17008_, _17006_, _17003_);
  or (_17009_, _17008_, _02994_);
  or (_17010_, _17009_, _17002_);
  nor (_17011_, _11127_, _08395_);
  or (_17012_, _16927_, _07120_);
  or (_17013_, _17012_, _17011_);
  and (_17014_, _17013_, _07118_);
  and (_17015_, _17014_, _17010_);
  nor (_17016_, _11133_, _08395_);
  or (_17017_, _17016_, _16927_);
  and (_17019_, _17017_, _03099_);
  or (_17020_, _17019_, _03133_);
  or (_17021_, _17020_, _17015_);
  or (_17022_, _16942_, _03138_);
  and (_17023_, _17022_, _03142_);
  and (_17024_, _17023_, _17021_);
  and (_17025_, _16965_, _02778_);
  or (_17026_, _17025_, _02852_);
  or (_17027_, _17026_, _17024_);
  and (_17028_, _11185_, _04673_);
  or (_17030_, _16927_, _02853_);
  or (_17031_, _17030_, _17028_);
  and (_17032_, _17031_, _34446_);
  and (_17033_, _17032_, _17027_);
  or (_35621_[3], _17033_, _16926_);
  not (_17034_, \oc8051_golden_model_1.P0 [4]);
  nor (_17035_, _34446_, _17034_);
  or (_17036_, _17035_, rst);
  nor (_17037_, _04673_, _17034_);
  and (_17038_, _11333_, _04673_);
  or (_17040_, _17038_, _17037_);
  and (_17041_, _17040_, _03107_);
  nor (_17042_, _05143_, _08395_);
  or (_17043_, _17042_, _17037_);
  or (_17044_, _17043_, _03860_);
  nor (_17045_, _04613_, _17034_);
  and (_17046_, _11224_, _04613_);
  or (_17047_, _17046_, _17045_);
  or (_17048_, _17045_, _11239_);
  and (_17049_, _17048_, _02790_);
  and (_17051_, _17049_, _17047_);
  nor (_17052_, _11207_, _08395_);
  or (_17053_, _17052_, _17037_);
  or (_17054_, _17053_, _06162_);
  and (_17055_, _04673_, \oc8051_golden_model_1.ACC [4]);
  or (_17056_, _17055_, _17037_);
  and (_17057_, _17056_, _02837_);
  nor (_17058_, _02837_, _17034_);
  or (_17059_, _17058_, _02932_);
  or (_17060_, _17059_, _17057_);
  and (_17062_, _17060_, _02939_);
  and (_17063_, _17062_, _17054_);
  and (_17064_, _17043_, _02930_);
  and (_17065_, _17047_, _02799_);
  or (_17066_, _17065_, _17064_);
  or (_17067_, _17066_, _02928_);
  or (_17068_, _17067_, _17063_);
  or (_17069_, _17056_, _02943_);
  and (_17070_, _17069_, _17068_);
  or (_17071_, _17070_, _02796_);
  and (_17073_, _11203_, _04613_);
  or (_17074_, _17073_, _17045_);
  or (_17075_, _17074_, _02927_);
  and (_17076_, _17075_, _06189_);
  and (_17077_, _17076_, _17071_);
  or (_17078_, _17077_, _17051_);
  and (_17079_, _17078_, _02966_);
  or (_17080_, _11256_, _11203_);
  and (_17081_, _17080_, _04613_);
  or (_17082_, _17081_, _17045_);
  and (_17083_, _17082_, _02785_);
  or (_17084_, _17083_, _03861_);
  or (_17085_, _17084_, _17079_);
  and (_17086_, _17085_, _17044_);
  or (_17087_, _17086_, _03850_);
  and (_17088_, _06121_, _04673_);
  or (_17089_, _17037_, _06726_);
  or (_17090_, _17089_, _17088_);
  and (_17091_, _17090_, _02970_);
  and (_17092_, _17091_, _17087_);
  nor (_17095_, _11313_, _08395_);
  or (_17096_, _17095_, _17037_);
  and (_17097_, _17096_, _02524_);
  or (_17098_, _17097_, _02974_);
  or (_17099_, _17098_, _17092_);
  and (_17100_, _05629_, _04673_);
  or (_17101_, _17100_, _17037_);
  or (_17102_, _17101_, _05261_);
  and (_17103_, _17102_, _17099_);
  or (_17104_, _17103_, _02977_);
  and (_17105_, _11327_, _04673_);
  or (_17106_, _17037_, _07092_);
  or (_17107_, _17106_, _17105_);
  and (_17108_, _17107_, _07104_);
  and (_17109_, _17108_, _17104_);
  or (_17110_, _17109_, _17041_);
  and (_17111_, _17110_, _03095_);
  or (_17112_, _17037_, _05190_);
  and (_17113_, _17056_, _03094_);
  and (_17114_, _17101_, _02991_);
  or (_17117_, _17114_, _17113_);
  and (_17118_, _17117_, _17112_);
  or (_17119_, _17118_, _02994_);
  or (_17120_, _17119_, _17111_);
  nor (_17121_, _11326_, _08395_);
  or (_17122_, _17037_, _07120_);
  or (_17123_, _17122_, _17121_);
  and (_17124_, _17123_, _07118_);
  and (_17125_, _17124_, _17120_);
  nor (_17126_, _11332_, _08395_);
  or (_17128_, _17126_, _17037_);
  and (_17129_, _17128_, _03099_);
  or (_17130_, _17129_, _03133_);
  or (_17131_, _17130_, _17125_);
  or (_17132_, _17053_, _03138_);
  and (_17133_, _17132_, _03142_);
  and (_17134_, _17133_, _17131_);
  and (_17135_, _17074_, _02778_);
  or (_17136_, _17135_, _02852_);
  or (_17137_, _17136_, _17134_);
  and (_17139_, _11383_, _04673_);
  or (_17140_, _17037_, _02853_);
  or (_17141_, _17140_, _17139_);
  and (_17142_, _17141_, _34446_);
  and (_17143_, _17142_, _17137_);
  or (_35621_[4], _17143_, _17036_);
  not (_17144_, \oc8051_golden_model_1.P0 [5]);
  nor (_17145_, _34446_, _17144_);
  or (_17146_, _17145_, rst);
  nor (_17147_, _04673_, _17144_);
  and (_17149_, _11531_, _04673_);
  or (_17150_, _17149_, _17147_);
  and (_17151_, _17150_, _03107_);
  nor (_17152_, _11408_, _08395_);
  or (_17153_, _17152_, _17147_);
  or (_17154_, _17153_, _06162_);
  and (_17155_, _04673_, \oc8051_golden_model_1.ACC [5]);
  or (_17156_, _17155_, _17147_);
  and (_17157_, _17156_, _02837_);
  nor (_17158_, _02837_, _17144_);
  or (_17160_, _17158_, _02932_);
  or (_17161_, _17160_, _17157_);
  and (_17162_, _17161_, _02939_);
  and (_17163_, _17162_, _17154_);
  nor (_17164_, _04839_, _08395_);
  or (_17165_, _17164_, _17147_);
  and (_17166_, _17165_, _02930_);
  nor (_17167_, _04613_, _17144_);
  and (_17168_, _11422_, _04613_);
  or (_17169_, _17168_, _17167_);
  and (_17171_, _17169_, _02799_);
  or (_17172_, _17171_, _17166_);
  or (_17173_, _17172_, _02928_);
  or (_17174_, _17173_, _17163_);
  or (_17175_, _17156_, _02943_);
  and (_17176_, _17175_, _17174_);
  or (_17177_, _17176_, _02796_);
  and (_17178_, _11405_, _04613_);
  or (_17179_, _17178_, _17167_);
  or (_17180_, _17179_, _02927_);
  and (_17182_, _17180_, _06189_);
  and (_17183_, _17182_, _17177_);
  and (_17184_, _11438_, _04613_);
  or (_17185_, _17184_, _17167_);
  and (_17186_, _17185_, _02790_);
  or (_17187_, _17186_, _17183_);
  and (_17188_, _17187_, _02966_);
  or (_17189_, _11454_, _11405_);
  and (_17190_, _17189_, _04613_);
  or (_17191_, _17190_, _17167_);
  and (_17193_, _17191_, _02785_);
  or (_17194_, _17193_, _03861_);
  or (_17195_, _17194_, _17188_);
  or (_17196_, _17165_, _03860_);
  and (_17197_, _17196_, _17195_);
  or (_17198_, _17197_, _03850_);
  and (_17199_, _06120_, _04673_);
  or (_17200_, _17147_, _06726_);
  or (_17201_, _17200_, _17199_);
  and (_17202_, _17201_, _02970_);
  and (_17204_, _17202_, _17198_);
  nor (_17205_, _11511_, _08395_);
  or (_17206_, _17205_, _17147_);
  and (_17207_, _17206_, _02524_);
  or (_17208_, _17207_, _02974_);
  or (_17209_, _17208_, _17204_);
  and (_17210_, _05633_, _04673_);
  or (_17211_, _17210_, _17147_);
  or (_17212_, _17211_, _05261_);
  and (_17213_, _17212_, _17209_);
  or (_17215_, _17213_, _02977_);
  and (_17216_, _11525_, _04673_);
  or (_17217_, _17147_, _07092_);
  or (_17218_, _17217_, _17216_);
  and (_17219_, _17218_, _07104_);
  and (_17220_, _17219_, _17215_);
  or (_17221_, _17220_, _17151_);
  and (_17222_, _17221_, _03095_);
  or (_17223_, _17147_, _04890_);
  and (_17224_, _17156_, _03094_);
  and (_17226_, _17211_, _02991_);
  or (_17227_, _17226_, _17224_);
  and (_17228_, _17227_, _17223_);
  or (_17229_, _17228_, _02994_);
  or (_17230_, _17229_, _17222_);
  nor (_17231_, _11524_, _08395_);
  or (_17232_, _17147_, _07120_);
  or (_17233_, _17232_, _17231_);
  and (_17234_, _17233_, _07118_);
  and (_17235_, _17234_, _17230_);
  nor (_17237_, _11530_, _08395_);
  or (_17238_, _17237_, _17147_);
  and (_17239_, _17238_, _03099_);
  or (_17240_, _17239_, _03133_);
  or (_17241_, _17240_, _17235_);
  or (_17242_, _17153_, _03138_);
  and (_17243_, _17242_, _03142_);
  and (_17244_, _17243_, _17241_);
  and (_17245_, _17179_, _02778_);
  or (_17246_, _17245_, _02852_);
  or (_17248_, _17246_, _17244_);
  and (_17249_, _11580_, _04673_);
  or (_17250_, _17147_, _02853_);
  or (_17251_, _17250_, _17249_);
  and (_17252_, _17251_, _34446_);
  and (_17253_, _17252_, _17248_);
  or (_35621_[5], _17253_, _17146_);
  not (_17254_, \oc8051_golden_model_1.P0 [6]);
  nor (_17255_, _34446_, _17254_);
  or (_17256_, _17255_, rst);
  nor (_17258_, _04673_, _17254_);
  and (_17259_, _11601_, _04673_);
  or (_17260_, _17259_, _17258_);
  and (_17261_, _17260_, _03107_);
  nor (_17262_, _04735_, _08395_);
  or (_17263_, _17262_, _17258_);
  or (_17264_, _17263_, _03860_);
  nor (_17265_, _04613_, _17254_);
  and (_17266_, _11604_, _04613_);
  or (_17267_, _17266_, _17265_);
  or (_17269_, _17265_, _11603_);
  and (_17270_, _17269_, _02790_);
  and (_17271_, _17270_, _17267_);
  nor (_17272_, _11610_, _08395_);
  or (_17273_, _17272_, _17258_);
  or (_17274_, _17273_, _06162_);
  and (_17275_, _04673_, \oc8051_golden_model_1.ACC [6]);
  or (_17276_, _17275_, _17258_);
  and (_17277_, _17276_, _02837_);
  nor (_17278_, _02837_, _17254_);
  or (_17280_, _17278_, _02932_);
  or (_17281_, _17280_, _17277_);
  and (_17282_, _17281_, _02939_);
  and (_17283_, _17282_, _17274_);
  and (_17284_, _17263_, _02930_);
  and (_17285_, _17267_, _02799_);
  or (_17286_, _17285_, _17284_);
  or (_17287_, _17286_, _02928_);
  or (_17288_, _17287_, _17283_);
  or (_17289_, _17276_, _02943_);
  and (_17291_, _17289_, _17288_);
  or (_17292_, _17291_, _02796_);
  and (_17293_, _11633_, _04613_);
  or (_17294_, _17293_, _17265_);
  or (_17295_, _17294_, _02927_);
  and (_17296_, _17295_, _06189_);
  and (_17297_, _17296_, _17292_);
  or (_17298_, _17297_, _17271_);
  and (_17299_, _17298_, _02966_);
  or (_17300_, _11654_, _11633_);
  and (_17302_, _17300_, _04613_);
  or (_17303_, _17302_, _17265_);
  and (_17304_, _17303_, _02785_);
  or (_17305_, _17304_, _03861_);
  or (_17306_, _17305_, _17299_);
  and (_17307_, _17306_, _17264_);
  or (_17308_, _17307_, _03850_);
  and (_17309_, _05798_, _04673_);
  or (_17310_, _17258_, _06726_);
  or (_17311_, _17310_, _17309_);
  and (_17313_, _17311_, _02970_);
  and (_17314_, _17313_, _17308_);
  nor (_17315_, _11711_, _08395_);
  or (_17316_, _17315_, _17258_);
  and (_17317_, _17316_, _02524_);
  or (_17318_, _17317_, _02974_);
  or (_17319_, _17318_, _17314_);
  and (_17320_, _11718_, _04673_);
  or (_17321_, _17320_, _17258_);
  or (_17322_, _17321_, _05261_);
  and (_17324_, _17322_, _17319_);
  or (_17325_, _17324_, _02977_);
  and (_17326_, _11728_, _04673_);
  or (_17327_, _17258_, _07092_);
  or (_17328_, _17327_, _17326_);
  and (_17329_, _17328_, _07104_);
  and (_17330_, _17329_, _17325_);
  or (_17331_, _17330_, _17261_);
  and (_17332_, _17331_, _03095_);
  or (_17333_, _17258_, _04784_);
  and (_17335_, _17276_, _03094_);
  and (_17336_, _17321_, _02991_);
  or (_17337_, _17336_, _17335_);
  and (_17338_, _17337_, _17333_);
  or (_17339_, _17338_, _02994_);
  or (_17340_, _17339_, _17332_);
  nor (_17341_, _11726_, _08395_);
  or (_17342_, _17258_, _07120_);
  or (_17343_, _17342_, _17341_);
  and (_17344_, _17343_, _07118_);
  and (_17346_, _17344_, _17340_);
  nor (_17347_, _11600_, _08395_);
  or (_17348_, _17347_, _17258_);
  and (_17349_, _17348_, _03099_);
  or (_17350_, _17349_, _03133_);
  or (_17351_, _17350_, _17346_);
  or (_17352_, _17273_, _03138_);
  and (_17353_, _17352_, _03142_);
  and (_17354_, _17353_, _17351_);
  and (_17355_, _17294_, _02778_);
  or (_17357_, _17355_, _02852_);
  or (_17358_, _17357_, _17354_);
  and (_17359_, _11778_, _04673_);
  or (_17360_, _17258_, _02853_);
  or (_17361_, _17360_, _17359_);
  and (_17362_, _17361_, _34446_);
  and (_17363_, _17362_, _17358_);
  or (_35621_[6], _17363_, _17256_);
  not (_17364_, \oc8051_golden_model_1.P1 [0]);
  nor (_17365_, _34446_, _17364_);
  or (_17367_, _17365_, rst);
  nor (_17368_, _04676_, _17364_);
  and (_17369_, _10546_, _04676_);
  or (_17370_, _17369_, _17368_);
  and (_17371_, _17370_, _03107_);
  and (_17372_, _04676_, _03805_);
  or (_17373_, _17372_, _17368_);
  or (_17374_, _17373_, _03860_);
  nor (_17375_, _05300_, _17364_);
  and (_17376_, _10441_, _05300_);
  or (_17378_, _17376_, _17375_);
  and (_17379_, _17378_, _02799_);
  nor (_17380_, _05036_, _08490_);
  or (_17381_, _17380_, _17368_);
  or (_17382_, _17381_, _06162_);
  and (_17383_, _04676_, \oc8051_golden_model_1.ACC [0]);
  or (_17384_, _17383_, _17368_);
  and (_17385_, _17384_, _02837_);
  nor (_17386_, _02837_, _17364_);
  or (_17387_, _17386_, _02932_);
  or (_17389_, _17387_, _17385_);
  and (_17390_, _17389_, _02939_);
  and (_17391_, _17390_, _17382_);
  and (_17392_, _17373_, _02930_);
  or (_17393_, _17392_, _02928_);
  or (_17394_, _17393_, _17391_);
  or (_17395_, _17394_, _17379_);
  or (_17396_, _17384_, _02943_);
  and (_17397_, _17396_, _02927_);
  and (_17398_, _17397_, _17395_);
  and (_17400_, _17368_, _02796_);
  or (_17401_, _17400_, _02790_);
  or (_17402_, _17401_, _17398_);
  or (_17403_, _17381_, _06189_);
  and (_17404_, _17403_, _02966_);
  and (_17405_, _17404_, _17402_);
  and (_17406_, _16640_, _05300_);
  or (_17407_, _17406_, _17375_);
  and (_17408_, _17407_, _02785_);
  or (_17409_, _17408_, _03861_);
  or (_17411_, _17409_, _17405_);
  and (_17412_, _17411_, _17374_);
  or (_17413_, _17412_, _03850_);
  and (_17414_, _06114_, _04676_);
  or (_17415_, _17368_, _06726_);
  or (_17416_, _17415_, _17414_);
  and (_17417_, _17416_, _02970_);
  and (_17418_, _17417_, _17413_);
  nor (_17419_, _10530_, _08490_);
  or (_17420_, _17419_, _17368_);
  and (_17422_, _17420_, _02524_);
  or (_17423_, _17422_, _02974_);
  or (_17424_, _17423_, _17418_);
  and (_17425_, _04676_, _05647_);
  or (_17426_, _17425_, _17368_);
  or (_17427_, _17426_, _05261_);
  and (_17428_, _17427_, _17424_);
  or (_17429_, _17428_, _02977_);
  and (_17430_, _10427_, _04676_);
  or (_17431_, _17368_, _07092_);
  or (_17433_, _17431_, _17430_);
  and (_17434_, _17433_, _07104_);
  and (_17435_, _17434_, _17429_);
  or (_17436_, _17435_, _17371_);
  and (_17437_, _17436_, _03095_);
  nand (_17438_, _17426_, _02991_);
  nor (_17439_, _17438_, _17380_);
  or (_17440_, _17368_, _05036_);
  and (_17441_, _17384_, _03094_);
  and (_17442_, _17441_, _17440_);
  or (_17444_, _17442_, _02994_);
  or (_17445_, _17444_, _17439_);
  or (_17446_, _17445_, _17437_);
  nor (_17447_, _10425_, _08490_);
  or (_17448_, _17368_, _07120_);
  or (_17449_, _17448_, _17447_);
  and (_17450_, _17449_, _07118_);
  and (_17451_, _17450_, _17446_);
  nor (_17452_, _10423_, _08490_);
  or (_17453_, _17452_, _17368_);
  and (_17455_, _17453_, _03099_);
  or (_17456_, _17455_, _03133_);
  or (_17457_, _17456_, _17451_);
  or (_17458_, _17381_, _03138_);
  and (_17459_, _17458_, _03142_);
  and (_17460_, _17459_, _17457_);
  and (_17461_, _17368_, _02778_);
  or (_17462_, _17461_, _02852_);
  or (_17463_, _17462_, _17460_);
  or (_17464_, _17381_, _02853_);
  and (_17466_, _17464_, _34446_);
  and (_17467_, _17466_, _17463_);
  or (_35623_[0], _17467_, _17367_);
  not (_17468_, \oc8051_golden_model_1.P1 [1]);
  nor (_17469_, _34446_, _17468_);
  or (_17470_, _17469_, rst);
  nand (_17471_, _04676_, _03660_);
  or (_17472_, _04676_, \oc8051_golden_model_1.P1 [1]);
  and (_17473_, _17472_, _02974_);
  and (_17474_, _17473_, _17471_);
  nand (_17476_, _10719_, _04676_);
  and (_17477_, _17472_, _02524_);
  and (_17478_, _17477_, _17476_);
  and (_17479_, _16710_, _05300_);
  nor (_17480_, _05300_, _17468_);
  or (_17481_, _17480_, _02966_);
  or (_17482_, _17481_, _17479_);
  and (_17483_, _10622_, _04676_);
  not (_17484_, _17483_);
  and (_17485_, _17484_, _17472_);
  or (_17487_, _17485_, _06162_);
  nand (_17488_, _04676_, _02477_);
  and (_17489_, _17488_, _17472_);
  and (_17490_, _17489_, _02837_);
  nor (_17491_, _02837_, _17468_);
  or (_17492_, _17491_, _02932_);
  or (_17493_, _17492_, _17490_);
  and (_17494_, _17493_, _02939_);
  and (_17495_, _17494_, _17487_);
  nor (_17496_, _04676_, _17468_);
  nor (_17498_, _08490_, _03989_);
  or (_17499_, _17498_, _17496_);
  and (_17500_, _17499_, _02930_);
  and (_17501_, _10617_, _05300_);
  or (_17502_, _17501_, _17480_);
  and (_17503_, _17502_, _02799_);
  or (_17504_, _17503_, _17500_);
  or (_17505_, _17504_, _02928_);
  or (_17506_, _17505_, _17495_);
  or (_17507_, _17489_, _02943_);
  and (_17509_, _17507_, _17506_);
  or (_17510_, _17509_, _02796_);
  and (_17511_, _10620_, _05300_);
  or (_17512_, _17511_, _17480_);
  or (_17513_, _17512_, _02927_);
  and (_17514_, _17513_, _06189_);
  and (_17515_, _17514_, _17510_);
  and (_17516_, _17501_, _10616_);
  or (_17517_, _17516_, _17480_);
  and (_17518_, _17517_, _02790_);
  or (_17520_, _17518_, _02785_);
  or (_17521_, _17520_, _17515_);
  and (_17522_, _17521_, _17482_);
  or (_17523_, _17522_, _03861_);
  or (_17524_, _17499_, _03860_);
  and (_17525_, _17524_, _17523_);
  or (_17526_, _17525_, _03850_);
  and (_17527_, _06113_, _04676_);
  or (_17528_, _17496_, _06726_);
  or (_17529_, _17528_, _17527_);
  and (_17531_, _17529_, _02970_);
  and (_17532_, _17531_, _17526_);
  or (_17533_, _17532_, _17478_);
  and (_17534_, _17533_, _05261_);
  or (_17535_, _17534_, _17474_);
  and (_17536_, _17535_, _03882_);
  or (_17537_, _10613_, _08490_);
  and (_17538_, _17472_, _02991_);
  and (_17539_, _17538_, _17537_);
  or (_17540_, _10610_, _08490_);
  and (_17542_, _17472_, _03107_);
  and (_17543_, _17542_, _17540_);
  or (_17544_, _10614_, _08490_);
  and (_17545_, _17472_, _02977_);
  and (_17546_, _17545_, _17544_);
  or (_17547_, _17546_, _17543_);
  or (_17548_, _17547_, _17539_);
  or (_17549_, _17548_, _17536_);
  and (_17550_, _17549_, _06161_);
  or (_17551_, _17496_, _04988_);
  and (_17553_, _17489_, _03094_);
  and (_17554_, _17553_, _17551_);
  or (_17555_, _17554_, _17550_);
  and (_17556_, _17555_, _03100_);
  or (_17557_, _17471_, _04988_);
  and (_17558_, _17472_, _02994_);
  and (_17559_, _17558_, _17557_);
  or (_17560_, _17488_, _04988_);
  and (_17561_, _17472_, _03099_);
  and (_17562_, _17561_, _17560_);
  or (_17564_, _17562_, _03133_);
  or (_17565_, _17564_, _17559_);
  or (_17566_, _17565_, _17556_);
  or (_17567_, _17485_, _03138_);
  and (_17568_, _17567_, _03142_);
  and (_17569_, _17568_, _17566_);
  and (_17570_, _17512_, _02778_);
  or (_17571_, _17570_, _02852_);
  or (_17572_, _17571_, _17569_);
  or (_17573_, _17496_, _02853_);
  or (_17575_, _17573_, _17483_);
  and (_17576_, _17575_, _34446_);
  and (_17577_, _17576_, _17572_);
  or (_35623_[1], _17577_, _17470_);
  not (_17578_, \oc8051_golden_model_1.P1 [2]);
  nor (_17579_, _34446_, _17578_);
  or (_17580_, _17579_, rst);
  nor (_17581_, _04676_, _17578_);
  and (_17582_, _10942_, _04676_);
  or (_17583_, _17582_, _17581_);
  and (_17585_, _17583_, _03107_);
  nor (_17586_, _08490_, _04413_);
  or (_17587_, _17586_, _17581_);
  or (_17588_, _17587_, _03860_);
  nor (_17589_, _10824_, _08490_);
  or (_17590_, _17589_, _17581_);
  or (_17591_, _17590_, _06162_);
  and (_17592_, _04676_, \oc8051_golden_model_1.ACC [2]);
  or (_17593_, _17592_, _17581_);
  and (_17594_, _17593_, _02837_);
  nor (_17596_, _02837_, _17578_);
  or (_17597_, _17596_, _02932_);
  or (_17598_, _17597_, _17594_);
  and (_17599_, _17598_, _02939_);
  and (_17600_, _17599_, _17591_);
  and (_17601_, _17587_, _02930_);
  nor (_17602_, _05300_, _17578_);
  and (_17603_, _10815_, _05300_);
  or (_17604_, _17603_, _17602_);
  and (_17605_, _17604_, _02799_);
  or (_17607_, _17605_, _17601_);
  or (_17608_, _17607_, _02928_);
  or (_17609_, _17608_, _17600_);
  or (_17610_, _17593_, _02943_);
  and (_17611_, _17610_, _17609_);
  or (_17612_, _17611_, _02796_);
  and (_17613_, _10818_, _05300_);
  or (_17614_, _17613_, _17602_);
  or (_17615_, _17614_, _02927_);
  and (_17616_, _17615_, _06189_);
  and (_17618_, _17616_, _17612_);
  and (_17619_, _17603_, _10814_);
  or (_17620_, _17619_, _17602_);
  and (_17621_, _17620_, _02790_);
  or (_17622_, _17621_, _17618_);
  and (_17623_, _17622_, _02966_);
  and (_17624_, _16860_, _05300_);
  or (_17625_, _17602_, _17624_);
  and (_17626_, _17625_, _02785_);
  or (_17627_, _17626_, _03861_);
  or (_17629_, _17627_, _17623_);
  and (_17630_, _17629_, _17588_);
  or (_17631_, _17630_, _03850_);
  and (_17632_, _06117_, _04676_);
  or (_17633_, _17581_, _06726_);
  or (_17634_, _17633_, _17632_);
  and (_17635_, _17634_, _02970_);
  and (_17636_, _17635_, _17631_);
  nor (_17637_, _10922_, _08490_);
  or (_17638_, _17637_, _17581_);
  and (_17640_, _17638_, _02524_);
  or (_17641_, _17640_, _02974_);
  or (_17642_, _17641_, _17636_);
  and (_17643_, _04676_, _05690_);
  or (_17644_, _17643_, _17581_);
  or (_17645_, _17644_, _05261_);
  and (_17646_, _17645_, _17642_);
  or (_17647_, _17646_, _02977_);
  and (_17648_, _10936_, _04676_);
  or (_17649_, _17581_, _07092_);
  or (_17651_, _17649_, _17648_);
  and (_17652_, _17651_, _07104_);
  and (_17653_, _17652_, _17647_);
  or (_17654_, _17653_, _17585_);
  and (_17655_, _17654_, _03095_);
  or (_17656_, _17581_, _05086_);
  and (_17657_, _17593_, _03094_);
  and (_17658_, _17644_, _02991_);
  or (_17659_, _17658_, _17657_);
  and (_17660_, _17659_, _17656_);
  or (_17662_, _17660_, _02994_);
  or (_17663_, _17662_, _17655_);
  nor (_17664_, _10935_, _08490_);
  or (_17665_, _17581_, _07120_);
  or (_17666_, _17665_, _17664_);
  and (_17667_, _17666_, _07118_);
  and (_17668_, _17667_, _17663_);
  nor (_17669_, _10941_, _08490_);
  or (_17670_, _17669_, _17581_);
  and (_17671_, _17670_, _03099_);
  or (_17673_, _17671_, _03133_);
  or (_17674_, _17673_, _17668_);
  or (_17675_, _17590_, _03138_);
  and (_17676_, _17675_, _03142_);
  and (_17677_, _17676_, _17674_);
  and (_17678_, _17614_, _02778_);
  or (_17679_, _17678_, _02852_);
  or (_17680_, _17679_, _17677_);
  and (_17681_, _10988_, _04676_);
  or (_17682_, _17581_, _02853_);
  or (_17684_, _17682_, _17681_);
  and (_17685_, _17684_, _34446_);
  and (_17686_, _17685_, _17680_);
  or (_35623_[2], _17686_, _17580_);
  nor (_17687_, \oc8051_golden_model_1.P1 [3], rst);
  nor (_17688_, _17687_, _04509_);
  and (_17689_, _08490_, \oc8051_golden_model_1.P1 [3]);
  and (_17690_, _11134_, _04676_);
  or (_17691_, _17690_, _17689_);
  and (_17692_, _17691_, _03107_);
  nor (_17694_, _08490_, _04226_);
  or (_17695_, _17694_, _17689_);
  or (_17696_, _17695_, _03860_);
  and (_17697_, _16935_, _05300_);
  not (_17698_, _05300_);
  and (_17699_, _17698_, \oc8051_golden_model_1.P1 [3]);
  or (_17700_, _17699_, _02966_);
  or (_17701_, _17700_, _17697_);
  nor (_17702_, _11014_, _08490_);
  or (_17703_, _17702_, _17689_);
  or (_17705_, _17703_, _06162_);
  and (_17706_, _04676_, \oc8051_golden_model_1.ACC [3]);
  or (_17707_, _17706_, _17689_);
  and (_17708_, _17707_, _02837_);
  and (_17709_, _09167_, \oc8051_golden_model_1.P1 [3]);
  or (_17710_, _17709_, _02932_);
  or (_17711_, _17710_, _17708_);
  and (_17712_, _17711_, _02939_);
  and (_17713_, _17712_, _17705_);
  and (_17714_, _17695_, _02930_);
  and (_17716_, _11011_, _05300_);
  or (_17717_, _17716_, _17699_);
  and (_17718_, _17717_, _02799_);
  or (_17719_, _17718_, _17714_);
  or (_17720_, _17719_, _02928_);
  or (_17721_, _17720_, _17713_);
  or (_17722_, _17707_, _02943_);
  and (_17723_, _17722_, _17721_);
  or (_17724_, _17723_, _02796_);
  and (_17725_, _11009_, _05300_);
  or (_17727_, _17725_, _17699_);
  or (_17728_, _17727_, _02927_);
  and (_17729_, _17728_, _06189_);
  and (_17730_, _17729_, _17724_);
  or (_17731_, _17699_, _11040_);
  and (_17732_, _17731_, _02790_);
  and (_17733_, _17732_, _17717_);
  or (_17734_, _17733_, _02785_);
  or (_17735_, _17734_, _17730_);
  and (_17736_, _17735_, _17701_);
  or (_17738_, _17736_, _03861_);
  and (_17739_, _17738_, _17696_);
  or (_17740_, _17739_, _03850_);
  and (_17741_, _06116_, _04676_);
  or (_17742_, _17689_, _06726_);
  or (_17743_, _17742_, _17741_);
  and (_17744_, _17743_, _02970_);
  and (_17745_, _17744_, _17740_);
  nor (_17746_, _11114_, _08490_);
  or (_17747_, _17746_, _17689_);
  and (_17749_, _17747_, _02524_);
  or (_17750_, _17749_, _02974_);
  or (_17751_, _17750_, _17745_);
  and (_17752_, _04676_, _05616_);
  or (_17753_, _17752_, _17689_);
  or (_17754_, _17753_, _05261_);
  and (_17755_, _17754_, _17751_);
  or (_17756_, _17755_, _02977_);
  and (_17757_, _11128_, _04676_);
  or (_17758_, _17689_, _07092_);
  or (_17760_, _17758_, _17757_);
  and (_17761_, _17760_, _07104_);
  and (_17762_, _17761_, _17756_);
  or (_17763_, _17762_, _17692_);
  and (_17764_, _17763_, _03095_);
  or (_17765_, _17689_, _04939_);
  and (_17766_, _17707_, _03094_);
  and (_17767_, _17753_, _02991_);
  or (_17768_, _17767_, _17766_);
  and (_17769_, _17768_, _17765_);
  or (_17771_, _17769_, _02994_);
  or (_17772_, _17771_, _17764_);
  nor (_17773_, _11127_, _08490_);
  or (_17774_, _17689_, _07120_);
  or (_17775_, _17774_, _17773_);
  and (_17776_, _17775_, _07118_);
  and (_17777_, _17776_, _17772_);
  nor (_17778_, _11133_, _08490_);
  or (_17779_, _17778_, _17689_);
  and (_17780_, _17779_, _03099_);
  or (_17782_, _17780_, _03133_);
  or (_17783_, _17782_, _17777_);
  or (_17784_, _17703_, _03138_);
  and (_17785_, _17784_, _03142_);
  and (_17786_, _17785_, _17783_);
  and (_17787_, _17727_, _02778_);
  or (_17788_, _17787_, _02852_);
  or (_17789_, _17788_, _17786_);
  and (_17790_, _11185_, _04676_);
  or (_17791_, _17689_, _02853_);
  or (_17793_, _17791_, _17790_);
  and (_17794_, _17793_, _34446_);
  and (_17795_, _17794_, _17789_);
  or (_35623_[3], _17795_, _17688_);
  nor (_17796_, \oc8051_golden_model_1.P1 [4], rst);
  nor (_17797_, _17796_, _04509_);
  and (_17798_, _08490_, \oc8051_golden_model_1.P1 [4]);
  and (_17799_, _11333_, _04676_);
  or (_17800_, _17799_, _17798_);
  and (_17801_, _17800_, _03107_);
  nor (_17803_, _05143_, _08490_);
  or (_17804_, _17803_, _17798_);
  or (_17805_, _17804_, _03860_);
  and (_17806_, _17698_, \oc8051_golden_model_1.P1 [4]);
  and (_17807_, _11224_, _05300_);
  or (_17808_, _17807_, _17806_);
  or (_17809_, _17806_, _11239_);
  and (_17810_, _17809_, _02790_);
  and (_17811_, _17810_, _17808_);
  nor (_17812_, _11207_, _08490_);
  or (_17814_, _17812_, _17798_);
  or (_17815_, _17814_, _06162_);
  and (_17816_, _04676_, \oc8051_golden_model_1.ACC [4]);
  or (_17817_, _17816_, _17798_);
  and (_17818_, _17817_, _02837_);
  and (_17819_, _09167_, \oc8051_golden_model_1.P1 [4]);
  or (_17820_, _17819_, _02932_);
  or (_17821_, _17820_, _17818_);
  and (_17822_, _17821_, _02939_);
  and (_17823_, _17822_, _17815_);
  and (_17825_, _17804_, _02930_);
  and (_17826_, _17808_, _02799_);
  or (_17827_, _17826_, _17825_);
  or (_17828_, _17827_, _02928_);
  or (_17829_, _17828_, _17823_);
  or (_17830_, _17817_, _02943_);
  and (_17831_, _17830_, _17829_);
  or (_17832_, _17831_, _02796_);
  and (_17833_, _11203_, _05300_);
  or (_17834_, _17833_, _17806_);
  or (_17836_, _17834_, _02927_);
  and (_17837_, _17836_, _06189_);
  and (_17838_, _17837_, _17832_);
  or (_17839_, _17838_, _17811_);
  and (_17840_, _17839_, _02966_);
  and (_17841_, _17080_, _05300_);
  or (_17842_, _17841_, _17806_);
  and (_17843_, _17842_, _02785_);
  or (_17844_, _17843_, _03861_);
  or (_17845_, _17844_, _17840_);
  and (_17847_, _17845_, _17805_);
  or (_17848_, _17847_, _03850_);
  and (_17849_, _06121_, _04676_);
  or (_17850_, _17798_, _06726_);
  or (_17851_, _17850_, _17849_);
  and (_17852_, _17851_, _02970_);
  and (_17853_, _17852_, _17848_);
  nor (_17854_, _11313_, _08490_);
  or (_17855_, _17854_, _17798_);
  and (_17856_, _17855_, _02524_);
  or (_17858_, _17856_, _02974_);
  or (_17859_, _17858_, _17853_);
  and (_17860_, _05629_, _04676_);
  or (_17861_, _17860_, _17798_);
  or (_17862_, _17861_, _05261_);
  and (_17863_, _17862_, _17859_);
  or (_17864_, _17863_, _02977_);
  and (_17865_, _11327_, _04676_);
  or (_17866_, _17798_, _07092_);
  or (_17867_, _17866_, _17865_);
  and (_17869_, _17867_, _07104_);
  and (_17870_, _17869_, _17864_);
  or (_17871_, _17870_, _17801_);
  and (_17872_, _17871_, _03095_);
  or (_17873_, _17798_, _05190_);
  and (_17874_, _17817_, _03094_);
  and (_17875_, _17861_, _02991_);
  or (_17876_, _17875_, _17874_);
  and (_17877_, _17876_, _17873_);
  or (_17878_, _17877_, _02994_);
  or (_17880_, _17878_, _17872_);
  nor (_17881_, _11326_, _08490_);
  or (_17882_, _17798_, _07120_);
  or (_17883_, _17882_, _17881_);
  and (_17884_, _17883_, _07118_);
  and (_17885_, _17884_, _17880_);
  nor (_17886_, _11332_, _08490_);
  or (_17887_, _17886_, _17798_);
  and (_17888_, _17887_, _03099_);
  or (_17889_, _17888_, _03133_);
  or (_17891_, _17889_, _17885_);
  or (_17892_, _17814_, _03138_);
  and (_17893_, _17892_, _03142_);
  and (_17894_, _17893_, _17891_);
  and (_17895_, _17834_, _02778_);
  or (_17896_, _17895_, _02852_);
  or (_17897_, _17896_, _17894_);
  and (_17898_, _11383_, _04676_);
  or (_17899_, _17798_, _02853_);
  or (_17900_, _17899_, _17898_);
  and (_17902_, _17900_, _34446_);
  and (_17903_, _17902_, _17897_);
  or (_35623_[4], _17903_, _17797_);
  nor (_17904_, \oc8051_golden_model_1.P1 [5], rst);
  nor (_17905_, _17904_, _04509_);
  and (_17906_, _08490_, \oc8051_golden_model_1.P1 [5]);
  and (_17907_, _11531_, _04676_);
  or (_17908_, _17907_, _17906_);
  and (_17909_, _17908_, _03107_);
  nor (_17910_, _11408_, _08490_);
  or (_17912_, _17910_, _17906_);
  or (_17913_, _17912_, _06162_);
  and (_17914_, _04676_, \oc8051_golden_model_1.ACC [5]);
  or (_17915_, _17914_, _17906_);
  and (_17916_, _17915_, _02837_);
  and (_17917_, _09167_, \oc8051_golden_model_1.P1 [5]);
  or (_17918_, _17917_, _02932_);
  or (_17919_, _17918_, _17916_);
  and (_17920_, _17919_, _02939_);
  and (_17921_, _17920_, _17913_);
  nor (_17923_, _04839_, _08490_);
  or (_17924_, _17923_, _17906_);
  and (_17925_, _17924_, _02930_);
  and (_17926_, _17698_, \oc8051_golden_model_1.P1 [5]);
  and (_17927_, _11422_, _05300_);
  or (_17928_, _17927_, _17926_);
  and (_17929_, _17928_, _02799_);
  or (_17930_, _17929_, _17925_);
  or (_17931_, _17930_, _02928_);
  or (_17932_, _17931_, _17921_);
  or (_17934_, _17915_, _02943_);
  and (_17935_, _17934_, _17932_);
  or (_17936_, _17935_, _02796_);
  and (_17937_, _11405_, _05300_);
  or (_17938_, _17937_, _17926_);
  or (_17939_, _17938_, _02927_);
  and (_17940_, _17939_, _06189_);
  and (_17941_, _17940_, _17936_);
  and (_17942_, _11438_, _05300_);
  or (_17943_, _17942_, _17926_);
  and (_17945_, _17943_, _02790_);
  or (_17946_, _17945_, _17941_);
  and (_17947_, _17946_, _02966_);
  and (_17948_, _17189_, _05300_);
  or (_17949_, _17948_, _17926_);
  and (_17950_, _17949_, _02785_);
  or (_17951_, _17950_, _03861_);
  or (_17952_, _17951_, _17947_);
  or (_17953_, _17924_, _03860_);
  and (_17954_, _17953_, _17952_);
  or (_17956_, _17954_, _03850_);
  and (_17957_, _06120_, _04676_);
  or (_17958_, _17906_, _06726_);
  or (_17959_, _17958_, _17957_);
  and (_17960_, _17959_, _02970_);
  and (_17961_, _17960_, _17956_);
  nor (_17962_, _11511_, _08490_);
  or (_17963_, _17962_, _17906_);
  and (_17964_, _17963_, _02524_);
  or (_17965_, _17964_, _02974_);
  or (_17967_, _17965_, _17961_);
  and (_17968_, _05633_, _04676_);
  or (_17969_, _17968_, _17906_);
  or (_17970_, _17969_, _05261_);
  and (_17971_, _17970_, _17967_);
  or (_17972_, _17971_, _02977_);
  and (_17973_, _11525_, _04676_);
  or (_17974_, _17906_, _07092_);
  or (_17975_, _17974_, _17973_);
  and (_17976_, _17975_, _07104_);
  and (_17978_, _17976_, _17972_);
  or (_17979_, _17978_, _17909_);
  and (_17980_, _17979_, _03095_);
  or (_17981_, _17906_, _04890_);
  and (_17982_, _17915_, _03094_);
  and (_17983_, _17969_, _02991_);
  or (_17984_, _17983_, _17982_);
  and (_17985_, _17984_, _17981_);
  or (_17986_, _17985_, _02994_);
  or (_17987_, _17986_, _17980_);
  nor (_17989_, _11524_, _08490_);
  or (_17990_, _17906_, _07120_);
  or (_17991_, _17990_, _17989_);
  and (_17992_, _17991_, _07118_);
  and (_17993_, _17992_, _17987_);
  nor (_17994_, _11530_, _08490_);
  or (_17995_, _17994_, _17906_);
  and (_17996_, _17995_, _03099_);
  or (_17997_, _17996_, _03133_);
  or (_17998_, _17997_, _17993_);
  or (_18000_, _17912_, _03138_);
  and (_18001_, _18000_, _03142_);
  and (_18002_, _18001_, _17998_);
  and (_18003_, _17938_, _02778_);
  or (_18004_, _18003_, _02852_);
  or (_18005_, _18004_, _18002_);
  and (_18006_, _11580_, _04676_);
  or (_18007_, _17906_, _02853_);
  or (_18008_, _18007_, _18006_);
  and (_18009_, _18008_, _34446_);
  and (_18011_, _18009_, _18005_);
  or (_35623_[5], _18011_, _17905_);
  not (_18012_, \oc8051_golden_model_1.P1 [6]);
  nor (_18013_, _34446_, _18012_);
  or (_18014_, _18013_, rst);
  nor (_18015_, _04676_, _18012_);
  and (_18016_, _11601_, _04676_);
  or (_18017_, _18016_, _18015_);
  and (_18018_, _18017_, _03107_);
  nor (_18019_, _04735_, _08490_);
  or (_18021_, _18019_, _18015_);
  or (_18022_, _18021_, _03860_);
  nor (_18023_, _05300_, _18012_);
  and (_18024_, _11604_, _05300_);
  or (_18025_, _18024_, _18023_);
  or (_18026_, _18023_, _11603_);
  and (_18027_, _18026_, _02790_);
  and (_18028_, _18027_, _18025_);
  nor (_18029_, _11610_, _08490_);
  or (_18030_, _18029_, _18015_);
  or (_18032_, _18030_, _06162_);
  and (_18033_, _04676_, \oc8051_golden_model_1.ACC [6]);
  or (_18034_, _18033_, _18015_);
  and (_18035_, _18034_, _02837_);
  nor (_18036_, _02837_, _18012_);
  or (_18037_, _18036_, _02932_);
  or (_18038_, _18037_, _18035_);
  and (_18039_, _18038_, _02939_);
  and (_18040_, _18039_, _18032_);
  and (_18041_, _18021_, _02930_);
  and (_18043_, _18025_, _02799_);
  or (_18044_, _18043_, _18041_);
  or (_18045_, _18044_, _02928_);
  or (_18046_, _18045_, _18040_);
  or (_18047_, _18034_, _02943_);
  and (_18048_, _18047_, _18046_);
  or (_18049_, _18048_, _02796_);
  and (_18050_, _11633_, _05300_);
  or (_18051_, _18050_, _18023_);
  or (_18052_, _18051_, _02927_);
  and (_18054_, _18052_, _06189_);
  and (_18055_, _18054_, _18049_);
  or (_18056_, _18055_, _18028_);
  and (_18057_, _18056_, _02966_);
  and (_18058_, _17300_, _05300_);
  or (_18059_, _18058_, _18023_);
  and (_18060_, _18059_, _02785_);
  or (_18061_, _18060_, _03861_);
  or (_18062_, _18061_, _18057_);
  and (_18063_, _18062_, _18022_);
  or (_18065_, _18063_, _03850_);
  and (_18066_, _05798_, _04676_);
  or (_18067_, _18015_, _06726_);
  or (_18068_, _18067_, _18066_);
  and (_18069_, _18068_, _02970_);
  and (_18070_, _18069_, _18065_);
  nor (_18071_, _11711_, _08490_);
  or (_18072_, _18071_, _18015_);
  and (_18073_, _18072_, _02524_);
  or (_18074_, _18073_, _02974_);
  or (_18076_, _18074_, _18070_);
  and (_18077_, _11718_, _04676_);
  or (_18078_, _18077_, _18015_);
  or (_18079_, _18078_, _05261_);
  and (_18080_, _18079_, _18076_);
  or (_18081_, _18080_, _02977_);
  and (_18082_, _11728_, _04676_);
  or (_18083_, _18015_, _07092_);
  or (_18084_, _18083_, _18082_);
  and (_18085_, _18084_, _07104_);
  and (_18087_, _18085_, _18081_);
  or (_18088_, _18087_, _18018_);
  and (_18089_, _18088_, _03095_);
  or (_18090_, _18015_, _04784_);
  and (_18091_, _18034_, _03094_);
  and (_18092_, _18078_, _02991_);
  or (_18093_, _18092_, _18091_);
  and (_18094_, _18093_, _18090_);
  or (_18095_, _18094_, _02994_);
  or (_18096_, _18095_, _18089_);
  nor (_18098_, _11726_, _08490_);
  or (_18099_, _18015_, _07120_);
  or (_18100_, _18099_, _18098_);
  and (_18101_, _18100_, _07118_);
  and (_18102_, _18101_, _18096_);
  nor (_18103_, _11600_, _08490_);
  or (_18104_, _18103_, _18015_);
  and (_18105_, _18104_, _03099_);
  or (_18106_, _18105_, _03133_);
  or (_18107_, _18106_, _18102_);
  or (_18109_, _18030_, _03138_);
  and (_18110_, _18109_, _03142_);
  and (_18111_, _18110_, _18107_);
  and (_18112_, _18051_, _02778_);
  or (_18113_, _18112_, _02852_);
  or (_18114_, _18113_, _18111_);
  and (_18115_, _11778_, _04676_);
  or (_18116_, _18015_, _02853_);
  or (_18117_, _18116_, _18115_);
  and (_18118_, _18117_, _34446_);
  and (_18120_, _18118_, _18114_);
  or (_35623_[6], _18120_, _18014_);
  not (_18121_, \oc8051_golden_model_1.P2 [0]);
  nor (_18122_, _34446_, _18121_);
  or (_18123_, _18122_, rst);
  nor (_18124_, _04679_, _18121_);
  and (_18125_, _10546_, _04679_);
  or (_18126_, _18125_, _18124_);
  and (_18127_, _18126_, _03107_);
  and (_18128_, _04679_, _03805_);
  or (_18130_, _18128_, _18124_);
  or (_18131_, _18130_, _03860_);
  nor (_18132_, _05278_, _18121_);
  and (_18133_, _10441_, _05278_);
  or (_18134_, _18133_, _18132_);
  and (_18135_, _18134_, _02799_);
  nor (_18136_, _05036_, _08596_);
  or (_18137_, _18136_, _18124_);
  or (_18138_, _18137_, _06162_);
  and (_18139_, _04679_, \oc8051_golden_model_1.ACC [0]);
  or (_18141_, _18139_, _18124_);
  and (_18142_, _18141_, _02837_);
  nor (_18143_, _02837_, _18121_);
  or (_18144_, _18143_, _02932_);
  or (_18145_, _18144_, _18142_);
  and (_18146_, _18145_, _02939_);
  and (_18147_, _18146_, _18138_);
  and (_18148_, _18130_, _02930_);
  or (_18149_, _18148_, _02928_);
  or (_18150_, _18149_, _18147_);
  or (_18152_, _18150_, _18135_);
  or (_18153_, _18141_, _02943_);
  and (_18154_, _18153_, _02927_);
  and (_18155_, _18154_, _18152_);
  and (_18156_, _18124_, _02796_);
  or (_18157_, _18156_, _02790_);
  or (_18158_, _18157_, _18155_);
  or (_18159_, _18137_, _06189_);
  and (_18160_, _18159_, _02966_);
  and (_18161_, _18160_, _18158_);
  and (_18163_, _16640_, _05278_);
  or (_18164_, _18163_, _18132_);
  and (_18165_, _18164_, _02785_);
  or (_18166_, _18165_, _03861_);
  or (_18167_, _18166_, _18161_);
  and (_18168_, _18167_, _18131_);
  or (_18169_, _18168_, _03850_);
  and (_18170_, _06114_, _04679_);
  or (_18171_, _18124_, _06726_);
  or (_18172_, _18171_, _18170_);
  and (_18174_, _18172_, _02970_);
  and (_18175_, _18174_, _18169_);
  nor (_18176_, _10530_, _08596_);
  or (_18177_, _18176_, _18124_);
  and (_18178_, _18177_, _02524_);
  or (_18179_, _18178_, _02974_);
  or (_18180_, _18179_, _18175_);
  and (_18181_, _04679_, _05647_);
  or (_18182_, _18181_, _18124_);
  or (_18183_, _18182_, _05261_);
  and (_18185_, _18183_, _18180_);
  or (_18186_, _18185_, _02977_);
  and (_18187_, _10427_, _04679_);
  or (_18188_, _18124_, _07092_);
  or (_18189_, _18188_, _18187_);
  and (_18190_, _18189_, _07104_);
  and (_18191_, _18190_, _18186_);
  or (_18192_, _18191_, _18127_);
  and (_18193_, _18192_, _03095_);
  nand (_18194_, _18182_, _02991_);
  nor (_18196_, _18194_, _18136_);
  or (_18197_, _18124_, _05036_);
  and (_18198_, _18141_, _03094_);
  and (_18199_, _18198_, _18197_);
  or (_18200_, _18199_, _02994_);
  or (_18201_, _18200_, _18196_);
  or (_18202_, _18201_, _18193_);
  nor (_18203_, _10425_, _08596_);
  or (_18204_, _18124_, _07120_);
  or (_18205_, _18204_, _18203_);
  and (_18207_, _18205_, _07118_);
  and (_18208_, _18207_, _18202_);
  nor (_18209_, _10423_, _08596_);
  or (_18210_, _18209_, _18124_);
  and (_18211_, _18210_, _03099_);
  or (_18212_, _18211_, _03133_);
  or (_18213_, _18212_, _18208_);
  or (_18214_, _18137_, _03138_);
  and (_18215_, _18214_, _03142_);
  and (_18216_, _18215_, _18213_);
  and (_18218_, _18124_, _02778_);
  or (_18219_, _18218_, _02852_);
  or (_18220_, _18219_, _18216_);
  or (_18221_, _18137_, _02853_);
  and (_18222_, _18221_, _34446_);
  and (_18223_, _18222_, _18220_);
  or (_35625_[0], _18223_, _18123_);
  not (_18224_, \oc8051_golden_model_1.P2 [1]);
  nor (_18225_, _34446_, _18224_);
  or (_18226_, _18225_, rst);
  nand (_18228_, _04679_, _03660_);
  or (_18229_, _04679_, \oc8051_golden_model_1.P2 [1]);
  and (_18230_, _18229_, _02974_);
  and (_18231_, _18230_, _18228_);
  nand (_18232_, _10719_, _04679_);
  and (_18233_, _18229_, _02524_);
  and (_18234_, _18233_, _18232_);
  and (_18235_, _16710_, _05278_);
  nor (_18236_, _05278_, _18224_);
  or (_18237_, _18236_, _02966_);
  or (_18239_, _18237_, _18235_);
  and (_18240_, _10622_, _04679_);
  not (_18241_, _18240_);
  and (_18242_, _18241_, _18229_);
  or (_18243_, _18242_, _06162_);
  nand (_18244_, _04679_, _02477_);
  and (_18245_, _18244_, _18229_);
  and (_18246_, _18245_, _02837_);
  nor (_18247_, _02837_, _18224_);
  or (_18248_, _18247_, _02932_);
  or (_18250_, _18248_, _18246_);
  and (_18251_, _18250_, _02939_);
  and (_18252_, _18251_, _18243_);
  nor (_18253_, _04679_, _18224_);
  nor (_18254_, _08596_, _03989_);
  or (_18255_, _18254_, _18253_);
  and (_18256_, _18255_, _02930_);
  and (_18257_, _10617_, _05278_);
  or (_18258_, _18257_, _18236_);
  and (_18259_, _18258_, _02799_);
  or (_18261_, _18259_, _18256_);
  or (_18262_, _18261_, _02928_);
  or (_18263_, _18262_, _18252_);
  or (_18264_, _18245_, _02943_);
  and (_18265_, _18264_, _18263_);
  or (_18266_, _18265_, _02796_);
  and (_18267_, _10620_, _05278_);
  or (_18268_, _18267_, _18236_);
  or (_18269_, _18268_, _02927_);
  and (_18270_, _18269_, _06189_);
  and (_18272_, _18270_, _18266_);
  and (_18273_, _18257_, _10616_);
  or (_18274_, _18273_, _18236_);
  and (_18275_, _18274_, _02790_);
  or (_18276_, _18275_, _02785_);
  or (_18277_, _18276_, _18272_);
  and (_18278_, _18277_, _18239_);
  or (_18279_, _18278_, _03861_);
  or (_18280_, _18255_, _03860_);
  and (_18281_, _18280_, _18279_);
  or (_18283_, _18281_, _03850_);
  and (_18284_, _06113_, _04679_);
  or (_18285_, _18253_, _06726_);
  or (_18286_, _18285_, _18284_);
  and (_18287_, _18286_, _02970_);
  and (_18288_, _18287_, _18283_);
  or (_18289_, _18288_, _18234_);
  and (_18290_, _18289_, _05261_);
  or (_18291_, _18290_, _18231_);
  and (_18292_, _18291_, _03882_);
  or (_18294_, _10613_, _08596_);
  and (_18295_, _18229_, _02991_);
  and (_18296_, _18295_, _18294_);
  or (_18297_, _10610_, _08596_);
  and (_18298_, _18229_, _03107_);
  and (_18299_, _18298_, _18297_);
  or (_18300_, _10614_, _08596_);
  and (_18301_, _18229_, _02977_);
  and (_18302_, _18301_, _18300_);
  or (_18303_, _18302_, _18299_);
  or (_18305_, _18303_, _18296_);
  or (_18306_, _18305_, _18292_);
  and (_18307_, _18306_, _06161_);
  or (_18308_, _18253_, _04988_);
  and (_18309_, _18245_, _03094_);
  and (_18310_, _18309_, _18308_);
  or (_18311_, _18310_, _18307_);
  and (_18312_, _18311_, _03100_);
  or (_18313_, _18228_, _04988_);
  and (_18314_, _18229_, _02994_);
  and (_18316_, _18314_, _18313_);
  or (_18317_, _18244_, _04988_);
  and (_18318_, _18229_, _03099_);
  and (_18319_, _18318_, _18317_);
  or (_18320_, _18319_, _03133_);
  or (_18321_, _18320_, _18316_);
  or (_18322_, _18321_, _18312_);
  or (_18323_, _18242_, _03138_);
  and (_18324_, _18323_, _03142_);
  and (_18325_, _18324_, _18322_);
  and (_18327_, _18268_, _02778_);
  or (_18328_, _18327_, _02852_);
  or (_18329_, _18328_, _18325_);
  or (_18330_, _18253_, _02853_);
  or (_18331_, _18330_, _18240_);
  and (_18332_, _18331_, _34446_);
  and (_18333_, _18332_, _18329_);
  or (_35625_[1], _18333_, _18226_);
  not (_18334_, \oc8051_golden_model_1.P2 [2]);
  nor (_18335_, _34446_, _18334_);
  or (_18337_, _18335_, rst);
  nor (_18338_, _04679_, _18334_);
  and (_18339_, _10942_, _04679_);
  or (_18340_, _18339_, _18338_);
  and (_18341_, _18340_, _03107_);
  nor (_18342_, _08596_, _04413_);
  or (_18343_, _18342_, _18338_);
  or (_18344_, _18343_, _03860_);
  nor (_18345_, _05278_, _18334_);
  and (_18346_, _10818_, _05278_);
  or (_18348_, _18346_, _18345_);
  or (_18349_, _18348_, _02927_);
  and (_18350_, _18349_, _06189_);
  nor (_18351_, _10824_, _08596_);
  or (_18352_, _18351_, _18338_);
  or (_18353_, _18352_, _06162_);
  and (_18354_, _04679_, \oc8051_golden_model_1.ACC [2]);
  or (_18355_, _18354_, _18338_);
  and (_18356_, _18355_, _02837_);
  nor (_18357_, _02837_, _18334_);
  or (_18359_, _18357_, _02932_);
  or (_18360_, _18359_, _18356_);
  and (_18361_, _18360_, _02939_);
  and (_18362_, _18361_, _18353_);
  and (_18363_, _10815_, _05278_);
  or (_18364_, _18363_, _18345_);
  and (_18365_, _18364_, _02799_);
  and (_18366_, _18343_, _02930_);
  or (_18367_, _18366_, _02928_);
  or (_18368_, _18367_, _18365_);
  or (_18370_, _18368_, _18362_);
  or (_18371_, _18355_, _02943_);
  and (_18372_, _18371_, _18370_);
  or (_18373_, _18372_, _02796_);
  and (_18374_, _18373_, _18350_);
  or (_18375_, _18345_, _10814_);
  and (_18376_, _18375_, _02790_);
  and (_18377_, _18376_, _18364_);
  or (_18378_, _18377_, _18374_);
  and (_18379_, _18378_, _02966_);
  and (_18381_, _16860_, _05278_);
  or (_18382_, _18381_, _18345_);
  and (_18383_, _18382_, _02785_);
  or (_18384_, _18383_, _03861_);
  or (_18385_, _18384_, _18379_);
  and (_18386_, _18385_, _18344_);
  or (_18387_, _18386_, _03850_);
  and (_18388_, _06117_, _04679_);
  or (_18389_, _18338_, _06726_);
  or (_18390_, _18389_, _18388_);
  and (_18392_, _18390_, _02970_);
  and (_18393_, _18392_, _18387_);
  nor (_18394_, _10922_, _08596_);
  or (_18395_, _18394_, _18338_);
  and (_18396_, _18395_, _02524_);
  or (_18397_, _18396_, _02974_);
  or (_18398_, _18397_, _18393_);
  and (_18399_, _04679_, _05690_);
  or (_18400_, _18399_, _18338_);
  or (_18401_, _18400_, _05261_);
  and (_18403_, _18401_, _18398_);
  or (_18404_, _18403_, _02977_);
  and (_18405_, _10936_, _04679_);
  or (_18406_, _18338_, _07092_);
  or (_18407_, _18406_, _18405_);
  and (_18408_, _18407_, _07104_);
  and (_18409_, _18408_, _18404_);
  or (_18410_, _18409_, _18341_);
  and (_18411_, _18410_, _03095_);
  or (_18412_, _18338_, _05086_);
  and (_18414_, _18355_, _03094_);
  and (_18415_, _18400_, _02991_);
  or (_18416_, _18415_, _18414_);
  and (_18417_, _18416_, _18412_);
  or (_18418_, _18417_, _02994_);
  or (_18419_, _18418_, _18411_);
  nor (_18420_, _10935_, _08596_);
  or (_18421_, _18338_, _07120_);
  or (_18422_, _18421_, _18420_);
  and (_18423_, _18422_, _07118_);
  and (_18425_, _18423_, _18419_);
  nor (_18426_, _10941_, _08596_);
  or (_18427_, _18426_, _18338_);
  and (_18428_, _18427_, _03099_);
  or (_18429_, _18428_, _03133_);
  or (_18430_, _18429_, _18425_);
  or (_18431_, _18352_, _03138_);
  and (_18432_, _18431_, _03142_);
  and (_18433_, _18432_, _18430_);
  and (_18434_, _18348_, _02778_);
  or (_18436_, _18434_, _02852_);
  or (_18437_, _18436_, _18433_);
  and (_18438_, _10988_, _04679_);
  or (_18439_, _18338_, _02853_);
  or (_18440_, _18439_, _18438_);
  and (_18441_, _18440_, _34446_);
  and (_18442_, _18441_, _18437_);
  or (_35625_[2], _18442_, _18337_);
  nor (_18443_, \oc8051_golden_model_1.P2 [3], rst);
  nor (_18444_, _18443_, _04509_);
  and (_18446_, _08596_, \oc8051_golden_model_1.P2 [3]);
  and (_18447_, _11134_, _04679_);
  or (_18448_, _18447_, _18446_);
  and (_18449_, _18448_, _03107_);
  nor (_18450_, _08596_, _04226_);
  or (_18451_, _18450_, _18446_);
  or (_18452_, _18451_, _03860_);
  and (_18453_, _16935_, _05278_);
  not (_18454_, _05278_);
  and (_18455_, _18454_, \oc8051_golden_model_1.P2 [3]);
  or (_18457_, _18455_, _02966_);
  or (_18458_, _18457_, _18453_);
  nor (_18459_, _11014_, _08596_);
  or (_18460_, _18459_, _18446_);
  or (_18461_, _18460_, _06162_);
  and (_18462_, _04679_, \oc8051_golden_model_1.ACC [3]);
  or (_18463_, _18462_, _18446_);
  and (_18464_, _18463_, _02837_);
  and (_18465_, _09167_, \oc8051_golden_model_1.P2 [3]);
  or (_18466_, _18465_, _02932_);
  or (_18468_, _18466_, _18464_);
  and (_18469_, _18468_, _02939_);
  and (_18470_, _18469_, _18461_);
  and (_18471_, _18451_, _02930_);
  and (_18472_, _11011_, _05278_);
  or (_18473_, _18472_, _18455_);
  and (_18474_, _18473_, _02799_);
  or (_18475_, _18474_, _18471_);
  or (_18476_, _18475_, _02928_);
  or (_18477_, _18476_, _18470_);
  or (_18479_, _18463_, _02943_);
  and (_18480_, _18479_, _18477_);
  or (_18481_, _18480_, _02796_);
  and (_18482_, _11009_, _05278_);
  or (_18483_, _18482_, _18455_);
  or (_18484_, _18483_, _02927_);
  and (_18485_, _18484_, _06189_);
  and (_18486_, _18485_, _18481_);
  or (_18487_, _18455_, _11040_);
  and (_18488_, _18473_, _02790_);
  and (_18490_, _18488_, _18487_);
  or (_18491_, _18490_, _02785_);
  or (_18492_, _18491_, _18486_);
  and (_18493_, _18492_, _18458_);
  or (_18494_, _18493_, _03861_);
  and (_18495_, _18494_, _18452_);
  or (_18496_, _18495_, _03850_);
  and (_18497_, _06116_, _04679_);
  or (_18498_, _18446_, _06726_);
  or (_18499_, _18498_, _18497_);
  and (_18501_, _18499_, _02970_);
  and (_18502_, _18501_, _18496_);
  nor (_18503_, _11114_, _08596_);
  or (_18504_, _18503_, _18446_);
  and (_18505_, _18504_, _02524_);
  or (_18506_, _18505_, _02974_);
  or (_18507_, _18506_, _18502_);
  and (_18508_, _04679_, _05616_);
  or (_18509_, _18508_, _18446_);
  or (_18510_, _18509_, _05261_);
  and (_18512_, _18510_, _18507_);
  or (_18513_, _18512_, _02977_);
  and (_18514_, _11128_, _04679_);
  or (_18515_, _18446_, _07092_);
  or (_18516_, _18515_, _18514_);
  and (_18517_, _18516_, _07104_);
  and (_18518_, _18517_, _18513_);
  or (_18519_, _18518_, _18449_);
  and (_18520_, _18519_, _03095_);
  or (_18521_, _18446_, _04939_);
  and (_18523_, _18463_, _03094_);
  and (_18524_, _18509_, _02991_);
  or (_18525_, _18524_, _18523_);
  and (_18526_, _18525_, _18521_);
  or (_18527_, _18526_, _02994_);
  or (_18528_, _18527_, _18520_);
  nor (_18529_, _11127_, _08596_);
  or (_18530_, _18446_, _07120_);
  or (_18531_, _18530_, _18529_);
  and (_18532_, _18531_, _07118_);
  and (_18534_, _18532_, _18528_);
  nor (_18535_, _11133_, _08596_);
  or (_18536_, _18535_, _18446_);
  and (_18537_, _18536_, _03099_);
  or (_18538_, _18537_, _03133_);
  or (_18539_, _18538_, _18534_);
  or (_18540_, _18460_, _03138_);
  and (_18541_, _18540_, _03142_);
  and (_18542_, _18541_, _18539_);
  and (_18543_, _18483_, _02778_);
  or (_18545_, _18543_, _02852_);
  or (_18546_, _18545_, _18542_);
  and (_18547_, _11185_, _04679_);
  or (_18548_, _18446_, _02853_);
  or (_18549_, _18548_, _18547_);
  and (_18550_, _18549_, _34446_);
  and (_18551_, _18550_, _18546_);
  or (_35625_[3], _18551_, _18444_);
  nor (_18552_, \oc8051_golden_model_1.P2 [4], rst);
  nor (_18553_, _18552_, _04509_);
  and (_18555_, _08596_, \oc8051_golden_model_1.P2 [4]);
  and (_18556_, _11333_, _04679_);
  or (_18557_, _18556_, _18555_);
  and (_18558_, _18557_, _03107_);
  nor (_18559_, _05143_, _08596_);
  or (_18560_, _18559_, _18555_);
  or (_18561_, _18560_, _03860_);
  and (_18562_, _18454_, \oc8051_golden_model_1.P2 [4]);
  and (_18563_, _11224_, _05278_);
  or (_18564_, _18563_, _18562_);
  or (_18566_, _18562_, _11239_);
  and (_18567_, _18566_, _02790_);
  and (_18568_, _18567_, _18564_);
  nor (_18569_, _11207_, _08596_);
  or (_18570_, _18569_, _18555_);
  or (_18571_, _18570_, _06162_);
  and (_18572_, _04679_, \oc8051_golden_model_1.ACC [4]);
  or (_18573_, _18572_, _18555_);
  and (_18574_, _18573_, _02837_);
  and (_18575_, _09167_, \oc8051_golden_model_1.P2 [4]);
  or (_18577_, _18575_, _02932_);
  or (_18578_, _18577_, _18574_);
  and (_18579_, _18578_, _02939_);
  and (_18580_, _18579_, _18571_);
  and (_18581_, _18560_, _02930_);
  and (_18582_, _18564_, _02799_);
  or (_18583_, _18582_, _18581_);
  or (_18584_, _18583_, _02928_);
  or (_18585_, _18584_, _18580_);
  or (_18586_, _18573_, _02943_);
  and (_18588_, _18586_, _18585_);
  or (_18589_, _18588_, _02796_);
  and (_18590_, _11203_, _05278_);
  or (_18591_, _18590_, _18562_);
  or (_18592_, _18591_, _02927_);
  and (_18593_, _18592_, _06189_);
  and (_18594_, _18593_, _18589_);
  or (_18595_, _18594_, _18568_);
  and (_18596_, _18595_, _02966_);
  and (_18597_, _17080_, _05278_);
  or (_18599_, _18597_, _18562_);
  and (_18600_, _18599_, _02785_);
  or (_18601_, _18600_, _03861_);
  or (_18602_, _18601_, _18596_);
  and (_18603_, _18602_, _18561_);
  or (_18604_, _18603_, _03850_);
  and (_18605_, _06121_, _04679_);
  or (_18606_, _18555_, _06726_);
  or (_18607_, _18606_, _18605_);
  and (_18608_, _18607_, _02970_);
  and (_18610_, _18608_, _18604_);
  nor (_18611_, _11313_, _08596_);
  or (_18612_, _18611_, _18555_);
  and (_18613_, _18612_, _02524_);
  or (_18614_, _18613_, _02974_);
  or (_18615_, _18614_, _18610_);
  and (_18616_, _05629_, _04679_);
  or (_18617_, _18616_, _18555_);
  or (_18618_, _18617_, _05261_);
  and (_18619_, _18618_, _18615_);
  or (_18621_, _18619_, _02977_);
  and (_18622_, _11327_, _04679_);
  or (_18623_, _18555_, _07092_);
  or (_18624_, _18623_, _18622_);
  and (_18625_, _18624_, _07104_);
  and (_18626_, _18625_, _18621_);
  or (_18627_, _18626_, _18558_);
  and (_18628_, _18627_, _03095_);
  or (_18629_, _18555_, _05190_);
  and (_18630_, _18573_, _03094_);
  and (_18632_, _18617_, _02991_);
  or (_18633_, _18632_, _18630_);
  and (_18634_, _18633_, _18629_);
  or (_18635_, _18634_, _02994_);
  or (_18636_, _18635_, _18628_);
  nor (_18637_, _11326_, _08596_);
  or (_18638_, _18555_, _07120_);
  or (_18639_, _18638_, _18637_);
  and (_18640_, _18639_, _07118_);
  and (_18641_, _18640_, _18636_);
  nor (_18643_, _11332_, _08596_);
  or (_18644_, _18643_, _18555_);
  and (_18645_, _18644_, _03099_);
  or (_18646_, _18645_, _03133_);
  or (_18647_, _18646_, _18641_);
  or (_18648_, _18570_, _03138_);
  and (_18649_, _18648_, _03142_);
  and (_18650_, _18649_, _18647_);
  and (_18651_, _18591_, _02778_);
  or (_18652_, _18651_, _02852_);
  or (_18654_, _18652_, _18650_);
  and (_18655_, _11383_, _04679_);
  or (_18656_, _18555_, _02853_);
  or (_18657_, _18656_, _18655_);
  and (_18658_, _18657_, _34446_);
  and (_18659_, _18658_, _18654_);
  or (_35625_[4], _18659_, _18553_);
  nor (_18660_, \oc8051_golden_model_1.P2 [5], rst);
  nor (_18661_, _18660_, _04509_);
  and (_18662_, _08596_, \oc8051_golden_model_1.P2 [5]);
  and (_18664_, _11531_, _04679_);
  or (_18665_, _18664_, _18662_);
  and (_18666_, _18665_, _03107_);
  nor (_18667_, _11408_, _08596_);
  or (_18668_, _18667_, _18662_);
  or (_18669_, _18668_, _06162_);
  and (_18670_, _04679_, \oc8051_golden_model_1.ACC [5]);
  or (_18671_, _18670_, _18662_);
  and (_18672_, _18671_, _02837_);
  and (_18673_, _09167_, \oc8051_golden_model_1.P2 [5]);
  or (_18675_, _18673_, _02932_);
  or (_18676_, _18675_, _18672_);
  and (_18677_, _18676_, _02939_);
  and (_18678_, _18677_, _18669_);
  nor (_18679_, _04839_, _08596_);
  or (_18680_, _18679_, _18662_);
  and (_18681_, _18680_, _02930_);
  and (_18682_, _18454_, \oc8051_golden_model_1.P2 [5]);
  and (_18683_, _11422_, _05278_);
  or (_18684_, _18683_, _18682_);
  and (_18686_, _18684_, _02799_);
  or (_18687_, _18686_, _18681_);
  or (_18688_, _18687_, _02928_);
  or (_18689_, _18688_, _18678_);
  or (_18690_, _18671_, _02943_);
  and (_18691_, _18690_, _18689_);
  or (_18692_, _18691_, _02796_);
  and (_18693_, _11405_, _05278_);
  or (_18694_, _18693_, _18682_);
  or (_18695_, _18694_, _02927_);
  and (_18697_, _18695_, _06189_);
  and (_18698_, _18697_, _18692_);
  and (_18699_, _11438_, _05278_);
  or (_18700_, _18699_, _18682_);
  and (_18701_, _18700_, _02790_);
  or (_18702_, _18701_, _18698_);
  and (_18703_, _18702_, _02966_);
  and (_18704_, _17189_, _05278_);
  or (_18705_, _18704_, _18682_);
  and (_18706_, _18705_, _02785_);
  or (_18708_, _18706_, _03861_);
  or (_18709_, _18708_, _18703_);
  or (_18710_, _18680_, _03860_);
  and (_18711_, _18710_, _18709_);
  or (_18712_, _18711_, _03850_);
  and (_18713_, _06120_, _04679_);
  or (_18714_, _18662_, _06726_);
  or (_18715_, _18714_, _18713_);
  and (_18716_, _18715_, _02970_);
  and (_18717_, _18716_, _18712_);
  nor (_18719_, _11511_, _08596_);
  or (_18720_, _18719_, _18662_);
  and (_18721_, _18720_, _02524_);
  or (_18722_, _18721_, _02974_);
  or (_18723_, _18722_, _18717_);
  and (_18724_, _05633_, _04679_);
  or (_18725_, _18724_, _18662_);
  or (_18726_, _18725_, _05261_);
  and (_18727_, _18726_, _18723_);
  or (_18728_, _18727_, _02977_);
  and (_18730_, _11525_, _04679_);
  or (_18731_, _18662_, _07092_);
  or (_18732_, _18731_, _18730_);
  and (_18733_, _18732_, _07104_);
  and (_18734_, _18733_, _18728_);
  or (_18735_, _18734_, _18666_);
  and (_18736_, _18735_, _03095_);
  or (_18737_, _18662_, _04890_);
  and (_18738_, _18671_, _03094_);
  and (_18739_, _18725_, _02991_);
  or (_18741_, _18739_, _18738_);
  and (_18742_, _18741_, _18737_);
  or (_18743_, _18742_, _02994_);
  or (_18744_, _18743_, _18736_);
  nor (_18745_, _11524_, _08596_);
  or (_18746_, _18662_, _07120_);
  or (_18747_, _18746_, _18745_);
  and (_18748_, _18747_, _07118_);
  and (_18749_, _18748_, _18744_);
  nor (_18750_, _11530_, _08596_);
  or (_18752_, _18750_, _18662_);
  and (_18753_, _18752_, _03099_);
  or (_18754_, _18753_, _03133_);
  or (_18755_, _18754_, _18749_);
  or (_18756_, _18668_, _03138_);
  and (_18757_, _18756_, _03142_);
  and (_18758_, _18757_, _18755_);
  and (_18759_, _18694_, _02778_);
  or (_18760_, _18759_, _02852_);
  or (_18761_, _18760_, _18758_);
  and (_18763_, _11580_, _04679_);
  or (_18764_, _18662_, _02853_);
  or (_18765_, _18764_, _18763_);
  and (_18766_, _18765_, _34446_);
  and (_18767_, _18766_, _18761_);
  or (_35625_[5], _18767_, _18661_);
  not (_18768_, \oc8051_golden_model_1.P2 [6]);
  nor (_18769_, _34446_, _18768_);
  or (_18770_, _18769_, rst);
  nor (_18771_, _04679_, _18768_);
  and (_18773_, _11601_, _04679_);
  or (_18774_, _18773_, _18771_);
  and (_18775_, _18774_, _03107_);
  nor (_18776_, _04735_, _08596_);
  or (_18777_, _18776_, _18771_);
  or (_18778_, _18777_, _03860_);
  nor (_18779_, _11610_, _08596_);
  or (_18780_, _18779_, _18771_);
  or (_18781_, _18780_, _06162_);
  and (_18782_, _04679_, \oc8051_golden_model_1.ACC [6]);
  or (_18784_, _18782_, _18771_);
  and (_18785_, _18784_, _02837_);
  nor (_18786_, _02837_, _18768_);
  or (_18787_, _18786_, _02932_);
  or (_18788_, _18787_, _18785_);
  and (_18789_, _18788_, _02939_);
  and (_18790_, _18789_, _18781_);
  and (_18791_, _18777_, _02930_);
  nor (_18792_, _05278_, _18768_);
  and (_18793_, _11604_, _05278_);
  or (_18795_, _18793_, _18792_);
  and (_18796_, _18795_, _02799_);
  or (_18797_, _18796_, _18791_);
  or (_18798_, _18797_, _02928_);
  or (_18799_, _18798_, _18790_);
  or (_18800_, _18784_, _02943_);
  and (_18801_, _18800_, _18799_);
  or (_18802_, _18801_, _02796_);
  and (_18803_, _11633_, _05278_);
  or (_18804_, _18803_, _18792_);
  or (_18806_, _18804_, _02927_);
  and (_18807_, _18806_, _06189_);
  and (_18808_, _18807_, _18802_);
  and (_18809_, _11605_, _05278_);
  or (_18810_, _18809_, _18792_);
  and (_18811_, _18810_, _02790_);
  or (_18812_, _18811_, _18808_);
  and (_18813_, _18812_, _02966_);
  and (_18814_, _17300_, _05278_);
  or (_18815_, _18814_, _18792_);
  and (_18817_, _18815_, _02785_);
  or (_18818_, _18817_, _03861_);
  or (_18819_, _18818_, _18813_);
  and (_18820_, _18819_, _18778_);
  or (_18821_, _18820_, _03850_);
  and (_18822_, _05798_, _04679_);
  or (_18823_, _18771_, _06726_);
  or (_18824_, _18823_, _18822_);
  and (_18825_, _18824_, _02970_);
  and (_18826_, _18825_, _18821_);
  nor (_18828_, _11711_, _08596_);
  or (_18829_, _18828_, _18771_);
  and (_18830_, _18829_, _02524_);
  or (_18831_, _18830_, _02974_);
  or (_18832_, _18831_, _18826_);
  and (_18833_, _11718_, _04679_);
  or (_18834_, _18833_, _18771_);
  or (_18835_, _18834_, _05261_);
  and (_18836_, _18835_, _18832_);
  or (_18837_, _18836_, _02977_);
  and (_18839_, _11728_, _04679_);
  or (_18840_, _18771_, _07092_);
  or (_18841_, _18840_, _18839_);
  and (_18842_, _18841_, _07104_);
  and (_18843_, _18842_, _18837_);
  or (_18844_, _18843_, _18775_);
  and (_18845_, _18844_, _03095_);
  or (_18846_, _18771_, _04784_);
  and (_18847_, _18784_, _03094_);
  and (_18848_, _18834_, _02991_);
  or (_18850_, _18848_, _18847_);
  and (_18851_, _18850_, _18846_);
  or (_18852_, _18851_, _02994_);
  or (_18853_, _18852_, _18845_);
  nor (_18854_, _11726_, _08596_);
  or (_18855_, _18771_, _07120_);
  or (_18856_, _18855_, _18854_);
  and (_18857_, _18856_, _07118_);
  and (_18858_, _18857_, _18853_);
  nor (_18859_, _11600_, _08596_);
  or (_18861_, _18859_, _18771_);
  and (_18862_, _18861_, _03099_);
  or (_18863_, _18862_, _03133_);
  or (_18864_, _18863_, _18858_);
  or (_18865_, _18780_, _03138_);
  and (_18866_, _18865_, _03142_);
  and (_18867_, _18866_, _18864_);
  and (_18868_, _18804_, _02778_);
  or (_18869_, _18868_, _02852_);
  or (_18870_, _18869_, _18867_);
  and (_18872_, _11778_, _04679_);
  or (_18873_, _18771_, _02853_);
  or (_18874_, _18873_, _18872_);
  and (_18875_, _18874_, _34446_);
  and (_18876_, _18875_, _18870_);
  or (_35625_[6], _18876_, _18770_);
  not (_18877_, \oc8051_golden_model_1.P3 [0]);
  nor (_18878_, _34446_, _18877_);
  or (_18879_, _18878_, rst);
  nor (_18880_, _04681_, _18877_);
  and (_18882_, _10546_, _04681_);
  or (_18883_, _18882_, _18880_);
  and (_18884_, _18883_, _03107_);
  and (_18885_, _04681_, _03805_);
  or (_18886_, _18885_, _18880_);
  or (_18887_, _18886_, _03860_);
  nor (_18888_, _05280_, _18877_);
  and (_18889_, _10441_, _05280_);
  or (_18890_, _18889_, _18888_);
  and (_18891_, _18890_, _02799_);
  nor (_18893_, _05036_, _08690_);
  or (_18894_, _18893_, _18880_);
  or (_18895_, _18894_, _06162_);
  and (_18896_, _04681_, \oc8051_golden_model_1.ACC [0]);
  or (_18897_, _18896_, _18880_);
  and (_18898_, _18897_, _02837_);
  nor (_18899_, _02837_, _18877_);
  or (_18900_, _18899_, _02932_);
  or (_18901_, _18900_, _18898_);
  and (_18902_, _18901_, _02939_);
  and (_18904_, _18902_, _18895_);
  and (_18905_, _18886_, _02930_);
  or (_18906_, _18905_, _02928_);
  or (_18907_, _18906_, _18904_);
  or (_18908_, _18907_, _18891_);
  or (_18909_, _18897_, _02943_);
  and (_18910_, _18909_, _02927_);
  and (_18911_, _18910_, _18908_);
  and (_18912_, _18880_, _02796_);
  or (_18913_, _18912_, _02790_);
  or (_18915_, _18913_, _18911_);
  or (_18916_, _18894_, _06189_);
  and (_18917_, _18916_, _02966_);
  and (_18918_, _18917_, _18915_);
  and (_18919_, _16640_, _05280_);
  or (_18920_, _18919_, _18888_);
  and (_18921_, _18920_, _02785_);
  or (_18922_, _18921_, _03861_);
  or (_18923_, _18922_, _18918_);
  and (_18924_, _18923_, _18887_);
  or (_18926_, _18924_, _03850_);
  and (_18927_, _06114_, _04681_);
  or (_18928_, _18880_, _06726_);
  or (_18929_, _18928_, _18927_);
  and (_18930_, _18929_, _02970_);
  and (_18931_, _18930_, _18926_);
  nor (_18932_, _10530_, _08690_);
  or (_18933_, _18932_, _18880_);
  and (_18934_, _18933_, _02524_);
  or (_18935_, _18934_, _02974_);
  or (_18937_, _18935_, _18931_);
  and (_18938_, _04681_, _05647_);
  or (_18939_, _18938_, _18880_);
  or (_18940_, _18939_, _05261_);
  and (_18941_, _18940_, _18937_);
  or (_18942_, _18941_, _02977_);
  and (_18943_, _10427_, _04681_);
  or (_18944_, _18880_, _07092_);
  or (_18945_, _18944_, _18943_);
  and (_18946_, _18945_, _07104_);
  and (_18948_, _18946_, _18942_);
  or (_18949_, _18948_, _18884_);
  and (_18950_, _18949_, _03095_);
  nand (_18951_, _18939_, _02991_);
  nor (_18952_, _18951_, _18893_);
  or (_18953_, _18880_, _05036_);
  and (_18954_, _18897_, _03094_);
  and (_18955_, _18954_, _18953_);
  or (_18956_, _18955_, _02994_);
  or (_18957_, _18956_, _18952_);
  or (_18959_, _18957_, _18950_);
  nor (_18960_, _10425_, _08690_);
  or (_18961_, _18880_, _07120_);
  or (_18962_, _18961_, _18960_);
  and (_18963_, _18962_, _07118_);
  and (_18964_, _18963_, _18959_);
  nor (_18965_, _10423_, _08690_);
  or (_18966_, _18965_, _18880_);
  and (_18967_, _18966_, _03099_);
  or (_18968_, _18967_, _03133_);
  or (_18970_, _18968_, _18964_);
  or (_18971_, _18894_, _03138_);
  and (_18972_, _18971_, _03142_);
  and (_18973_, _18972_, _18970_);
  and (_18974_, _18880_, _02778_);
  or (_18975_, _18974_, _02852_);
  or (_18976_, _18975_, _18973_);
  or (_18977_, _18894_, _02853_);
  and (_18978_, _18977_, _34446_);
  and (_18979_, _18978_, _18976_);
  or (_35627_[0], _18979_, _18879_);
  not (_18981_, \oc8051_golden_model_1.P3 [1]);
  nor (_18982_, _34446_, _18981_);
  or (_18983_, _18982_, rst);
  nand (_18984_, _04681_, _03660_);
  or (_18985_, _04681_, \oc8051_golden_model_1.P3 [1]);
  and (_18986_, _18985_, _02974_);
  and (_18987_, _18986_, _18984_);
  nand (_18988_, _10719_, _04681_);
  and (_18989_, _18985_, _02524_);
  and (_18991_, _18989_, _18988_);
  and (_18992_, _16710_, _05280_);
  nor (_18993_, _05280_, _18981_);
  or (_18994_, _18993_, _02966_);
  or (_18995_, _18994_, _18992_);
  and (_18996_, _10622_, _04681_);
  not (_18997_, _18996_);
  and (_18998_, _18997_, _18985_);
  or (_18999_, _18998_, _06162_);
  nand (_19000_, _04681_, _02477_);
  and (_19002_, _19000_, _18985_);
  and (_19003_, _19002_, _02837_);
  nor (_19004_, _02837_, _18981_);
  or (_19005_, _19004_, _02932_);
  or (_19006_, _19005_, _19003_);
  and (_19007_, _19006_, _02939_);
  and (_19008_, _19007_, _18999_);
  nor (_19009_, _04681_, _18981_);
  nor (_19010_, _08690_, _03989_);
  or (_19011_, _19010_, _19009_);
  and (_19013_, _19011_, _02930_);
  and (_19014_, _10617_, _05280_);
  or (_19015_, _19014_, _18993_);
  and (_19016_, _19015_, _02799_);
  or (_19017_, _19016_, _19013_);
  or (_19018_, _19017_, _02928_);
  or (_19019_, _19018_, _19008_);
  or (_19020_, _19002_, _02943_);
  and (_19021_, _19020_, _19019_);
  or (_19022_, _19021_, _02796_);
  and (_19024_, _10620_, _05280_);
  or (_19025_, _19024_, _18993_);
  or (_19026_, _19025_, _02927_);
  and (_19027_, _19026_, _06189_);
  and (_19028_, _19027_, _19022_);
  and (_19029_, _19014_, _10616_);
  or (_19030_, _19029_, _18993_);
  and (_19031_, _19030_, _02790_);
  or (_19032_, _19031_, _02785_);
  or (_19033_, _19032_, _19028_);
  and (_19035_, _19033_, _18995_);
  or (_19036_, _19035_, _03861_);
  or (_19037_, _19011_, _03860_);
  and (_19038_, _19037_, _19036_);
  or (_19039_, _19038_, _03850_);
  and (_19040_, _06113_, _04681_);
  or (_19041_, _19009_, _06726_);
  or (_19042_, _19041_, _19040_);
  and (_19043_, _19042_, _02970_);
  and (_19044_, _19043_, _19039_);
  or (_19046_, _19044_, _18991_);
  and (_19047_, _19046_, _05261_);
  or (_19048_, _19047_, _18987_);
  and (_19049_, _19048_, _03882_);
  or (_19050_, _10613_, _08690_);
  and (_19051_, _18985_, _02991_);
  and (_19052_, _19051_, _19050_);
  or (_19053_, _10610_, _08690_);
  and (_19054_, _18985_, _03107_);
  and (_19055_, _19054_, _19053_);
  or (_19057_, _10614_, _08690_);
  and (_19058_, _18985_, _02977_);
  and (_19059_, _19058_, _19057_);
  or (_19060_, _19059_, _19055_);
  or (_19061_, _19060_, _19052_);
  or (_19062_, _19061_, _19049_);
  and (_19063_, _19062_, _06161_);
  or (_19064_, _19009_, _04988_);
  and (_19065_, _19002_, _03094_);
  and (_19066_, _19065_, _19064_);
  or (_19068_, _19066_, _19063_);
  and (_19069_, _19068_, _03100_);
  or (_19070_, _18984_, _04988_);
  and (_19071_, _18985_, _02994_);
  and (_19072_, _19071_, _19070_);
  or (_19073_, _19000_, _04988_);
  and (_19074_, _18985_, _03099_);
  and (_19075_, _19074_, _19073_);
  or (_19076_, _19075_, _03133_);
  or (_19077_, _19076_, _19072_);
  or (_19079_, _19077_, _19069_);
  or (_19080_, _18998_, _03138_);
  and (_19081_, _19080_, _03142_);
  and (_19082_, _19081_, _19079_);
  and (_19083_, _19025_, _02778_);
  or (_19084_, _19083_, _02852_);
  or (_19085_, _19084_, _19082_);
  or (_19086_, _19009_, _02853_);
  or (_19087_, _19086_, _18996_);
  and (_19088_, _19087_, _34446_);
  and (_19090_, _19088_, _19085_);
  or (_35627_[1], _19090_, _18983_);
  not (_19091_, \oc8051_golden_model_1.P3 [2]);
  nor (_19092_, _34446_, _19091_);
  or (_19093_, _19092_, rst);
  nor (_19094_, _04681_, _19091_);
  and (_19095_, _10942_, _04681_);
  or (_19096_, _19095_, _19094_);
  and (_19097_, _19096_, _03107_);
  nor (_19098_, _08690_, _04413_);
  or (_19100_, _19098_, _19094_);
  or (_19101_, _19100_, _03860_);
  nor (_19102_, _10824_, _08690_);
  or (_19103_, _19102_, _19094_);
  or (_19104_, _19103_, _06162_);
  and (_19105_, _04681_, \oc8051_golden_model_1.ACC [2]);
  or (_19106_, _19105_, _19094_);
  and (_19107_, _19106_, _02837_);
  nor (_19108_, _02837_, _19091_);
  or (_19109_, _19108_, _02932_);
  or (_19111_, _19109_, _19107_);
  and (_19112_, _19111_, _02939_);
  and (_19113_, _19112_, _19104_);
  and (_19114_, _19100_, _02930_);
  nor (_19115_, _05280_, _19091_);
  and (_19116_, _10815_, _05280_);
  or (_19117_, _19116_, _19115_);
  and (_19118_, _19117_, _02799_);
  or (_19119_, _19118_, _19114_);
  or (_19120_, _19119_, _02928_);
  or (_19122_, _19120_, _19113_);
  or (_19123_, _19106_, _02943_);
  and (_19124_, _19123_, _19122_);
  or (_19125_, _19124_, _02796_);
  and (_19126_, _10818_, _05280_);
  or (_19127_, _19126_, _19115_);
  or (_19128_, _19127_, _02927_);
  and (_19129_, _19128_, _06189_);
  and (_19130_, _19129_, _19125_);
  and (_19131_, _19116_, _10814_);
  or (_19133_, _19131_, _19115_);
  and (_19134_, _19133_, _02790_);
  or (_19135_, _19134_, _19130_);
  and (_19136_, _19135_, _02966_);
  and (_19137_, _16860_, _05280_);
  or (_19138_, _19115_, _19137_);
  and (_19139_, _19138_, _02785_);
  or (_19140_, _19139_, _03861_);
  or (_19141_, _19140_, _19136_);
  and (_19142_, _19141_, _19101_);
  or (_19144_, _19142_, _03850_);
  and (_19145_, _06117_, _04681_);
  or (_19146_, _19094_, _06726_);
  or (_19147_, _19146_, _19145_);
  and (_19148_, _19147_, _02970_);
  and (_19149_, _19148_, _19144_);
  nor (_19150_, _10922_, _08690_);
  or (_19151_, _19150_, _19094_);
  and (_19152_, _19151_, _02524_);
  or (_19153_, _19152_, _02974_);
  or (_19155_, _19153_, _19149_);
  and (_19156_, _04681_, _05690_);
  or (_19157_, _19156_, _19094_);
  or (_19158_, _19157_, _05261_);
  and (_19159_, _19158_, _19155_);
  or (_19160_, _19159_, _02977_);
  and (_19161_, _10936_, _04681_);
  or (_19162_, _19094_, _07092_);
  or (_19163_, _19162_, _19161_);
  and (_19164_, _19163_, _07104_);
  and (_19166_, _19164_, _19160_);
  or (_19167_, _19166_, _19097_);
  and (_19168_, _19167_, _03095_);
  or (_19169_, _19094_, _05086_);
  and (_19170_, _19106_, _03094_);
  and (_19171_, _19157_, _02991_);
  or (_19172_, _19171_, _19170_);
  and (_19173_, _19172_, _19169_);
  or (_19174_, _19173_, _02994_);
  or (_19175_, _19174_, _19168_);
  nor (_19177_, _10935_, _08690_);
  or (_19178_, _19094_, _07120_);
  or (_19179_, _19178_, _19177_);
  and (_19180_, _19179_, _07118_);
  and (_19181_, _19180_, _19175_);
  nor (_19182_, _10941_, _08690_);
  or (_19183_, _19182_, _19094_);
  and (_19184_, _19183_, _03099_);
  or (_19185_, _19184_, _03133_);
  or (_19186_, _19185_, _19181_);
  or (_19188_, _19103_, _03138_);
  and (_19189_, _19188_, _03142_);
  and (_19190_, _19189_, _19186_);
  and (_19191_, _19127_, _02778_);
  or (_19192_, _19191_, _02852_);
  or (_19193_, _19192_, _19190_);
  and (_19194_, _10988_, _04681_);
  or (_19195_, _19094_, _02853_);
  or (_19196_, _19195_, _19194_);
  and (_19197_, _19196_, _34446_);
  and (_19199_, _19197_, _19193_);
  or (_35627_[2], _19199_, _19093_);
  nor (_19200_, \oc8051_golden_model_1.P3 [3], rst);
  nor (_19201_, _19200_, _04509_);
  and (_19202_, _08690_, \oc8051_golden_model_1.P3 [3]);
  and (_19203_, _11134_, _04681_);
  or (_19204_, _19203_, _19202_);
  and (_19205_, _19204_, _03107_);
  nor (_19206_, _08690_, _04226_);
  or (_19207_, _19206_, _19202_);
  or (_19209_, _19207_, _03860_);
  and (_19210_, _16935_, _05280_);
  not (_19211_, _05280_);
  and (_19212_, _19211_, \oc8051_golden_model_1.P3 [3]);
  or (_19213_, _19212_, _02966_);
  or (_19214_, _19213_, _19210_);
  nor (_19215_, _11014_, _08690_);
  or (_19216_, _19215_, _19202_);
  or (_19217_, _19216_, _06162_);
  and (_19218_, _04681_, \oc8051_golden_model_1.ACC [3]);
  or (_19220_, _19218_, _19202_);
  and (_19221_, _19220_, _02837_);
  and (_19222_, _09167_, \oc8051_golden_model_1.P3 [3]);
  or (_19223_, _19222_, _02932_);
  or (_19224_, _19223_, _19221_);
  and (_19225_, _19224_, _02939_);
  and (_19226_, _19225_, _19217_);
  and (_19227_, _19207_, _02930_);
  and (_19228_, _11011_, _05280_);
  or (_19229_, _19228_, _19212_);
  and (_19231_, _19229_, _02799_);
  or (_19232_, _19231_, _19227_);
  or (_19233_, _19232_, _02928_);
  or (_19234_, _19233_, _19226_);
  or (_19235_, _19220_, _02943_);
  and (_19236_, _19235_, _19234_);
  or (_19237_, _19236_, _02796_);
  and (_19238_, _11009_, _05280_);
  or (_19239_, _19238_, _19212_);
  or (_19240_, _19239_, _02927_);
  and (_19242_, _19240_, _06189_);
  and (_19243_, _19242_, _19237_);
  or (_19244_, _19212_, _11040_);
  and (_19245_, _19229_, _02790_);
  and (_19246_, _19245_, _19244_);
  or (_19247_, _19246_, _02785_);
  or (_19248_, _19247_, _19243_);
  and (_19249_, _19248_, _19214_);
  or (_19250_, _19249_, _03861_);
  and (_19251_, _19250_, _19209_);
  or (_19253_, _19251_, _03850_);
  and (_19254_, _06116_, _04681_);
  or (_19255_, _19202_, _06726_);
  or (_19256_, _19255_, _19254_);
  and (_19257_, _19256_, _02970_);
  and (_19258_, _19257_, _19253_);
  nor (_19259_, _11114_, _08690_);
  or (_19260_, _19259_, _19202_);
  and (_19261_, _19260_, _02524_);
  or (_19262_, _19261_, _02974_);
  or (_19264_, _19262_, _19258_);
  and (_19265_, _04681_, _05616_);
  or (_19266_, _19265_, _19202_);
  or (_19267_, _19266_, _05261_);
  and (_19268_, _19267_, _19264_);
  or (_19269_, _19268_, _02977_);
  and (_19270_, _11128_, _04681_);
  or (_19271_, _19202_, _07092_);
  or (_19272_, _19271_, _19270_);
  and (_19273_, _19272_, _07104_);
  and (_19275_, _19273_, _19269_);
  or (_19276_, _19275_, _19205_);
  and (_19277_, _19276_, _03095_);
  or (_19278_, _19202_, _04939_);
  and (_19279_, _19220_, _03094_);
  and (_19280_, _19266_, _02991_);
  or (_19281_, _19280_, _19279_);
  and (_19282_, _19281_, _19278_);
  or (_19283_, _19282_, _02994_);
  or (_19284_, _19283_, _19277_);
  nor (_19286_, _11127_, _08690_);
  or (_19287_, _19202_, _07120_);
  or (_19288_, _19287_, _19286_);
  and (_19289_, _19288_, _07118_);
  and (_19290_, _19289_, _19284_);
  nor (_19291_, _11133_, _08690_);
  or (_19292_, _19291_, _19202_);
  and (_19293_, _19292_, _03099_);
  or (_19294_, _19293_, _03133_);
  or (_19295_, _19294_, _19290_);
  or (_19297_, _19216_, _03138_);
  and (_19298_, _19297_, _03142_);
  and (_19299_, _19298_, _19295_);
  and (_19300_, _19239_, _02778_);
  or (_19301_, _19300_, _02852_);
  or (_19302_, _19301_, _19299_);
  and (_19303_, _11185_, _04681_);
  or (_19304_, _19202_, _02853_);
  or (_19305_, _19304_, _19303_);
  and (_19306_, _19305_, _34446_);
  and (_19308_, _19306_, _19302_);
  or (_35627_[3], _19308_, _19201_);
  nor (_19309_, \oc8051_golden_model_1.P3 [4], rst);
  nor (_19310_, _19309_, _04509_);
  and (_19311_, _08690_, \oc8051_golden_model_1.P3 [4]);
  and (_19312_, _11333_, _04681_);
  or (_19313_, _19312_, _19311_);
  and (_19314_, _19313_, _03107_);
  nor (_19315_, _05143_, _08690_);
  or (_19316_, _19315_, _19311_);
  or (_19318_, _19316_, _03860_);
  and (_19319_, _19211_, \oc8051_golden_model_1.P3 [4]);
  and (_19320_, _11224_, _05280_);
  or (_19321_, _19320_, _19319_);
  or (_19322_, _19319_, _11239_);
  and (_19323_, _19322_, _02790_);
  and (_19324_, _19323_, _19321_);
  nor (_19325_, _11207_, _08690_);
  or (_19326_, _19325_, _19311_);
  or (_19327_, _19326_, _06162_);
  and (_19329_, _04681_, \oc8051_golden_model_1.ACC [4]);
  or (_19330_, _19329_, _19311_);
  and (_19331_, _19330_, _02837_);
  and (_19332_, _09167_, \oc8051_golden_model_1.P3 [4]);
  or (_19333_, _19332_, _02932_);
  or (_19334_, _19333_, _19331_);
  and (_19335_, _19334_, _02939_);
  and (_19336_, _19335_, _19327_);
  and (_19337_, _19316_, _02930_);
  and (_19338_, _19321_, _02799_);
  or (_19340_, _19338_, _19337_);
  or (_19341_, _19340_, _02928_);
  or (_19342_, _19341_, _19336_);
  or (_19343_, _19330_, _02943_);
  and (_19344_, _19343_, _19342_);
  or (_19345_, _19344_, _02796_);
  and (_19346_, _11203_, _05280_);
  or (_19347_, _19346_, _19319_);
  or (_19348_, _19347_, _02927_);
  and (_19349_, _19348_, _06189_);
  and (_19351_, _19349_, _19345_);
  or (_19352_, _19351_, _19324_);
  and (_19353_, _19352_, _02966_);
  and (_19354_, _17080_, _05280_);
  or (_19355_, _19354_, _19319_);
  and (_19356_, _19355_, _02785_);
  or (_19357_, _19356_, _03861_);
  or (_19358_, _19357_, _19353_);
  and (_19359_, _19358_, _19318_);
  or (_19360_, _19359_, _03850_);
  and (_19362_, _06121_, _04681_);
  or (_19363_, _19311_, _06726_);
  or (_19364_, _19363_, _19362_);
  and (_19365_, _19364_, _02970_);
  and (_19366_, _19365_, _19360_);
  nor (_19367_, _11313_, _08690_);
  or (_19368_, _19367_, _19311_);
  and (_19369_, _19368_, _02524_);
  or (_19370_, _19369_, _02974_);
  or (_19371_, _19370_, _19366_);
  and (_19373_, _05629_, _04681_);
  or (_19374_, _19373_, _19311_);
  or (_19375_, _19374_, _05261_);
  and (_19376_, _19375_, _19371_);
  or (_19377_, _19376_, _02977_);
  and (_19378_, _11327_, _04681_);
  or (_19379_, _19311_, _07092_);
  or (_19380_, _19379_, _19378_);
  and (_19381_, _19380_, _07104_);
  and (_19382_, _19381_, _19377_);
  or (_19384_, _19382_, _19314_);
  and (_19385_, _19384_, _03095_);
  or (_19386_, _19311_, _05190_);
  and (_19387_, _19330_, _03094_);
  and (_19388_, _19374_, _02991_);
  or (_19389_, _19388_, _19387_);
  and (_19390_, _19389_, _19386_);
  or (_19391_, _19390_, _02994_);
  or (_19392_, _19391_, _19385_);
  nor (_19393_, _11326_, _08690_);
  or (_19395_, _19311_, _07120_);
  or (_19396_, _19395_, _19393_);
  and (_19397_, _19396_, _07118_);
  and (_19398_, _19397_, _19392_);
  nor (_19399_, _11332_, _08690_);
  or (_19400_, _19399_, _19311_);
  and (_19401_, _19400_, _03099_);
  or (_19402_, _19401_, _03133_);
  or (_19403_, _19402_, _19398_);
  or (_19404_, _19326_, _03138_);
  and (_19406_, _19404_, _03142_);
  and (_19407_, _19406_, _19403_);
  and (_19408_, _19347_, _02778_);
  or (_19409_, _19408_, _02852_);
  or (_19410_, _19409_, _19407_);
  and (_19411_, _11383_, _04681_);
  or (_19412_, _19311_, _02853_);
  or (_19413_, _19412_, _19411_);
  and (_19414_, _19413_, _34446_);
  and (_19415_, _19414_, _19410_);
  or (_35627_[4], _19415_, _19310_);
  nor (_19417_, \oc8051_golden_model_1.P3 [5], rst);
  nor (_19418_, _19417_, _04509_);
  and (_19419_, _08690_, \oc8051_golden_model_1.P3 [5]);
  and (_19420_, _11531_, _04681_);
  or (_19421_, _19420_, _19419_);
  and (_19422_, _19421_, _03107_);
  and (_19423_, _19211_, \oc8051_golden_model_1.P3 [5]);
  and (_19424_, _11422_, _05280_);
  or (_19425_, _19424_, _19423_);
  or (_19427_, _19423_, _11437_);
  and (_19428_, _19427_, _02790_);
  and (_19429_, _19428_, _19425_);
  nor (_19430_, _11408_, _08690_);
  or (_19431_, _19430_, _19419_);
  or (_19432_, _19431_, _06162_);
  and (_19433_, _04681_, \oc8051_golden_model_1.ACC [5]);
  or (_19434_, _19433_, _19419_);
  and (_19435_, _19434_, _02837_);
  and (_19436_, _09167_, \oc8051_golden_model_1.P3 [5]);
  or (_19438_, _19436_, _02932_);
  or (_19439_, _19438_, _19435_);
  and (_19440_, _19439_, _02939_);
  and (_19441_, _19440_, _19432_);
  nor (_19442_, _04839_, _08690_);
  or (_19443_, _19442_, _19419_);
  and (_19444_, _19443_, _02930_);
  and (_19445_, _19425_, _02799_);
  or (_19446_, _19445_, _19444_);
  or (_19447_, _19446_, _02928_);
  or (_19449_, _19447_, _19441_);
  or (_19450_, _19434_, _02943_);
  and (_19451_, _19450_, _19449_);
  or (_19452_, _19451_, _02796_);
  and (_19453_, _11405_, _05280_);
  or (_19454_, _19453_, _19423_);
  or (_19455_, _19454_, _02927_);
  and (_19456_, _19455_, _06189_);
  and (_19457_, _19456_, _19452_);
  or (_19458_, _19457_, _19429_);
  and (_19460_, _19458_, _02966_);
  and (_19461_, _17189_, _05280_);
  or (_19462_, _19461_, _19423_);
  and (_19463_, _19462_, _02785_);
  or (_19464_, _19463_, _03861_);
  or (_19465_, _19464_, _19460_);
  or (_19466_, _19443_, _03860_);
  and (_19467_, _19466_, _19465_);
  or (_19468_, _19467_, _03850_);
  and (_19469_, _06120_, _04681_);
  or (_19471_, _19419_, _06726_);
  or (_19472_, _19471_, _19469_);
  and (_19473_, _19472_, _02970_);
  and (_19474_, _19473_, _19468_);
  nor (_19475_, _11511_, _08690_);
  or (_19476_, _19475_, _19419_);
  and (_19477_, _19476_, _02524_);
  or (_19478_, _19477_, _02974_);
  or (_19479_, _19478_, _19474_);
  and (_19480_, _05633_, _04681_);
  or (_19482_, _19480_, _19419_);
  or (_19483_, _19482_, _05261_);
  and (_19484_, _19483_, _19479_);
  or (_19485_, _19484_, _02977_);
  and (_19486_, _11525_, _04681_);
  or (_19487_, _19419_, _07092_);
  or (_19488_, _19487_, _19486_);
  and (_19489_, _19488_, _07104_);
  and (_19490_, _19489_, _19485_);
  or (_19491_, _19490_, _19422_);
  and (_19493_, _19491_, _03095_);
  or (_19494_, _19419_, _04890_);
  and (_19495_, _19434_, _03094_);
  and (_19496_, _19482_, _02991_);
  or (_19497_, _19496_, _19495_);
  and (_19498_, _19497_, _19494_);
  or (_19499_, _19498_, _02994_);
  or (_19500_, _19499_, _19493_);
  nor (_19501_, _11524_, _08690_);
  or (_19502_, _19419_, _07120_);
  or (_19504_, _19502_, _19501_);
  and (_19505_, _19504_, _07118_);
  and (_19506_, _19505_, _19500_);
  nor (_19507_, _11530_, _08690_);
  or (_19508_, _19507_, _19419_);
  and (_19509_, _19508_, _03099_);
  or (_19510_, _19509_, _03133_);
  or (_19511_, _19510_, _19506_);
  or (_19512_, _19431_, _03138_);
  and (_19513_, _19512_, _03142_);
  and (_19515_, _19513_, _19511_);
  and (_19516_, _19454_, _02778_);
  or (_19517_, _19516_, _02852_);
  or (_19518_, _19517_, _19515_);
  and (_19519_, _11580_, _04681_);
  or (_19520_, _19419_, _02853_);
  or (_19521_, _19520_, _19519_);
  and (_19522_, _19521_, _34446_);
  and (_19523_, _19522_, _19518_);
  or (_35627_[5], _19523_, _19418_);
  not (_19525_, \oc8051_golden_model_1.P3 [6]);
  nor (_19526_, _34446_, _19525_);
  or (_19527_, _19526_, rst);
  nor (_19528_, _04681_, _19525_);
  and (_19529_, _11601_, _04681_);
  or (_19530_, _19529_, _19528_);
  and (_19531_, _19530_, _03107_);
  nor (_19532_, _04735_, _08690_);
  or (_19533_, _19532_, _19528_);
  or (_19534_, _19533_, _03860_);
  nor (_19536_, _11610_, _08690_);
  or (_19537_, _19536_, _19528_);
  or (_19538_, _19537_, _06162_);
  and (_19539_, _04681_, \oc8051_golden_model_1.ACC [6]);
  or (_19540_, _19539_, _19528_);
  and (_19541_, _19540_, _02837_);
  nor (_19542_, _02837_, _19525_);
  or (_19543_, _19542_, _02932_);
  or (_19544_, _19543_, _19541_);
  and (_19545_, _19544_, _02939_);
  and (_19547_, _19545_, _19538_);
  and (_19548_, _19533_, _02930_);
  nor (_19549_, _05280_, _19525_);
  and (_19550_, _11604_, _05280_);
  or (_19551_, _19550_, _19549_);
  and (_19552_, _19551_, _02799_);
  or (_19553_, _19552_, _19548_);
  or (_19554_, _19553_, _02928_);
  or (_19555_, _19554_, _19547_);
  or (_19556_, _19540_, _02943_);
  and (_19558_, _19556_, _19555_);
  or (_19559_, _19558_, _02796_);
  and (_19560_, _11633_, _05280_);
  or (_19561_, _19560_, _19549_);
  or (_19562_, _19561_, _02927_);
  and (_19563_, _19562_, _06189_);
  and (_19564_, _19563_, _19559_);
  and (_19565_, _11605_, _05280_);
  or (_19566_, _19565_, _19549_);
  and (_19567_, _19566_, _02790_);
  or (_19569_, _19567_, _19564_);
  and (_19570_, _19569_, _02966_);
  and (_19571_, _17300_, _05280_);
  or (_19572_, _19571_, _19549_);
  and (_19573_, _19572_, _02785_);
  or (_19574_, _19573_, _03861_);
  or (_19575_, _19574_, _19570_);
  and (_19576_, _19575_, _19534_);
  or (_19577_, _19576_, _03850_);
  and (_19578_, _05798_, _04681_);
  or (_19580_, _19528_, _06726_);
  or (_19581_, _19580_, _19578_);
  and (_19582_, _19581_, _02970_);
  and (_19583_, _19582_, _19577_);
  nor (_19584_, _11711_, _08690_);
  or (_19585_, _19584_, _19528_);
  and (_19586_, _19585_, _02524_);
  or (_19587_, _19586_, _02974_);
  or (_19588_, _19587_, _19583_);
  and (_19589_, _11718_, _04681_);
  or (_19591_, _19589_, _19528_);
  or (_19592_, _19591_, _05261_);
  and (_19593_, _19592_, _19588_);
  or (_19594_, _19593_, _02977_);
  and (_19595_, _11728_, _04681_);
  or (_19596_, _19528_, _07092_);
  or (_19597_, _19596_, _19595_);
  and (_19598_, _19597_, _07104_);
  and (_19599_, _19598_, _19594_);
  or (_19600_, _19599_, _19531_);
  and (_19602_, _19600_, _03095_);
  or (_19603_, _19528_, _04784_);
  and (_19604_, _19540_, _03094_);
  and (_19605_, _19591_, _02991_);
  or (_19606_, _19605_, _19604_);
  and (_19607_, _19606_, _19603_);
  or (_19608_, _19607_, _02994_);
  or (_19609_, _19608_, _19602_);
  nor (_19610_, _11726_, _08690_);
  or (_19611_, _19528_, _07120_);
  or (_19613_, _19611_, _19610_);
  and (_19614_, _19613_, _07118_);
  and (_19615_, _19614_, _19609_);
  nor (_19616_, _11600_, _08690_);
  or (_19617_, _19616_, _19528_);
  and (_19618_, _19617_, _03099_);
  or (_19619_, _19618_, _03133_);
  or (_19620_, _19619_, _19615_);
  or (_19621_, _19537_, _03138_);
  and (_19622_, _19621_, _03142_);
  and (_19624_, _19622_, _19620_);
  and (_19625_, _19561_, _02778_);
  or (_19626_, _19625_, _02852_);
  or (_19627_, _19626_, _19624_);
  and (_19628_, _11778_, _04681_);
  or (_19629_, _19528_, _02853_);
  or (_19630_, _19629_, _19628_);
  and (_19631_, _19630_, _34446_);
  and (_19632_, _19631_, _19627_);
  or (_35627_[6], _19632_, _19527_);
  not (_19634_, _10310_);
  and (_19635_, _19634_, _03471_);
  and (_19636_, _09696_, _09688_);
  nor (_19637_, _19636_, _02225_);
  and (_19638_, _09675_, _09667_);
  nor (_19639_, _19638_, _02225_);
  not (_19640_, _02575_);
  and (_19641_, _08795_, _09650_);
  nor (_19642_, _19641_, _02225_);
  nor (_19643_, _07743_, _02225_);
  and (_19645_, _07743_, _02225_);
  nor (_19646_, _19645_, _19643_);
  nor (_19647_, _19646_, _08800_);
  and (_19648_, _08805_, _07120_);
  nor (_19649_, _19648_, _02225_);
  and (_19650_, _08812_, _03881_);
  nor (_19651_, _19650_, _02225_);
  not (_19652_, _02582_);
  and (_19653_, _08822_, _07092_);
  nor (_19654_, _19653_, _02225_);
  and (_19656_, _02974_, _02225_);
  and (_19657_, _10325_, _08194_);
  nor (_19658_, _19657_, _02225_);
  nor (_19659_, _03471_, _02530_);
  nor (_19660_, _09273_, _02225_);
  nor (_19661_, _03471_, _02533_);
  nor (_19662_, _03471_, _02538_);
  nor (_19663_, _03471_, _02547_);
  not (_19664_, _07428_);
  and (_19665_, _09159_, _19664_);
  nor (_19667_, _19665_, _02225_);
  nor (_19668_, _19667_, _09178_);
  and (_19669_, _09164_, _02225_);
  nor (_19670_, _09164_, _02225_);
  nor (_19671_, _19670_, _19669_);
  and (_19672_, _19671_, _02546_);
  not (_19673_, _19672_);
  and (_19674_, _19673_, _19665_);
  not (_19675_, _19674_);
  and (_19676_, _19675_, _19668_);
  nor (_19678_, _19676_, _19663_);
  nor (_19679_, _19678_, _07425_);
  and (_19680_, _07425_, _02225_);
  nor (_19681_, _19680_, _05327_);
  not (_19682_, _19681_);
  nor (_19683_, _19682_, _19679_);
  and (_19684_, _02835_, _02225_);
  nor (_19685_, _19684_, _09095_);
  and (_19686_, _19685_, _09148_);
  and (_19687_, _05330_, _09146_);
  and (_19689_, _05328_, _05207_);
  and (_19690_, _19689_, _19687_);
  and (_19691_, _19690_, \oc8051_golden_model_1.PC [0]);
  or (_19692_, _19691_, _19686_);
  nor (_19693_, _19692_, _05325_);
  nor (_19694_, _19693_, _19683_);
  nor (_19695_, _19694_, _03806_);
  and (_19696_, _03806_, \oc8051_golden_model_1.PC [0]);
  nor (_19697_, _19696_, _02932_);
  not (_19698_, _19697_);
  nor (_19700_, _19698_, _19695_);
  not (_19701_, _19700_);
  and (_19702_, _03471_, \oc8051_golden_model_1.PC [0]);
  nor (_19703_, _19702_, _08911_);
  not (_19704_, _19703_);
  and (_19705_, _19704_, _09023_);
  and (_19706_, _09022_, _05036_);
  and (_19707_, _10821_, _04938_);
  and (_19708_, _19707_, _19706_);
  and (_19709_, _19708_, \oc8051_golden_model_1.PC [0]);
  or (_19711_, _19709_, _06162_);
  or (_19712_, _19711_, _19705_);
  and (_19713_, _19712_, _09018_);
  and (_19714_, _19713_, _19701_);
  nor (_19715_, _09018_, _02225_);
  nor (_19716_, _19715_, _04239_);
  not (_19717_, _19716_);
  nor (_19718_, _19717_, _19714_);
  nor (_19719_, _03471_, _02540_);
  and (_19720_, _09212_, _09199_);
  not (_19722_, _19720_);
  nor (_19723_, _19722_, _19719_);
  not (_19724_, _19723_);
  nor (_19725_, _19724_, _19718_);
  nor (_19726_, _19720_, _02225_);
  nor (_19727_, _19726_, _09209_);
  not (_19728_, _19727_);
  nor (_19729_, _19728_, _19725_);
  or (_19730_, _19729_, _09906_);
  nor (_19731_, _19730_, _19662_);
  and (_19733_, _09252_, _02225_);
  nor (_19734_, _19704_, _09252_);
  or (_19735_, _19734_, _09217_);
  nor (_19736_, _19735_, _19733_);
  nor (_19737_, _19736_, _02944_);
  not (_19738_, _19737_);
  nor (_19739_, _19738_, _19731_);
  nor (_19740_, _19739_, _02972_);
  and (_19741_, _09000_, _02225_);
  nor (_19742_, _19704_, _09000_);
  or (_19744_, _19742_, _09858_);
  nor (_19745_, _19744_, _19741_);
  nor (_19746_, _19745_, _19740_);
  and (_19747_, _09008_, _02225_);
  nor (_19748_, _19704_, _09008_);
  nor (_19749_, _19748_, _19747_);
  nor (_19750_, _19749_, _03397_);
  nor (_19751_, _19750_, _19746_);
  nor (_19752_, _19751_, _02979_);
  nor (_19753_, _19703_, _08839_);
  and (_19755_, _08839_, \oc8051_golden_model_1.PC [0]);
  or (_19756_, _19755_, _08969_);
  nor (_19757_, _19756_, _19753_);
  or (_19758_, _19757_, _19752_);
  and (_19759_, _19758_, _08828_);
  and (_19760_, _08827_, _02225_);
  or (_19761_, _19760_, _19759_);
  and (_19762_, _19761_, _02533_);
  or (_19763_, _19762_, _09281_);
  nor (_19764_, _19763_, _19661_);
  or (_19766_, _19764_, _09277_);
  nor (_19767_, _19766_, _19660_);
  and (_19768_, _09285_, _02499_);
  not (_19769_, _19768_);
  or (_19770_, _19769_, _19767_);
  nor (_19771_, _19770_, _19659_);
  nor (_19772_, _19768_, _02225_);
  nor (_19773_, _19772_, _02518_);
  not (_19774_, _19773_);
  nor (_19775_, _19774_, _19771_);
  nor (_19777_, _03471_, _04132_);
  not (_19778_, _19657_);
  nor (_19779_, _19778_, _19777_);
  not (_19780_, _19779_);
  nor (_19781_, _19780_, _19775_);
  or (_19782_, _19781_, _02578_);
  nor (_19783_, _19782_, _19658_);
  nor (_19784_, _03471_, _02579_);
  or (_19785_, _19784_, _09318_);
  nor (_19786_, _19785_, _19783_);
  nor (_19788_, _19685_, _09319_);
  nor (_19789_, _19788_, _19786_);
  and (_19790_, _19789_, _05261_);
  or (_19791_, _19790_, _19656_);
  and (_19792_, _19791_, _09335_);
  and (_19793_, _09334_, _02650_);
  or (_19794_, _19793_, _19792_);
  and (_19795_, _19794_, _04131_);
  nor (_19796_, _03471_, _04131_);
  or (_19797_, _19796_, _19795_);
  and (_19799_, _19797_, _09376_);
  not (_19800_, _19653_);
  and (_19801_, _08149_, \oc8051_golden_model_1.PC [0]);
  and (_19802_, _19685_, _09381_);
  or (_19803_, _19802_, _19801_);
  and (_19804_, _19803_, _09375_);
  nor (_19805_, _19804_, _19800_);
  not (_19806_, _19805_);
  nor (_19807_, _19806_, _19799_);
  nor (_19808_, _19807_, _19654_);
  and (_19810_, _19808_, _19652_);
  nor (_19811_, _03471_, _19652_);
  or (_19812_, _19811_, _19810_);
  and (_19813_, _19812_, _09398_);
  not (_19814_, _19650_);
  nor (_19815_, _19685_, _09381_);
  nor (_19816_, _08149_, \oc8051_golden_model_1.PC [0]);
  nor (_19817_, _19816_, _09398_);
  not (_19818_, _19817_);
  nor (_19819_, _19818_, _19815_);
  nor (_19821_, _19819_, _19814_);
  not (_19822_, _19821_);
  nor (_19823_, _19822_, _19813_);
  nor (_19824_, _19823_, _19651_);
  and (_19825_, _19824_, _10353_);
  nor (_19826_, _03471_, _10353_);
  or (_19827_, _19826_, _19825_);
  and (_19828_, _19827_, _08808_);
  not (_19829_, _19648_);
  and (_19830_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [0]);
  and (_19832_, _19685_, _07294_);
  or (_19833_, _19832_, _19830_);
  and (_19834_, _19833_, _08807_);
  nor (_19835_, _19834_, _19829_);
  not (_19836_, _19835_);
  nor (_19837_, _19836_, _19828_);
  nor (_19838_, _19837_, _19649_);
  and (_19839_, _19838_, _02590_);
  nor (_19840_, _03471_, _02590_);
  or (_19841_, _19840_, _19839_);
  and (_19843_, _19841_, _08800_);
  and (_19844_, _08797_, _08028_);
  not (_19845_, _19844_);
  or (_19846_, _19845_, _19843_);
  nor (_19847_, _19846_, _19647_);
  nor (_19848_, _19844_, _02225_);
  nor (_19849_, _19848_, _03113_);
  not (_19850_, _19849_);
  nor (_19851_, _19850_, _19847_);
  and (_19852_, _06114_, _03113_);
  or (_19854_, _19852_, _19851_);
  and (_19855_, _19854_, _05741_);
  nor (_19856_, _03471_, _05741_);
  or (_19857_, _19856_, _19855_);
  and (_19858_, _19857_, _03549_);
  and (_19859_, _19704_, _09640_);
  nor (_19860_, _09640_, _02225_);
  or (_19861_, _19860_, _03549_);
  or (_19862_, _19861_, _19859_);
  and (_19863_, _19862_, _19641_);
  not (_19865_, _19863_);
  nor (_19866_, _19865_, _19858_);
  nor (_19867_, _19866_, _19642_);
  and (_19868_, _19867_, _02855_);
  and (_19869_, _06114_, _02854_);
  or (_19870_, _19869_, _19868_);
  and (_19871_, _19870_, _19640_);
  nor (_19872_, _03471_, _19640_);
  nor (_19873_, _19872_, _19871_);
  nor (_19874_, _19873_, _02990_);
  not (_19876_, _19638_);
  and (_19877_, _09640_, \oc8051_golden_model_1.PC [0]);
  nor (_19878_, _19703_, _09640_);
  nor (_19879_, _19878_, _19877_);
  and (_19880_, _19879_, _02990_);
  nor (_19881_, _19880_, _19876_);
  not (_19882_, _19881_);
  nor (_19883_, _19882_, _19874_);
  nor (_19884_, _19883_, _19639_);
  nor (_19885_, _19884_, _04331_);
  and (_19887_, _04331_, _03471_);
  nor (_19888_, _19887_, _02778_);
  not (_19889_, _19888_);
  nor (_19890_, _19889_, _19885_);
  not (_19891_, _19636_);
  and (_19892_, _19879_, _02778_);
  nor (_19893_, _19892_, _19891_);
  not (_19894_, _19893_);
  nor (_19895_, _19894_, _19890_);
  nor (_19896_, _19895_, _19637_);
  nor (_19898_, _19896_, _19634_);
  or (_19899_, _19898_, _09706_);
  nor (_19900_, _19899_, _19635_);
  and (_19901_, _09706_, _02225_);
  nor (_19902_, _19901_, _19900_);
  nand (_19903_, _19902_, _34446_);
  or (_19904_, _34446_, \oc8051_golden_model_1.PC [0]);
  and (_19905_, _19904_, _35583_);
  and (_35629_[0], _19905_, _19903_);
  or (_19906_, _09675_, _08909_);
  or (_19907_, _08795_, _08909_);
  nor (_19908_, _07239_, _03518_);
  or (_19909_, _19908_, _08909_);
  or (_19910_, _08805_, _08909_);
  or (_19911_, _08812_, _08909_);
  and (_19912_, _14577_, _07828_);
  or (_19913_, _13411_, _08909_);
  or (_19914_, _05267_, _02198_);
  nand (_19915_, _02785_, \oc8051_golden_model_1.PC [1]);
  or (_19916_, _09285_, _08909_);
  or (_19918_, _03660_, _02533_);
  and (_19919_, _08827_, _02478_);
  nand (_19920_, _09252_, _02478_);
  nor (_19921_, _08913_, _08911_);
  nor (_19922_, _19921_, _08914_);
  not (_19923_, _19922_);
  or (_19924_, _19923_, _09252_);
  and (_19925_, _19924_, _19920_);
  and (_19926_, _19925_, _09906_);
  or (_19927_, _03660_, _02544_);
  and (_19929_, _09157_, _07413_);
  nor (_19930_, _19929_, _08909_);
  or (_19931_, _03660_, _02546_);
  nor (_19932_, _02837_, \oc8051_golden_model_1.PC [0]);
  or (_19933_, _19932_, _09168_);
  and (_19934_, _19933_, _02198_);
  nor (_19935_, _19933_, _02198_);
  or (_19936_, _19935_, _07415_);
  or (_19937_, _19936_, _19934_);
  nor (_19938_, _09162_, _08909_);
  or (_19940_, _19938_, _09163_);
  and (_19941_, _19940_, _19937_);
  and (_19942_, _09162_, _02478_);
  or (_19943_, _19942_, _02804_);
  or (_19944_, _19943_, _19941_);
  and (_19945_, _19944_, _19929_);
  and (_19946_, _19945_, _19931_);
  or (_19947_, _19946_, _19930_);
  and (_19948_, _19947_, _07408_);
  and (_19949_, _03343_, _02478_);
  or (_19950_, _19949_, _02934_);
  or (_19951_, _19950_, _19948_);
  and (_19952_, _02934_, _02198_);
  nor (_19953_, _19952_, _07428_);
  and (_19954_, _19953_, _19951_);
  and (_19955_, _07428_, _02478_);
  or (_19956_, _19955_, _09178_);
  or (_19957_, _19956_, _19954_);
  and (_19958_, _19957_, _19927_);
  or (_19959_, _19958_, _07425_);
  nand (_19961_, _07425_, _08909_);
  and (_19962_, _19961_, _05325_);
  and (_19963_, _19962_, _19959_);
  nor (_19964_, _09097_, _09095_);
  nor (_19965_, _19964_, _09098_);
  nand (_19966_, _19965_, _09148_);
  or (_19967_, _09148_, \oc8051_golden_model_1.PC [1]);
  and (_19968_, _19967_, _05327_);
  and (_19969_, _19968_, _19966_);
  or (_19970_, _19969_, _19963_);
  and (_19971_, _19970_, _05311_);
  and (_19972_, _03806_, _02478_);
  or (_19973_, _19972_, _02932_);
  or (_19974_, _19973_, _19971_);
  and (_19975_, _19923_, _09023_);
  and (_19976_, _09025_, _08909_);
  or (_19977_, _19976_, _06162_);
  or (_19978_, _19977_, _19975_);
  and (_19979_, _19978_, _09018_);
  and (_19980_, _19979_, _19974_);
  nor (_19982_, _09018_, _08909_);
  or (_19983_, _19982_, _02799_);
  or (_19984_, _19983_, _19980_);
  nand (_19985_, _02799_, _02198_);
  and (_19986_, _19985_, _02540_);
  and (_19987_, _19986_, _19984_);
  and (_19988_, _03660_, _04239_);
  or (_19989_, _19988_, _02930_);
  or (_19990_, _19989_, _19987_);
  nand (_19991_, _02930_, _02198_);
  and (_19993_, _19991_, _09199_);
  and (_19994_, _19993_, _19990_);
  nor (_19995_, _09199_, _08909_);
  or (_19996_, _19995_, _02928_);
  or (_19997_, _19996_, _19994_);
  and (_19998_, _02928_, _02198_);
  nor (_19999_, _19998_, _09206_);
  and (_20000_, _19999_, _19997_);
  and (_20001_, _09206_, _02478_);
  or (_20002_, _20001_, _02796_);
  or (_20003_, _20002_, _20000_);
  and (_20004_, _02538_, \oc8051_golden_model_1.PC [1]);
  or (_20005_, _20004_, _09210_);
  and (_20006_, _20005_, _20003_);
  and (_20007_, _03660_, _09209_);
  or (_20008_, _20007_, _02795_);
  or (_20009_, _20008_, _20006_);
  nand (_20010_, _02795_, _02198_);
  and (_20011_, _20010_, _09217_);
  and (_20012_, _20011_, _20009_);
  or (_20014_, _20012_, _19926_);
  and (_20015_, _20014_, _09858_);
  nand (_20016_, _09000_, _02478_);
  or (_20017_, _19923_, _09000_);
  and (_20018_, _20017_, _02972_);
  and (_20019_, _20018_, _20016_);
  or (_20020_, _20019_, _02944_);
  or (_20021_, _20020_, _20015_);
  or (_20022_, _19923_, _09008_);
  nand (_20023_, _09008_, _02478_);
  and (_20025_, _20023_, _20022_);
  or (_20026_, _20025_, _03397_);
  and (_20027_, _20026_, _20021_);
  or (_20028_, _20027_, _02979_);
  and (_20029_, _08839_, _08909_);
  nor (_20030_, _19922_, _08839_);
  or (_20031_, _20030_, _08969_);
  or (_20032_, _20031_, _20029_);
  and (_20033_, _20032_, _08828_);
  and (_20034_, _20033_, _20028_);
  or (_20035_, _20034_, _19919_);
  and (_20036_, _20035_, _06189_);
  and (_20037_, _02790_, \oc8051_golden_model_1.PC [1]);
  or (_20038_, _20037_, _04230_);
  or (_20039_, _20038_, _20036_);
  nand (_20040_, _20039_, _19918_);
  and (_20041_, _03231_, _02900_);
  nor (_20042_, _20041_, _02925_);
  and (_20043_, _03244_, _02900_);
  and (_20044_, _03680_, _02900_);
  nor (_20046_, _20044_, _20043_);
  and (_20047_, _20046_, _20042_);
  and (_20048_, _20047_, _04115_);
  and (_20049_, _20048_, _20040_);
  nor (_20050_, _20048_, \oc8051_golden_model_1.PC [1]);
  or (_20051_, _20050_, _09281_);
  or (_20052_, _20051_, _20049_);
  or (_20053_, _09273_, _08909_);
  and (_20054_, _20053_, _09276_);
  and (_20055_, _20054_, _20052_);
  and (_20057_, _02902_, _02198_);
  or (_20058_, _20057_, _09277_);
  or (_20059_, _20058_, _20055_);
  nand (_20060_, _03660_, _09277_);
  and (_20061_, _20060_, _09759_);
  and (_20062_, _20061_, _20059_);
  nand (_20063_, _02901_, _02198_);
  nand (_20064_, _20063_, _09285_);
  or (_20065_, _20064_, _20062_);
  and (_20066_, _20065_, _19916_);
  or (_20067_, _20066_, _09290_);
  or (_20068_, _09289_, _02198_);
  and (_20069_, _20068_, _02499_);
  and (_20070_, _20069_, _20067_);
  nor (_20071_, _02499_, _02478_);
  or (_20072_, _20071_, _02785_);
  or (_20073_, _20072_, _20070_);
  and (_20074_, _20073_, _19915_);
  or (_20075_, _20074_, _02518_);
  nand (_20076_, _03660_, _02518_);
  and (_20078_, _20076_, _08194_);
  and (_20079_, _20078_, _20075_);
  nand (_20080_, _02975_, _02478_);
  nand (_20081_, _20080_, _09305_);
  or (_20082_, _20081_, _20079_);
  or (_20083_, _09305_, _02198_);
  and (_20084_, _20083_, _02970_);
  and (_20085_, _20084_, _20082_);
  nor (_20086_, _08824_, _02478_);
  nor (_20087_, _20086_, _10325_);
  or (_20089_, _20087_, _20085_);
  nand (_20090_, _08824_, _02478_);
  and (_20091_, _20090_, _03474_);
  and (_20092_, _20091_, _20089_);
  and (_20093_, _02894_, _02198_);
  or (_20094_, _20093_, _02578_);
  or (_20095_, _20094_, _20092_);
  nand (_20096_, _03660_, _02578_);
  and (_20097_, _20096_, _09319_);
  and (_20098_, _20097_, _20095_);
  and (_20099_, _19965_, _09318_);
  or (_20100_, _20099_, _05516_);
  or (_20101_, _20100_, _20098_);
  and (_20102_, _20101_, _19914_);
  or (_20103_, _20102_, _02974_);
  nand (_20104_, _02974_, _08909_);
  and (_20105_, _20104_, _07808_);
  and (_20106_, _20105_, _20103_);
  and (_20107_, _07807_, _02198_);
  or (_20108_, _20107_, _09334_);
  or (_20110_, _20108_, _20106_);
  or (_20111_, _09335_, _02671_);
  and (_20112_, _20111_, _10067_);
  and (_20113_, _20112_, _20110_);
  and (_20114_, _02893_, _02198_);
  or (_20115_, _20114_, _02585_);
  or (_20116_, _20115_, _20113_);
  nand (_20117_, _03660_, _02585_);
  and (_20118_, _20117_, _09376_);
  and (_20119_, _20118_, _20116_);
  or (_20121_, _19965_, _08149_);
  nand (_20122_, _08149_, \oc8051_golden_model_1.PC [1]);
  and (_20123_, _20122_, _09375_);
  and (_20124_, _20123_, _20121_);
  or (_20125_, _20124_, _13413_);
  or (_20126_, _20125_, _20119_);
  nand (_20127_, _20126_, _19913_);
  nand (_20128_, _20127_, _19912_);
  or (_20129_, _19912_, _08909_);
  and (_20130_, _20129_, _03487_);
  and (_20131_, _20130_, _20128_);
  nand (_20132_, _03486_, _08909_);
  nand (_20133_, _20132_, _08814_);
  or (_20134_, _20133_, _20131_);
  or (_20135_, _08814_, _02198_);
  and (_20136_, _20135_, _07092_);
  and (_20137_, _20136_, _20134_);
  and (_20138_, _02977_, _02478_);
  or (_20139_, _20138_, _03107_);
  or (_20140_, _20139_, _20137_);
  nand (_20142_, _03107_, \oc8051_golden_model_1.PC [1]);
  and (_20143_, _20142_, _20140_);
  or (_20144_, _20143_, _02582_);
  nand (_20145_, _03660_, _02582_);
  and (_20146_, _20145_, _09398_);
  and (_20147_, _20146_, _20144_);
  or (_20148_, _19965_, _09381_);
  or (_20149_, _08149_, _02198_);
  and (_20150_, _20149_, _09397_);
  and (_20151_, _20150_, _20148_);
  or (_20153_, _20151_, _09406_);
  or (_20154_, _20153_, _20147_);
  and (_20155_, _20154_, _19911_);
  or (_20156_, _20155_, _07882_);
  or (_20157_, _07881_, _02198_);
  and (_20158_, _20157_, _03881_);
  and (_20159_, _20158_, _20156_);
  and (_20160_, _02991_, _02478_);
  or (_20161_, _20160_, _03094_);
  or (_20162_, _20161_, _20159_);
  nand (_20163_, _03094_, \oc8051_golden_model_1.PC [1]);
  and (_20164_, _20163_, _20162_);
  or (_20165_, _20164_, _02594_);
  nand (_20166_, _03660_, _02594_);
  and (_20167_, _20166_, _08808_);
  and (_20168_, _20167_, _20165_);
  or (_20169_, _19965_, \oc8051_golden_model_1.PSW [7]);
  nand (_20170_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.PC [1]);
  and (_20171_, _20170_, _08807_);
  and (_20172_, _20171_, _20169_);
  or (_20174_, _20172_, _09418_);
  or (_20175_, _20174_, _20168_);
  and (_20176_, _20175_, _19910_);
  or (_20177_, _20176_, _07901_);
  or (_20178_, _07900_, _02198_);
  and (_20179_, _20178_, _07120_);
  and (_20180_, _20179_, _20177_);
  and (_20181_, _02994_, _02478_);
  or (_20182_, _20181_, _03099_);
  or (_20183_, _20182_, _20180_);
  nand (_20185_, _03099_, \oc8051_golden_model_1.PC [1]);
  and (_20186_, _20185_, _20183_);
  or (_20187_, _20186_, _02589_);
  nand (_20188_, _03660_, _02589_);
  and (_20189_, _20188_, _08800_);
  and (_20190_, _20189_, _20187_);
  or (_20191_, _19965_, _07294_);
  or (_20192_, \oc8051_golden_model_1.PSW [7], _02198_);
  and (_20193_, _20192_, _08799_);
  nand (_20194_, _20193_, _20191_);
  nand (_20195_, _20194_, _19908_);
  or (_20196_, _20195_, _20190_);
  nand (_20197_, _20196_, _19909_);
  and (_20198_, _03495_, _02591_);
  and (_20199_, _10346_, _02591_);
  nor (_20200_, _20199_, _20198_);
  nand (_20201_, _20200_, _20197_);
  not (_20202_, _03512_);
  or (_20203_, _20200_, _08909_);
  and (_20204_, _20203_, _20202_);
  and (_20206_, _20204_, _20201_);
  nand (_20207_, _03512_, _08909_);
  nand (_20208_, _20207_, _07947_);
  or (_20209_, _20208_, _20206_);
  or (_20210_, _07947_, _02198_);
  and (_20211_, _20210_, _08028_);
  and (_20212_, _20211_, _20209_);
  and (_20213_, _08027_, _08909_);
  or (_20214_, _20213_, _03113_);
  or (_20215_, _20214_, _20212_);
  or (_20217_, _06113_, _10159_);
  and (_20218_, _20217_, _20215_);
  or (_20219_, _20218_, _02592_);
  nand (_20220_, _03660_, _02592_);
  and (_20221_, _20220_, _03549_);
  and (_20222_, _20221_, _20219_);
  nand (_20223_, _19923_, _09640_);
  or (_20224_, _09640_, _02478_);
  and (_20225_, _20224_, _02993_);
  and (_20226_, _20225_, _20223_);
  or (_20227_, _20226_, _09455_);
  or (_20228_, _20227_, _20222_);
  and (_20229_, _20228_, _19907_);
  or (_20230_, _20229_, _08772_);
  nand (_20231_, _08772_, \oc8051_golden_model_1.PC [1]);
  and (_20232_, _20231_, _09650_);
  and (_20233_, _20232_, _20230_);
  and (_20234_, _07143_, _08909_);
  or (_20235_, _20234_, _02854_);
  or (_20236_, _20235_, _20233_);
  or (_20238_, _06113_, _02855_);
  and (_20239_, _20238_, _20236_);
  or (_20240_, _20239_, _02575_);
  nand (_20241_, _03660_, _02575_);
  and (_20242_, _20241_, _03134_);
  and (_20243_, _20242_, _20240_);
  nand (_20244_, _09640_, _08909_);
  or (_20245_, _19922_, _09640_);
  and (_20246_, _20245_, _20244_);
  nand (_20247_, _20246_, _02990_);
  nand (_20249_, _20247_, _04109_);
  or (_20250_, _20249_, _20243_);
  nor (_20251_, _04109_, _08909_);
  and (_20252_, _04120_, _02571_);
  nor (_20253_, _20252_, _20251_);
  and (_20254_, _20253_, _20250_);
  nor (_20255_, _03898_, _03557_);
  nand (_20256_, _20252_, _08909_);
  nand (_20257_, _20256_, _20255_);
  or (_20258_, _20257_, _20254_);
  or (_20259_, _20255_, _08909_);
  and (_20260_, _20259_, _03138_);
  and (_20261_, _20260_, _20258_);
  nand (_20262_, _03133_, _02198_);
  nand (_20263_, _20262_, _09675_);
  or (_20264_, _20263_, _20261_);
  and (_20265_, _20264_, _19906_);
  or (_20266_, _20265_, _04331_);
  nand (_20267_, _04331_, _03660_);
  and (_20268_, _20267_, _03142_);
  and (_20270_, _20268_, _20266_);
  and (_20271_, _20246_, _02778_);
  or (_20272_, _20271_, _10780_);
  or (_20273_, _20272_, _20270_);
  nand (_20274_, _10780_, _02478_);
  nand (_20275_, _20274_, _20273_);
  nor (_20276_, _03581_, _03912_);
  nand (_20277_, _20276_, _20275_);
  or (_20278_, _20276_, _08909_);
  and (_20279_, _20278_, _02853_);
  and (_20281_, _20279_, _20277_);
  and (_20282_, _02852_, _02198_);
  or (_20283_, _20282_, _20281_);
  and (_20284_, _20283_, _09696_);
  nor (_20285_, _09696_, _02478_);
  or (_20286_, _20285_, _19634_);
  or (_20287_, _20286_, _20284_);
  and (_20288_, _19634_, _03660_);
  nor (_20289_, _20288_, _09706_);
  and (_20290_, _20289_, _20287_);
  and (_20291_, _09706_, _08909_);
  or (_20292_, _20291_, _20290_);
  or (_20293_, _20292_, _34450_);
  or (_20294_, _34446_, \oc8051_golden_model_1.PC [1]);
  and (_20295_, _20294_, _35583_);
  and (_35629_[1], _20295_, _20293_);
  and (_20296_, _03133_, _02555_);
  not (_20297_, _08772_);
  nor (_20298_, _08795_, _02487_);
  nor (_20299_, _08797_, _02487_);
  nor (_20301_, _08805_, _02487_);
  nor (_20302_, _08812_, _02487_);
  nor (_20303_, _08822_, _02487_);
  nor (_20304_, _05266_, _02555_);
  not (_20305_, _02487_);
  and (_20306_, _08824_, _20305_);
  not (_20307_, _03856_);
  nor (_20308_, _20307_, _03435_);
  nor (_20309_, _20308_, _02555_);
  and (_20310_, _02600_, _02785_);
  nor (_20312_, _20048_, _02555_);
  and (_20313_, _08827_, _20305_);
  and (_20314_, _08918_, _08915_);
  nor (_20315_, _20314_, _08919_);
  not (_20316_, _20315_);
  nor (_20317_, _20316_, _09000_);
  and (_20318_, _09000_, _08906_);
  nor (_20319_, _20318_, _20317_);
  nor (_20320_, _20319_, _09858_);
  not (_20321_, _20320_);
  nor (_20323_, _20316_, _09008_);
  and (_20324_, _09008_, _08906_);
  nor (_20325_, _20324_, _20323_);
  nor (_20326_, _20325_, _03397_);
  or (_20327_, _20316_, _09025_);
  or (_20328_, _09023_, _08907_);
  and (_20329_, _20328_, _02932_);
  and (_20330_, _20329_, _20327_);
  and (_20331_, _09102_, _09099_);
  nor (_20332_, _20331_, _09103_);
  and (_20333_, _20332_, _09148_);
  and (_20334_, _19690_, _02555_);
  nor (_20335_, _20334_, _20333_);
  nand (_20336_, _20335_, _05327_);
  nor (_20337_, _03223_, _02544_);
  and (_20338_, _02934_, _02555_);
  nor (_20339_, _03223_, _02546_);
  not (_20340_, _09159_);
  not (_20341_, _09163_);
  and (_20342_, _09168_, \oc8051_golden_model_1.PC [2]);
  and (_20344_, _02837_, _02555_);
  nor (_20345_, _20344_, _20342_);
  nor (_20346_, _20345_, _20341_);
  nor (_20347_, _09164_, _20305_);
  nor (_20348_, _20347_, _20346_);
  nor (_20349_, _20348_, _02804_);
  nor (_20350_, _20349_, _20340_);
  not (_20351_, _20350_);
  nor (_20352_, _20351_, _20339_);
  nor (_20353_, _09159_, _02487_);
  nor (_20355_, _20353_, _02934_);
  not (_20356_, _20355_);
  nor (_20357_, _20356_, _20352_);
  or (_20358_, _20357_, _07428_);
  nor (_20359_, _20358_, _20338_);
  and (_20360_, _07428_, _20305_);
  nor (_20361_, _20360_, _09178_);
  not (_20362_, _20361_);
  nor (_20363_, _20362_, _20359_);
  nor (_20364_, _20363_, _20337_);
  nor (_20365_, _20364_, _07425_);
  and (_20366_, _07425_, _02487_);
  nor (_20367_, _20366_, _05327_);
  not (_20368_, _20367_);
  nor (_20369_, _20368_, _20365_);
  nor (_20370_, _20369_, _03806_);
  nand (_20371_, _20370_, _20336_);
  nand (_20372_, _03806_, _02487_);
  and (_20373_, _20372_, _06162_);
  and (_20374_, _20373_, _20371_);
  or (_20376_, _20374_, _20330_);
  nand (_20377_, _20376_, _09018_);
  nor (_20378_, _09018_, _02487_);
  nor (_20379_, _20378_, _02799_);
  and (_20380_, _20379_, _20377_);
  and (_20381_, _02799_, _02555_);
  or (_20382_, _20381_, _04239_);
  or (_20383_, _20382_, _20380_);
  and (_20384_, _03223_, _04239_);
  nor (_20385_, _20384_, _02930_);
  nand (_20387_, _20385_, _20383_);
  and (_20388_, _02930_, _02555_);
  nor (_20389_, _20388_, _09200_);
  nand (_20390_, _20389_, _20387_);
  nor (_20391_, _09199_, _02487_);
  nor (_20392_, _20391_, _02928_);
  nand (_20393_, _20392_, _20390_);
  and (_20394_, _02928_, _02555_);
  nor (_20395_, _20394_, _09206_);
  nand (_20396_, _20395_, _20393_);
  and (_20398_, _09206_, _20305_);
  nor (_20399_, _20398_, _02796_);
  and (_20400_, _20399_, _20396_);
  and (_20401_, _02796_, _02555_);
  or (_20402_, _20401_, _09209_);
  or (_20403_, _20402_, _20400_);
  and (_20404_, _03223_, _09209_);
  nor (_20405_, _20404_, _02795_);
  nand (_20406_, _20405_, _20403_);
  and (_20407_, _02795_, _02555_);
  nor (_20408_, _20407_, _09906_);
  and (_20409_, _20408_, _20406_);
  nor (_20410_, _20316_, _09252_);
  and (_20411_, _09252_, _08906_);
  nor (_20412_, _20411_, _20410_);
  and (_20413_, _20412_, _09906_);
  nor (_20414_, _20413_, _20409_);
  and (_20415_, _20414_, _02973_);
  nor (_20416_, _20415_, _20326_);
  nand (_20417_, _20416_, _20321_);
  nand (_20419_, _20417_, _08969_);
  nor (_20420_, _20315_, _08839_);
  and (_20421_, _08907_, _08839_);
  or (_20422_, _20421_, _08969_);
  or (_20423_, _20422_, _20420_);
  and (_20424_, _20423_, _08828_);
  and (_20425_, _20424_, _20419_);
  or (_20426_, _20425_, _20313_);
  nand (_20427_, _20426_, _06189_);
  and (_20428_, _02790_, _02600_);
  nor (_20430_, _20428_, _04230_);
  nand (_20431_, _20430_, _20427_);
  not (_20432_, _20048_);
  nor (_20433_, _03223_, _02533_);
  nor (_20434_, _20433_, _20432_);
  and (_20435_, _20434_, _20431_);
  or (_20436_, _20435_, _20312_);
  nand (_20437_, _20436_, _09273_);
  nor (_20438_, _09273_, _02487_);
  nor (_20439_, _20438_, _02902_);
  nand (_20440_, _20439_, _20437_);
  and (_20441_, _02902_, _02555_);
  nor (_20442_, _20441_, _09277_);
  nand (_20443_, _20442_, _20440_);
  and (_20444_, _03223_, _09277_);
  nor (_20445_, _20444_, _02901_);
  nand (_20446_, _20445_, _20443_);
  not (_20447_, _09285_);
  and (_20448_, _02901_, _02555_);
  nor (_20449_, _20448_, _20447_);
  and (_20451_, _20449_, _20446_);
  nor (_20452_, _09285_, _02487_);
  or (_20453_, _20452_, _20451_);
  nand (_20454_, _20453_, _09289_);
  nor (_20455_, _09289_, _02555_);
  nor (_20456_, _20455_, _07700_);
  nand (_20457_, _20456_, _20454_);
  nor (_20458_, _02499_, _20305_);
  nor (_20459_, _20458_, _02785_);
  and (_20460_, _20459_, _20457_);
  or (_20462_, _20460_, _20310_);
  nand (_20463_, _20462_, _04132_);
  and (_20464_, _03223_, _02518_);
  nor (_20465_, _20464_, _02975_);
  nand (_20466_, _20465_, _20463_);
  and (_20467_, _08906_, _02975_);
  not (_20468_, _20467_);
  and (_20469_, _20468_, _20308_);
  and (_20470_, _20469_, _20466_);
  or (_20471_, _20470_, _20309_);
  nor (_20473_, _04158_, _03850_);
  nand (_20474_, _20473_, _20471_);
  nor (_20475_, _20473_, _02555_);
  nor (_20476_, _20475_, _02524_);
  and (_20477_, _20476_, _20474_);
  and (_20478_, _08906_, _02524_);
  or (_20479_, _20478_, _08824_);
  nor (_20480_, _20479_, _20477_);
  or (_20481_, _20480_, _20306_);
  nand (_20482_, _20481_, _03474_);
  and (_20484_, _02894_, _02600_);
  nor (_20485_, _20484_, _02578_);
  and (_20486_, _20485_, _20482_);
  nor (_20487_, _03223_, _02579_);
  or (_20488_, _20487_, _20486_);
  nand (_20489_, _20488_, _09319_);
  not (_20490_, _05266_);
  and (_20491_, _20332_, _09318_);
  nor (_20492_, _20491_, _20490_);
  and (_20493_, _20492_, _20489_);
  or (_20495_, _20493_, _20304_);
  nand (_20496_, _20495_, _05262_);
  and (_20497_, _03870_, _02600_);
  nor (_20498_, _20497_, _02974_);
  and (_20499_, _20498_, _20496_);
  and (_20500_, _08906_, _02974_);
  or (_20501_, _20500_, _07807_);
  nor (_20502_, _20501_, _20499_);
  and (_20503_, _07807_, _02600_);
  or (_20504_, _20503_, _20502_);
  nand (_20506_, _20504_, _09335_);
  and (_20507_, _09334_, _02513_);
  nor (_20508_, _20507_, _02893_);
  nand (_20509_, _20508_, _20506_);
  and (_20510_, _02893_, _02555_);
  nor (_20511_, _20510_, _02585_);
  nand (_20512_, _20511_, _20509_);
  and (_20513_, _03223_, _02585_);
  nor (_20514_, _20513_, _09375_);
  nand (_20515_, _20514_, _20512_);
  and (_20517_, _08149_, _02555_);
  and (_20518_, _20332_, _09381_);
  or (_20519_, _20518_, _20517_);
  and (_20520_, _20519_, _09375_);
  nor (_20521_, _20520_, _09385_);
  and (_20522_, _20521_, _20515_);
  or (_20523_, _20522_, _20303_);
  nand (_20524_, _20523_, _08814_);
  nor (_20525_, _08814_, _02555_);
  nor (_20526_, _20525_, _02977_);
  and (_20528_, _20526_, _20524_);
  and (_20529_, _08906_, _02977_);
  or (_20530_, _20529_, _03107_);
  nor (_20531_, _20530_, _20528_);
  and (_20532_, _03107_, _02600_);
  or (_20533_, _20532_, _20531_);
  nand (_20534_, _20533_, _19652_);
  and (_20535_, _03223_, _02582_);
  nor (_20536_, _20535_, _09397_);
  nand (_20537_, _20536_, _20534_);
  or (_20539_, _20332_, _09381_);
  or (_20540_, _08149_, _02555_);
  and (_20541_, _20540_, _09397_);
  and (_20542_, _20541_, _20539_);
  nor (_20543_, _20542_, _09406_);
  and (_20544_, _20543_, _20537_);
  or (_20545_, _20544_, _20302_);
  nand (_20546_, _20545_, _07881_);
  nor (_20547_, _07881_, _02555_);
  nor (_20548_, _20547_, _02991_);
  and (_20549_, _20548_, _20546_);
  and (_20550_, _08906_, _02991_);
  or (_20551_, _20550_, _03094_);
  nor (_20552_, _20551_, _20549_);
  and (_20553_, _03094_, _02600_);
  or (_20554_, _20553_, _20552_);
  nand (_20555_, _20554_, _10353_);
  and (_20556_, _03223_, _02594_);
  nor (_20557_, _20556_, _08807_);
  nand (_20558_, _20557_, _20555_);
  nor (_20559_, _20332_, \oc8051_golden_model_1.PSW [7]);
  nor (_20560_, _02555_, _07294_);
  nor (_20561_, _20560_, _08808_);
  not (_20562_, _20561_);
  nor (_20563_, _20562_, _20559_);
  nor (_20564_, _20563_, _09418_);
  and (_20565_, _20564_, _20558_);
  or (_20566_, _20565_, _20301_);
  nand (_20567_, _20566_, _07900_);
  nor (_20568_, _07900_, _02555_);
  nor (_20570_, _20568_, _02994_);
  nand (_20571_, _20570_, _20567_);
  and (_20572_, _08906_, _02994_);
  nor (_20573_, _20572_, _03099_);
  and (_20574_, _20573_, _20571_);
  and (_20575_, _03099_, _02600_);
  or (_20576_, _20575_, _20574_);
  nand (_20577_, _20576_, _02590_);
  and (_20578_, _03223_, _02589_);
  nor (_20579_, _20578_, _08799_);
  nand (_20581_, _20579_, _20577_);
  and (_20582_, _02555_, _07294_);
  and (_20583_, _20332_, \oc8051_golden_model_1.PSW [7]);
  or (_20584_, _20583_, _20582_);
  and (_20585_, _20584_, _08799_);
  nor (_20586_, _20585_, _09434_);
  and (_20587_, _20586_, _20581_);
  or (_20588_, _20587_, _20299_);
  nand (_20589_, _20588_, _07947_);
  nor (_20590_, _07947_, _02555_);
  nor (_20592_, _20590_, _08027_);
  nand (_20593_, _20592_, _20589_);
  and (_20594_, _08027_, _02487_);
  nor (_20595_, _20594_, _03113_);
  and (_20596_, _20595_, _20593_);
  and (_20597_, _05980_, _03113_);
  or (_20598_, _20597_, _20596_);
  nand (_20599_, _20598_, _05741_);
  and (_20600_, _03223_, _02592_);
  nor (_20601_, _20600_, _02993_);
  nand (_20603_, _20601_, _20599_);
  nor (_20604_, _09640_, _08906_);
  and (_20605_, _20316_, _09640_);
  or (_20606_, _20605_, _03549_);
  or (_20607_, _20606_, _20604_);
  and (_20608_, _20607_, _08795_);
  and (_20609_, _20608_, _20603_);
  or (_20610_, _20609_, _20298_);
  nand (_20611_, _20610_, _20297_);
  and (_20612_, _08772_, _02600_);
  nor (_20614_, _20612_, _07143_);
  nand (_20615_, _20614_, _20611_);
  and (_20616_, _07143_, _02487_);
  nor (_20617_, _20616_, _02854_);
  and (_20618_, _20617_, _20615_);
  and (_20619_, _05980_, _02854_);
  or (_20620_, _20619_, _20618_);
  nand (_20621_, _20620_, _19640_);
  and (_20622_, _03223_, _02575_);
  nor (_20623_, _20622_, _02990_);
  nand (_20625_, _20623_, _20621_);
  nor (_20626_, _20315_, _09640_);
  and (_20627_, _09640_, _08907_);
  nor (_20628_, _20627_, _20626_);
  and (_20629_, _20628_, _02990_);
  nor (_20630_, _20629_, _09668_);
  nand (_20631_, _20630_, _20625_);
  nor (_20632_, _09667_, _02487_);
  nor (_20633_, _20632_, _03133_);
  and (_20634_, _20633_, _20631_);
  or (_20636_, _20634_, _20296_);
  nand (_20637_, _20636_, _09675_);
  nor (_20638_, _09675_, _20305_);
  nor (_20639_, _20638_, _04331_);
  nand (_20640_, _20639_, _20637_);
  and (_20641_, _04331_, _03223_);
  nor (_20642_, _20641_, _02778_);
  and (_20643_, _20642_, _20640_);
  nor (_20644_, _20628_, _09689_);
  nor (_20645_, _20644_, _10370_);
  or (_20647_, _20645_, _20643_);
  nor (_20648_, _09688_, _02487_);
  nor (_20649_, _20648_, _02852_);
  and (_20650_, _20649_, _20647_);
  and (_20651_, _09696_, _02600_);
  nor (_20652_, _20651_, _10371_);
  nor (_20653_, _20652_, _20650_);
  nor (_20654_, _09696_, _02487_);
  or (_20655_, _20654_, _20653_);
  nand (_20656_, _20655_, _10310_);
  and (_20658_, _19634_, _03223_);
  nor (_20659_, _20658_, _09706_);
  and (_20660_, _20659_, _20656_);
  and (_20661_, _09706_, _02487_);
  or (_20662_, _20661_, _20660_);
  or (_20663_, _20662_, _34450_);
  or (_20664_, _34446_, \oc8051_golden_model_1.PC [2]);
  and (_20665_, _20664_, _35583_);
  and (_35629_[2], _20665_, _20663_);
  and (_20666_, _03133_, _02620_);
  and (_20668_, _05935_, _02854_);
  nor (_20669_, _08795_, _02616_);
  nor (_20670_, _08797_, _02616_);
  nor (_20671_, _08805_, _02616_);
  nor (_20672_, _08812_, _02616_);
  nor (_20673_, _08822_, _02616_);
  nor (_20674_, _05267_, _02620_);
  nor (_20675_, _20048_, _02620_);
  and (_20676_, _08827_, _02608_);
  and (_20677_, _09252_, _08901_);
  or (_20679_, _08904_, _08903_);
  and (_20680_, _20679_, _08920_);
  nor (_20681_, _20679_, _08920_);
  nor (_20682_, _20681_, _20680_);
  not (_20683_, _20682_);
  nor (_20684_, _20683_, _09252_);
  or (_20685_, _20684_, _20677_);
  nor (_20686_, _20685_, _09217_);
  or (_20687_, _09023_, _08901_);
  or (_20688_, _20682_, _09025_);
  and (_20690_, _20688_, _20687_);
  or (_20691_, _20690_, _06162_);
  or (_20692_, _09092_, _09091_);
  and (_20693_, _20692_, _09104_);
  nor (_20694_, _20692_, _09104_);
  nor (_20695_, _20694_, _20693_);
  and (_20696_, _20695_, _09148_);
  and (_20697_, _09150_, _02620_);
  nor (_20698_, _20697_, _20696_);
  nand (_20699_, _20698_, _05327_);
  nor (_20701_, _03087_, _02544_);
  nor (_20702_, _03087_, _02546_);
  and (_20703_, _09168_, \oc8051_golden_model_1.PC [3]);
  and (_20704_, _02837_, _02620_);
  nor (_20705_, _20704_, _20703_);
  nor (_20706_, _20705_, _20341_);
  nor (_20707_, _09164_, _02608_);
  nor (_20708_, _20707_, _20706_);
  nor (_20709_, _20708_, _02804_);
  nor (_20710_, _20709_, _20340_);
  not (_20712_, _20710_);
  nor (_20713_, _20712_, _20702_);
  nor (_20714_, _09159_, _02616_);
  nor (_20715_, _20714_, _02934_);
  not (_20716_, _20715_);
  nor (_20717_, _20716_, _20713_);
  nor (_20718_, _07428_, _02934_);
  nor (_20719_, _07428_, _02620_);
  nor (_20720_, _20719_, _20718_);
  nor (_20721_, _20720_, _20717_);
  and (_20723_, _07428_, _02608_);
  nor (_20724_, _20723_, _09178_);
  not (_20725_, _20724_);
  nor (_20726_, _20725_, _20721_);
  nor (_20727_, _20726_, _20701_);
  nor (_20728_, _20727_, _07425_);
  and (_20729_, _07425_, _02616_);
  nor (_20730_, _20729_, _05327_);
  not (_20731_, _20730_);
  nor (_20732_, _20731_, _20728_);
  nor (_20734_, _20732_, _03806_);
  and (_20735_, _20734_, _20699_);
  and (_20736_, _03806_, _02616_);
  or (_20737_, _20736_, _02932_);
  or (_20738_, _20737_, _20735_);
  nand (_20739_, _20738_, _20691_);
  nand (_20740_, _20739_, _09018_);
  nor (_20741_, _09018_, _02616_);
  nor (_20742_, _20741_, _02799_);
  and (_20743_, _20742_, _20740_);
  and (_20745_, _02799_, _02620_);
  or (_20746_, _20745_, _04239_);
  or (_20747_, _20746_, _20743_);
  and (_20748_, _03087_, _04239_);
  nor (_20749_, _20748_, _02930_);
  nand (_20750_, _20749_, _20747_);
  and (_20751_, _02930_, _02620_);
  nor (_20752_, _20751_, _09200_);
  nand (_20753_, _20752_, _20750_);
  nor (_20754_, _09199_, _02616_);
  nor (_20756_, _20754_, _02928_);
  nand (_20757_, _20756_, _20753_);
  and (_20758_, _02928_, _02620_);
  nor (_20759_, _20758_, _09206_);
  nand (_20760_, _20759_, _20757_);
  and (_20761_, _09206_, _02608_);
  nor (_20762_, _20761_, _02796_);
  nand (_20763_, _20762_, _20760_);
  and (_20764_, _02796_, _02620_);
  nor (_20765_, _20764_, _09209_);
  nand (_20767_, _20765_, _20763_);
  and (_20768_, _03087_, _09209_);
  nor (_20769_, _20768_, _02795_);
  nand (_20770_, _20769_, _20767_);
  and (_20771_, _02795_, _02620_);
  nor (_20772_, _20771_, _09906_);
  and (_20773_, _20772_, _20770_);
  or (_20774_, _20773_, _20686_);
  nand (_20775_, _20774_, _09858_);
  and (_20776_, _09000_, _08901_);
  nor (_20778_, _20683_, _09000_);
  nor (_20779_, _20778_, _20776_);
  nand (_20780_, _20779_, _02972_);
  and (_20781_, _20780_, _09927_);
  and (_20782_, _20781_, _20775_);
  and (_20783_, _09008_, _08901_);
  nor (_20784_, _20683_, _09008_);
  nor (_20785_, _20784_, _20783_);
  nor (_20786_, _20785_, _03397_);
  not (_20787_, _20786_);
  and (_20789_, _08902_, _08839_);
  nor (_20790_, _20682_, _08839_);
  or (_20791_, _20790_, _08969_);
  nor (_20792_, _20791_, _20789_);
  nor (_20793_, _20792_, _08827_);
  nand (_20794_, _20793_, _20787_);
  nor (_20795_, _20794_, _20782_);
  or (_20796_, _20795_, _20676_);
  nand (_20797_, _20796_, _06189_);
  and (_20798_, _02790_, _02641_);
  nor (_20800_, _20798_, _04230_);
  nand (_20801_, _20800_, _20797_);
  nor (_20802_, _03087_, _02533_);
  nor (_20803_, _20802_, _20432_);
  and (_20804_, _20803_, _20801_);
  or (_20805_, _20804_, _20675_);
  nand (_20806_, _20805_, _09273_);
  nor (_20807_, _09273_, _02616_);
  nor (_20808_, _20807_, _02902_);
  nand (_20809_, _20808_, _20806_);
  and (_20811_, _02902_, _02620_);
  nor (_20812_, _20811_, _09277_);
  nand (_20813_, _20812_, _20809_);
  and (_20814_, _03087_, _09277_);
  nor (_20815_, _20814_, _02901_);
  nand (_20816_, _20815_, _20813_);
  and (_20817_, _02901_, _02620_);
  nor (_20818_, _20817_, _20447_);
  and (_20819_, _20818_, _20816_);
  nor (_20820_, _09285_, _02616_);
  or (_20822_, _20820_, _20819_);
  nand (_20823_, _20822_, _09289_);
  nor (_20824_, _09289_, _02620_);
  nor (_20825_, _20824_, _07700_);
  and (_20826_, _20825_, _20823_);
  nor (_20827_, _02499_, _02608_);
  or (_20828_, _20827_, _02785_);
  nor (_20829_, _20828_, _20826_);
  and (_20830_, _02641_, _02785_);
  or (_20831_, _20830_, _20829_);
  nand (_20833_, _20831_, _04132_);
  and (_20834_, _03087_, _02518_);
  nor (_20835_, _20834_, _02975_);
  nand (_20836_, _20835_, _20833_);
  and (_20837_, _08901_, _02975_);
  not (_20838_, _20837_);
  and (_20839_, _20838_, _09305_);
  nand (_20840_, _20839_, _20836_);
  nor (_20841_, _09305_, _02620_);
  nor (_20842_, _20841_, _02524_);
  and (_20844_, _20842_, _20840_);
  nor (_20845_, _08901_, _08824_);
  nor (_20846_, _20845_, _10325_);
  or (_20847_, _20846_, _20844_);
  and (_20848_, _08824_, _02608_);
  nor (_20849_, _20848_, _02894_);
  nand (_20850_, _20849_, _20847_);
  and (_20851_, _02894_, _02620_);
  nor (_20852_, _20851_, _02578_);
  nand (_20853_, _20852_, _20850_);
  and (_20855_, _03087_, _02578_);
  nor (_20856_, _20855_, _09318_);
  nand (_20857_, _20856_, _20853_);
  and (_20858_, _20695_, _09318_);
  nor (_20859_, _20858_, _05516_);
  and (_20860_, _20859_, _20857_);
  or (_20861_, _20860_, _20674_);
  nand (_20862_, _20861_, _05261_);
  and (_20863_, _08902_, _02974_);
  nor (_20864_, _20863_, _07807_);
  nand (_20866_, _20864_, _20862_);
  and (_20867_, _07807_, _02620_);
  nor (_20868_, _20867_, _09334_);
  nand (_20869_, _20868_, _20866_);
  and (_20870_, _09334_, _02632_);
  nor (_20871_, _20870_, _02893_);
  and (_20872_, _20871_, _20869_);
  and (_20873_, _02893_, _02620_);
  or (_20874_, _20873_, _02585_);
  or (_20875_, _20874_, _20872_);
  and (_20877_, _03087_, _02585_);
  nor (_20878_, _20877_, _09375_);
  nand (_20879_, _20878_, _20875_);
  and (_20880_, _08149_, _02620_);
  and (_20881_, _20695_, _09381_);
  or (_20882_, _20881_, _20880_);
  and (_20883_, _20882_, _09375_);
  nor (_20884_, _20883_, _09385_);
  and (_20885_, _20884_, _20879_);
  or (_20886_, _20885_, _20673_);
  nand (_20888_, _20886_, _08814_);
  nor (_20889_, _08814_, _02620_);
  nor (_20890_, _20889_, _02977_);
  and (_20891_, _20890_, _20888_);
  and (_20892_, _08901_, _02977_);
  or (_20893_, _20892_, _03107_);
  nor (_20894_, _20893_, _20891_);
  and (_20895_, _03107_, _02641_);
  or (_20896_, _20895_, _20894_);
  nand (_20897_, _20896_, _19652_);
  and (_20899_, _03087_, _02582_);
  nor (_20900_, _20899_, _09397_);
  nand (_20901_, _20900_, _20897_);
  nor (_20902_, _08149_, _02641_);
  and (_20903_, _20695_, _08149_);
  or (_20904_, _20903_, _20902_);
  and (_20905_, _20904_, _09397_);
  nor (_20906_, _20905_, _09406_);
  and (_20907_, _20906_, _20901_);
  or (_20908_, _20907_, _20672_);
  nand (_20910_, _20908_, _07881_);
  nor (_20911_, _07881_, _02620_);
  nor (_20912_, _20911_, _02991_);
  and (_20913_, _20912_, _20910_);
  and (_20914_, _08901_, _02991_);
  or (_20915_, _20914_, _03094_);
  nor (_20916_, _20915_, _20913_);
  and (_20917_, _03094_, _02641_);
  or (_20918_, _20917_, _20916_);
  nand (_20919_, _20918_, _10353_);
  and (_20921_, _03087_, _02594_);
  nor (_20922_, _20921_, _08807_);
  nand (_20923_, _20922_, _20919_);
  nor (_20924_, _20695_, \oc8051_golden_model_1.PSW [7]);
  nor (_20925_, _02620_, _07294_);
  nor (_20926_, _20925_, _08808_);
  not (_20927_, _20926_);
  nor (_20928_, _20927_, _20924_);
  nor (_20929_, _20928_, _09418_);
  and (_20930_, _20929_, _20923_);
  or (_20932_, _20930_, _20671_);
  nand (_20933_, _20932_, _07900_);
  nor (_20934_, _07900_, _02620_);
  nor (_20935_, _20934_, _02994_);
  and (_20936_, _20935_, _20933_);
  and (_20937_, _08901_, _02994_);
  or (_20938_, _20937_, _03099_);
  nor (_20939_, _20938_, _20936_);
  and (_20940_, _03099_, _02641_);
  or (_20941_, _20940_, _20939_);
  nand (_20943_, _20941_, _02590_);
  and (_20944_, _03087_, _02589_);
  nor (_20945_, _20944_, _08799_);
  nand (_20946_, _20945_, _20943_);
  nor (_20947_, _20695_, _07294_);
  nor (_20948_, _02620_, \oc8051_golden_model_1.PSW [7]);
  nor (_20949_, _20948_, _08800_);
  not (_20950_, _20949_);
  nor (_20951_, _20950_, _20947_);
  nor (_20952_, _20951_, _09434_);
  and (_20954_, _20952_, _20946_);
  or (_20955_, _20954_, _20670_);
  nand (_20956_, _20955_, _07947_);
  nor (_20957_, _07947_, _02620_);
  nor (_20958_, _20957_, _08027_);
  nand (_20959_, _20958_, _20956_);
  and (_20960_, _08027_, _02616_);
  nor (_20961_, _20960_, _03113_);
  and (_20962_, _20961_, _20959_);
  and (_20963_, _05935_, _03113_);
  or (_20965_, _20963_, _20962_);
  nand (_20966_, _20965_, _05741_);
  and (_20967_, _03087_, _02592_);
  nor (_20968_, _20967_, _02993_);
  nand (_20969_, _20968_, _20966_);
  and (_20970_, _20683_, _09640_);
  nor (_20971_, _09640_, _08901_);
  or (_20972_, _20971_, _03549_);
  or (_20973_, _20972_, _20970_);
  and (_20974_, _20973_, _08795_);
  and (_20976_, _20974_, _20969_);
  or (_20977_, _20976_, _20669_);
  nand (_20978_, _20977_, _20297_);
  and (_20979_, _08772_, _02641_);
  nor (_20980_, _20979_, _07143_);
  nand (_20981_, _20980_, _20978_);
  and (_20982_, _07143_, _02616_);
  nor (_20983_, _20982_, _02854_);
  and (_20984_, _20983_, _20981_);
  or (_20985_, _20984_, _20668_);
  nand (_20987_, _20985_, _19640_);
  and (_20988_, _03087_, _02575_);
  nor (_20989_, _20988_, _02990_);
  nand (_20990_, _20989_, _20987_);
  and (_20991_, _09640_, _08902_);
  nor (_20992_, _20682_, _09640_);
  nor (_20993_, _20992_, _20991_);
  and (_20994_, _20993_, _02990_);
  nor (_20995_, _20994_, _09668_);
  nand (_20996_, _20995_, _20990_);
  nor (_20998_, _09667_, _02616_);
  nor (_20999_, _20998_, _03133_);
  and (_21000_, _20999_, _20996_);
  or (_21001_, _21000_, _20666_);
  nand (_21002_, _21001_, _09675_);
  nor (_21003_, _09675_, _02608_);
  nor (_21004_, _21003_, _04331_);
  nand (_21005_, _21004_, _21002_);
  and (_21006_, _04331_, _03087_);
  nor (_21007_, _21006_, _02778_);
  nand (_21009_, _21007_, _21005_);
  and (_21010_, _20993_, _02778_);
  nor (_21011_, _21010_, _09689_);
  nand (_21012_, _21011_, _21009_);
  nor (_21013_, _09688_, _02616_);
  nor (_21014_, _21013_, _02852_);
  and (_21015_, _21014_, _21012_);
  and (_21016_, _09696_, _02641_);
  nor (_21017_, _21016_, _10371_);
  nor (_21018_, _21017_, _21015_);
  nor (_21020_, _09696_, _02616_);
  or (_21021_, _21020_, _21018_);
  nand (_21022_, _21021_, _10310_);
  and (_21023_, _19634_, _03087_);
  nor (_21024_, _21023_, _09706_);
  and (_21025_, _21024_, _21022_);
  and (_21026_, _09706_, _02616_);
  or (_21027_, _21026_, _21025_);
  or (_21028_, _21027_, _34450_);
  or (_21029_, _34446_, \oc8051_golden_model_1.PC [3]);
  and (_21031_, _21029_, _35583_);
  and (_35629_[3], _21031_, _21028_);
  and (_21032_, _19634_, _05581_);
  not (_21033_, _09696_);
  and (_21034_, _09089_, _02852_);
  or (_21035_, _21034_, _21033_);
  and (_21036_, _05581_, _04331_);
  not (_21037_, \oc8051_golden_model_1.PC [4]);
  nor (_21038_, _02212_, _21037_);
  and (_21039_, _02212_, _21037_);
  nor (_21041_, _21039_, _21038_);
  not (_21042_, _21041_);
  nor (_21043_, _21042_, _08812_);
  nor (_21044_, _09089_, _08149_);
  and (_21045_, _09109_, _09106_);
  nor (_21046_, _21045_, _09110_);
  and (_21047_, _21046_, _08149_);
  or (_21048_, _21047_, _21044_);
  and (_21049_, _21048_, _09397_);
  nor (_21050_, _21042_, _08822_);
  and (_21052_, _09088_, _08149_);
  and (_21053_, _21046_, _09381_);
  or (_21054_, _21053_, _21052_);
  and (_21055_, _21054_, _09375_);
  nor (_21056_, _09088_, _05267_);
  and (_21057_, _09089_, _02785_);
  nor (_21058_, _20048_, _09088_);
  and (_21059_, _21042_, _08827_);
  and (_21060_, _08898_, _08839_);
  and (_21061_, _08925_, _08922_);
  nor (_21063_, _21061_, _08926_);
  nor (_21064_, _21063_, _08839_);
  or (_21065_, _21064_, _08969_);
  nor (_21066_, _21065_, _21060_);
  nor (_21067_, _21066_, _08827_);
  and (_21068_, _09000_, _08897_);
  not (_21069_, _21063_);
  nor (_21070_, _21069_, _09000_);
  nor (_21071_, _21070_, _21068_);
  nor (_21072_, _21071_, _09858_);
  and (_21074_, _09089_, _02796_);
  nor (_21075_, _21041_, _09199_);
  nand (_21076_, _21046_, _09148_);
  or (_21077_, _09148_, _09089_);
  and (_21078_, _21077_, _21076_);
  and (_21079_, _21078_, _05327_);
  not (_21080_, _07425_);
  nor (_21081_, _05581_, _02546_);
  nor (_21082_, _21042_, _09165_);
  not (_21083_, _21082_);
  and (_21085_, _10364_, _09158_);
  and (_21086_, _09088_, _02837_);
  and (_21087_, _09168_, \oc8051_golden_model_1.PC [4]);
  nor (_21088_, _21087_, _21086_);
  nor (_21089_, _21088_, _20341_);
  and (_21090_, _21089_, _21085_);
  nor (_21091_, _21090_, _02934_);
  and (_21092_, _21091_, _21083_);
  not (_21093_, _21092_);
  nor (_21094_, _21093_, _21081_);
  and (_21096_, _09089_, _02934_);
  nor (_21097_, _21096_, _21094_);
  nor (_21098_, _21097_, _07428_);
  and (_21099_, _21042_, _07428_);
  nor (_21100_, _21099_, _21098_);
  and (_21101_, _21100_, _02544_);
  nor (_21102_, _05581_, _02544_);
  or (_21103_, _21102_, _21101_);
  and (_21104_, _21103_, _21080_);
  and (_21105_, _21041_, _07425_);
  nor (_21107_, _21105_, _05327_);
  not (_21108_, _21107_);
  nor (_21109_, _21108_, _21104_);
  or (_21110_, _21109_, _21079_);
  nand (_21111_, _21110_, _05311_);
  and (_21112_, _21042_, _03806_);
  nor (_21113_, _21112_, _02932_);
  nand (_21114_, _21113_, _21111_);
  or (_21115_, _09023_, _08898_);
  or (_21116_, _21069_, _09025_);
  nand (_21118_, _21116_, _21115_);
  nand (_21119_, _21118_, _02932_);
  nand (_21120_, _21119_, _21114_);
  nand (_21121_, _21120_, _09018_);
  nor (_21122_, _21042_, _09018_);
  nor (_21123_, _21122_, _02799_);
  nand (_21124_, _21123_, _21121_);
  and (_21125_, _09089_, _02799_);
  nor (_21126_, _21125_, _04239_);
  and (_21127_, _21126_, _21124_);
  nor (_21129_, _05581_, _02540_);
  or (_21130_, _21129_, _02930_);
  nor (_21131_, _21130_, _21127_);
  and (_21132_, _09089_, _02930_);
  or (_21133_, _21132_, _21131_);
  and (_21134_, _21133_, _09199_);
  or (_21135_, _21134_, _21075_);
  nand (_21136_, _21135_, _02943_);
  and (_21137_, _09089_, _02928_);
  nor (_21138_, _21137_, _09206_);
  nand (_21140_, _21138_, _21136_);
  and (_21141_, _21041_, _09206_);
  nor (_21142_, _21141_, _02796_);
  and (_21143_, _21142_, _21140_);
  or (_21144_, _21143_, _21074_);
  nand (_21145_, _21144_, _02538_);
  and (_21146_, _05581_, _09209_);
  nor (_21147_, _21146_, _02795_);
  nand (_21148_, _21147_, _21145_);
  and (_21149_, _09088_, _02795_);
  nor (_21151_, _21149_, _09906_);
  nand (_21152_, _21151_, _21148_);
  and (_21153_, _09252_, _08897_);
  nor (_21154_, _21069_, _09252_);
  or (_21155_, _21154_, _21153_);
  nor (_21156_, _21155_, _09217_);
  nor (_21157_, _21156_, _02972_);
  and (_21158_, _21157_, _21152_);
  or (_21159_, _21158_, _21072_);
  nand (_21160_, _21159_, _03397_);
  nand (_21162_, _09008_, _08897_);
  or (_21163_, _21069_, _09008_);
  and (_21164_, _21163_, _21162_);
  or (_21165_, _21164_, _03397_);
  nand (_21166_, _21165_, _21160_);
  nand (_21167_, _21166_, _08969_);
  and (_21168_, _21167_, _21067_);
  or (_21169_, _21168_, _21059_);
  nand (_21170_, _21169_, _06189_);
  and (_21171_, _09089_, _02790_);
  nor (_21173_, _21171_, _04230_);
  nand (_21174_, _21173_, _21170_);
  nor (_21175_, _05581_, _02533_);
  nor (_21176_, _21175_, _20432_);
  and (_21177_, _21176_, _21174_);
  or (_21178_, _21177_, _21058_);
  nand (_21179_, _21178_, _09273_);
  nor (_21180_, _21041_, _09273_);
  nor (_21181_, _21180_, _02902_);
  nand (_21182_, _21181_, _21179_);
  and (_21184_, _09088_, _02902_);
  nor (_21185_, _21184_, _09277_);
  nand (_21186_, _21185_, _21182_);
  and (_21187_, _05581_, _09277_);
  nor (_21188_, _21187_, _02901_);
  and (_21189_, _21188_, _21186_);
  and (_21190_, _09088_, _02901_);
  or (_21191_, _21190_, _21189_);
  nand (_21192_, _21191_, _09285_);
  nor (_21193_, _21042_, _09285_);
  nor (_21195_, _21193_, _09290_);
  nand (_21196_, _21195_, _21192_);
  nor (_21197_, _09289_, _09088_);
  nor (_21198_, _21197_, _07700_);
  nand (_21199_, _21198_, _21196_);
  nor (_21200_, _21042_, _02499_);
  nor (_21201_, _21200_, _02785_);
  and (_21202_, _21201_, _21199_);
  or (_21203_, _21202_, _21057_);
  nand (_21204_, _21203_, _04132_);
  and (_21206_, _05581_, _02518_);
  nor (_21207_, _21206_, _02975_);
  nand (_21208_, _21207_, _21204_);
  and (_21209_, _08897_, _02975_);
  not (_21210_, _21209_);
  and (_21211_, _21210_, _09305_);
  nand (_21212_, _21211_, _21208_);
  nor (_21213_, _09305_, _09088_);
  nor (_21214_, _21213_, _02524_);
  nand (_21215_, _21214_, _21212_);
  nor (_21217_, _08897_, _08824_);
  or (_21218_, _21217_, _10325_);
  nand (_21219_, _21218_, _21215_);
  and (_21220_, _21042_, _08824_);
  nor (_21221_, _21220_, _02894_);
  nand (_21222_, _21221_, _21219_);
  and (_21223_, _09088_, _02894_);
  nor (_21224_, _21223_, _02578_);
  nand (_21225_, _21224_, _21222_);
  and (_21226_, _05581_, _02578_);
  nor (_21228_, _21226_, _09318_);
  nand (_21229_, _21228_, _21225_);
  and (_21230_, _21046_, _09318_);
  nor (_21231_, _21230_, _05516_);
  and (_21232_, _21231_, _21229_);
  or (_21233_, _21232_, _21056_);
  nand (_21234_, _21233_, _05261_);
  and (_21235_, _08898_, _02974_);
  nor (_21236_, _21235_, _07807_);
  nand (_21237_, _21236_, _21234_);
  and (_21239_, _09088_, _07807_);
  nor (_21240_, _21239_, _09334_);
  nand (_21241_, _21240_, _21237_);
  and (_21242_, _09351_, _09348_);
  nor (_21243_, _21242_, _09352_);
  nor (_21244_, _21243_, _09335_);
  nor (_21245_, _21244_, _02893_);
  and (_21246_, _21245_, _21241_);
  and (_21247_, _09088_, _02893_);
  or (_21248_, _21247_, _02585_);
  or (_21250_, _21248_, _21246_);
  and (_21251_, _05581_, _02585_);
  nor (_21252_, _21251_, _09375_);
  and (_21253_, _21252_, _21250_);
  or (_21254_, _21253_, _21055_);
  and (_21255_, _21254_, _08822_);
  or (_21256_, _21255_, _08815_);
  or (_21257_, _21256_, _21050_);
  nor (_21258_, _08814_, _09088_);
  nor (_21259_, _21258_, _02977_);
  and (_21261_, _21259_, _21257_);
  and (_21262_, _08897_, _02977_);
  or (_21263_, _21262_, _03107_);
  nor (_21264_, _21263_, _21261_);
  and (_21265_, _09089_, _03107_);
  or (_21266_, _21265_, _21264_);
  nand (_21267_, _21266_, _19652_);
  and (_21268_, _05581_, _02582_);
  nor (_21269_, _21268_, _09397_);
  and (_21270_, _21269_, _21267_);
  or (_21272_, _21270_, _21049_);
  and (_21273_, _21272_, _08812_);
  or (_21274_, _21273_, _07882_);
  or (_21275_, _21274_, _21043_);
  nor (_21276_, _09088_, _07881_);
  nor (_21277_, _21276_, _02991_);
  and (_21278_, _21277_, _21275_);
  and (_21279_, _08897_, _02991_);
  or (_21280_, _21279_, _03094_);
  nor (_21281_, _21280_, _21278_);
  and (_21283_, _09089_, _03094_);
  or (_21284_, _21283_, _21281_);
  nand (_21285_, _21284_, _10353_);
  and (_21286_, _05581_, _02594_);
  nor (_21287_, _21286_, _08807_);
  nand (_21288_, _21287_, _21285_);
  nand (_21289_, _09088_, \oc8051_golden_model_1.PSW [7]);
  nand (_21290_, _21046_, _07294_);
  and (_21291_, _21290_, _21289_);
  or (_21292_, _21291_, _08808_);
  nand (_21294_, _21292_, _21288_);
  nand (_21295_, _21294_, _08805_);
  nor (_21296_, _21042_, _08805_);
  nor (_21297_, _21296_, _07901_);
  nand (_21298_, _21297_, _21295_);
  nor (_21299_, _09088_, _07900_);
  nor (_21300_, _21299_, _02994_);
  nand (_21301_, _21300_, _21298_);
  and (_21302_, _08897_, _02994_);
  nor (_21303_, _21302_, _03099_);
  and (_21304_, _21303_, _21301_);
  and (_21305_, _09089_, _03099_);
  or (_21306_, _21305_, _21304_);
  nand (_21307_, _21306_, _02590_);
  not (_21308_, _10376_);
  and (_21309_, _05581_, _02589_);
  nor (_21310_, _21309_, _21308_);
  nand (_21311_, _21310_, _21307_);
  nor (_21312_, _21046_, _07294_);
  nor (_21313_, _09088_, \oc8051_golden_model_1.PSW [7]);
  nor (_21315_, _21313_, _08800_);
  not (_21316_, _21315_);
  nor (_21317_, _21316_, _21312_);
  nor (_21318_, _21042_, _08797_);
  nor (_21319_, _21318_, _07948_);
  not (_21320_, _21319_);
  nor (_21321_, _21320_, _21317_);
  nand (_21322_, _21321_, _21311_);
  nor (_21323_, _09088_, _07947_);
  nor (_21324_, _21323_, _08027_);
  nand (_21326_, _21324_, _21322_);
  and (_21327_, _21041_, _08027_);
  nor (_21328_, _21327_, _03113_);
  and (_21329_, _21328_, _21326_);
  and (_21330_, _06072_, _03113_);
  or (_21331_, _21330_, _21329_);
  nand (_21332_, _21331_, _05741_);
  and (_21333_, _05581_, _02592_);
  nor (_21334_, _21333_, _02993_);
  and (_21335_, _21334_, _21332_);
  nor (_21337_, _09640_, _08898_);
  and (_21338_, _21063_, _09640_);
  nor (_21339_, _21338_, _21337_);
  nor (_21340_, _21339_, _03549_);
  or (_21341_, _21340_, _21335_);
  nand (_21342_, _21341_, _08795_);
  nor (_21343_, _21041_, _08772_);
  or (_21344_, _21343_, _10297_);
  nand (_21345_, _21344_, _21342_);
  and (_21346_, _09089_, _08772_);
  nor (_21348_, _21346_, _07143_);
  nand (_21349_, _21348_, _21345_);
  and (_21350_, _21041_, _07143_);
  nor (_21351_, _21350_, _02854_);
  nand (_21352_, _21351_, _21349_);
  and (_21353_, _06072_, _02854_);
  nor (_21354_, _21353_, _02575_);
  nand (_21355_, _21354_, _21352_);
  nor (_21356_, _05581_, _19640_);
  nor (_21357_, _21356_, _02990_);
  nand (_21359_, _21357_, _21355_);
  and (_21360_, _09640_, _08898_);
  nor (_21361_, _21063_, _09640_);
  nor (_21362_, _21361_, _21360_);
  nor (_21363_, _21362_, _03134_);
  nor (_21364_, _21363_, _09668_);
  nand (_21365_, _21364_, _21359_);
  nor (_21366_, _21042_, _09667_);
  nor (_21367_, _21366_, _03133_);
  nand (_21368_, _21367_, _21365_);
  not (_21371_, _09675_);
  and (_21372_, _09089_, _03133_);
  nor (_21373_, _21372_, _21371_);
  nand (_21374_, _21373_, _21368_);
  nor (_21375_, _21042_, _09675_);
  nor (_21376_, _21375_, _04331_);
  and (_21377_, _21376_, _21374_);
  or (_21378_, _21377_, _21036_);
  nand (_21379_, _21378_, _03142_);
  nor (_21380_, _21362_, _03142_);
  nor (_21382_, _21380_, _09689_);
  nand (_21383_, _21382_, _21379_);
  nor (_21384_, _21042_, _09688_);
  nor (_21385_, _21384_, _02852_);
  and (_21386_, _21385_, _21383_);
  or (_21387_, _21386_, _21035_);
  nor (_21388_, _21042_, _09696_);
  nor (_21389_, _21388_, _19634_);
  and (_21390_, _21389_, _21387_);
  or (_21391_, _21390_, _21032_);
  and (_21393_, _21391_, _09707_);
  and (_21394_, _21042_, _09706_);
  nor (_21395_, _21394_, _21393_);
  or (_21396_, _21395_, _34450_);
  or (_21397_, _34446_, \oc8051_golden_model_1.PC [4]);
  and (_21398_, _21397_, _35583_);
  and (_35629_[4], _21398_, _21396_);
  nor (_21399_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor (_21400_, _09083_, _02225_);
  nor (_21401_, _21400_, _21399_);
  nor (_21403_, _21401_, _09696_);
  and (_21404_, _09083_, _03133_);
  and (_21405_, _06027_, _02854_);
  nor (_21406_, _21401_, _08795_);
  nor (_21407_, _21401_, _08797_);
  nor (_21408_, _21401_, _08805_);
  nor (_21409_, _21401_, _08812_);
  nor (_21410_, _21401_, _08822_);
  nor (_21411_, _09083_, _05267_);
  and (_21412_, _09084_, _02785_);
  nor (_21414_, _20048_, _09083_);
  not (_21415_, _21401_);
  and (_21416_, _21415_, _08827_);
  and (_21417_, _09000_, _08892_);
  or (_21418_, _08894_, _08895_);
  and (_21419_, _21418_, _08927_);
  nor (_21420_, _21418_, _08927_);
  nor (_21421_, _21420_, _21419_);
  not (_21422_, _21421_);
  nor (_21423_, _21422_, _09000_);
  or (_21425_, _21423_, _21417_);
  nor (_21426_, _21425_, _09858_);
  and (_21427_, _21421_, _09023_);
  and (_21428_, _09025_, _08892_);
  or (_21429_, _21428_, _06162_);
  or (_21430_, _21429_, _21427_);
  or (_21431_, _09085_, _09086_);
  and (_21432_, _21431_, _09111_);
  nor (_21433_, _21431_, _09111_);
  nor (_21434_, _21433_, _21432_);
  and (_21436_, _21434_, _09148_);
  and (_21437_, _19690_, _09083_);
  nor (_21438_, _21437_, _21436_);
  nand (_21439_, _21438_, _05327_);
  nor (_21440_, _05612_, _02544_);
  and (_21441_, _09083_, _02934_);
  nor (_21442_, _05612_, _02546_);
  and (_21443_, _09168_, \oc8051_golden_model_1.PC [5]);
  and (_21444_, _09083_, _02837_);
  nor (_21445_, _21444_, _21443_);
  nor (_21447_, _21445_, _20341_);
  nor (_21448_, _21415_, _09164_);
  nor (_21449_, _21448_, _21447_);
  nor (_21450_, _21449_, _02804_);
  nor (_21451_, _21450_, _20340_);
  not (_21452_, _21451_);
  nor (_21453_, _21452_, _21442_);
  nor (_21454_, _21401_, _09159_);
  nor (_21455_, _21454_, _02934_);
  not (_21456_, _21455_);
  nor (_21458_, _21456_, _21453_);
  or (_21459_, _21458_, _07428_);
  nor (_21460_, _21459_, _21441_);
  and (_21461_, _21415_, _07428_);
  nor (_21462_, _21461_, _09178_);
  not (_21463_, _21462_);
  nor (_21464_, _21463_, _21460_);
  nor (_21465_, _21464_, _21440_);
  nor (_21466_, _21465_, _07425_);
  and (_21467_, _21401_, _07425_);
  nor (_21469_, _21467_, _05327_);
  not (_21470_, _21469_);
  nor (_21471_, _21470_, _21466_);
  nor (_21472_, _21471_, _03806_);
  and (_21473_, _21472_, _21439_);
  and (_21474_, _21401_, _03806_);
  or (_21475_, _21474_, _02932_);
  or (_21476_, _21475_, _21473_);
  nand (_21477_, _21476_, _21430_);
  nand (_21478_, _21477_, _09018_);
  nor (_21480_, _21401_, _09018_);
  nor (_21481_, _21480_, _02799_);
  and (_21482_, _21481_, _21478_);
  and (_21483_, _09083_, _02799_);
  or (_21484_, _21483_, _04239_);
  or (_21485_, _21484_, _21482_);
  and (_21486_, _05612_, _04239_);
  nor (_21487_, _21486_, _02930_);
  nand (_21488_, _21487_, _21485_);
  and (_21489_, _09083_, _02930_);
  nor (_21491_, _21489_, _09200_);
  nand (_21492_, _21491_, _21488_);
  nor (_21493_, _21401_, _09199_);
  nor (_21494_, _21493_, _02928_);
  nand (_21495_, _21494_, _21492_);
  and (_21496_, _09083_, _02928_);
  nor (_21497_, _21496_, _09206_);
  nand (_21498_, _21497_, _21495_);
  and (_21499_, _21415_, _09206_);
  nor (_21500_, _21499_, _02796_);
  nand (_21502_, _21500_, _21498_);
  and (_21503_, _09083_, _02796_);
  nor (_21504_, _21503_, _09209_);
  nand (_21505_, _21504_, _21502_);
  and (_21506_, _05612_, _09209_);
  nor (_21507_, _21506_, _02795_);
  nand (_21508_, _21507_, _21505_);
  and (_21509_, _09083_, _02795_);
  nor (_21510_, _21509_, _09906_);
  and (_21511_, _21510_, _21508_);
  and (_21513_, _09252_, _08892_);
  nor (_21514_, _21422_, _09252_);
  or (_21515_, _21514_, _21513_);
  nor (_21516_, _21515_, _09217_);
  or (_21517_, _21516_, _21511_);
  and (_21518_, _21517_, _09858_);
  or (_21519_, _21518_, _21426_);
  or (_21520_, _21519_, _02944_);
  and (_21521_, _09008_, _08892_);
  nor (_21522_, _21422_, _09008_);
  nor (_21524_, _21522_, _21521_);
  or (_21525_, _21524_, _03397_);
  and (_21526_, _21525_, _21520_);
  or (_21527_, _21526_, _02979_);
  and (_21528_, _08893_, _08839_);
  nor (_21529_, _21421_, _08839_);
  or (_21530_, _21529_, _08969_);
  nor (_21531_, _21530_, _21528_);
  nor (_21532_, _21531_, _08827_);
  and (_21533_, _21532_, _21527_);
  or (_21535_, _21533_, _21416_);
  nand (_21536_, _21535_, _06189_);
  and (_21537_, _09084_, _02790_);
  nor (_21538_, _21537_, _04230_);
  nand (_21539_, _21538_, _21536_);
  nor (_21540_, _05612_, _02533_);
  nor (_21541_, _21540_, _20432_);
  and (_21542_, _21541_, _21539_);
  or (_21543_, _21542_, _21414_);
  nand (_21544_, _21543_, _09273_);
  nor (_21546_, _21401_, _09273_);
  nor (_21547_, _21546_, _02902_);
  nand (_21548_, _21547_, _21544_);
  and (_21549_, _09083_, _02902_);
  nor (_21550_, _21549_, _09277_);
  nand (_21551_, _21550_, _21548_);
  and (_21552_, _05612_, _09277_);
  nor (_21553_, _21552_, _02901_);
  nand (_21554_, _21553_, _21551_);
  and (_21555_, _09083_, _02901_);
  nor (_21557_, _21555_, _20447_);
  and (_21558_, _21557_, _21554_);
  nor (_21559_, _21401_, _09285_);
  or (_21560_, _21559_, _21558_);
  nand (_21561_, _21560_, _09289_);
  nor (_21562_, _09289_, _09083_);
  nor (_21563_, _21562_, _07700_);
  nand (_21564_, _21563_, _21561_);
  nor (_21565_, _21415_, _02499_);
  nor (_21566_, _21565_, _02785_);
  and (_21568_, _21566_, _21564_);
  or (_21569_, _21568_, _21412_);
  nand (_21570_, _21569_, _04132_);
  and (_21571_, _05612_, _02518_);
  nor (_21572_, _21571_, _02975_);
  nand (_21573_, _21572_, _21570_);
  and (_21574_, _08892_, _02975_);
  not (_21575_, _21574_);
  and (_21576_, _21575_, _09305_);
  nand (_21577_, _21576_, _21573_);
  nor (_21579_, _09305_, _09083_);
  nor (_21580_, _21579_, _02524_);
  and (_21581_, _21580_, _21577_);
  nor (_21582_, _08892_, _08824_);
  nor (_21583_, _21582_, _10325_);
  or (_21584_, _21583_, _21581_);
  and (_21585_, _21415_, _08824_);
  nor (_21586_, _21585_, _02894_);
  nand (_21587_, _21586_, _21584_);
  nor (_21588_, _09083_, _02578_);
  or (_21590_, _21588_, _09315_);
  nand (_21591_, _21590_, _21587_);
  and (_21592_, _05612_, _02578_);
  nor (_21593_, _21592_, _09318_);
  nand (_21594_, _21593_, _21591_);
  and (_21595_, _21434_, _09318_);
  nor (_21596_, _21595_, _05516_);
  and (_21597_, _21596_, _21594_);
  or (_21598_, _21597_, _21411_);
  nand (_21599_, _21598_, _05261_);
  and (_21601_, _08893_, _02974_);
  nor (_21602_, _21601_, _07807_);
  nand (_21603_, _21602_, _21599_);
  and (_21604_, _09083_, _07807_);
  nor (_21605_, _21604_, _09334_);
  nand (_21606_, _21605_, _21603_);
  or (_21607_, _09345_, _09346_);
  and (_21608_, _21607_, _09353_);
  nor (_21609_, _21607_, _09353_);
  nor (_21610_, _21609_, _21608_);
  nor (_21612_, _21610_, _09335_);
  nor (_21613_, _21612_, _02893_);
  nand (_21614_, _21613_, _21606_);
  and (_21615_, _09083_, _02893_);
  nor (_21616_, _21615_, _02585_);
  nand (_21617_, _21616_, _21614_);
  and (_21618_, _05612_, _02585_);
  nor (_21619_, _21618_, _09375_);
  nand (_21620_, _21619_, _21617_);
  and (_21621_, _09083_, _08149_);
  and (_21623_, _21434_, _09381_);
  or (_21624_, _21623_, _21621_);
  and (_21625_, _21624_, _09375_);
  nor (_21626_, _21625_, _09385_);
  and (_21627_, _21626_, _21620_);
  or (_21628_, _21627_, _21410_);
  nand (_21629_, _21628_, _08814_);
  nor (_21630_, _08814_, _09083_);
  nor (_21631_, _21630_, _02977_);
  and (_21632_, _21631_, _21629_);
  and (_21634_, _08892_, _02977_);
  or (_21635_, _21634_, _03107_);
  nor (_21636_, _21635_, _21632_);
  and (_21637_, _09084_, _03107_);
  or (_21638_, _21637_, _21636_);
  nand (_21639_, _21638_, _19652_);
  and (_21640_, _05612_, _02582_);
  nor (_21641_, _21640_, _09397_);
  nand (_21642_, _21641_, _21639_);
  or (_21643_, _21434_, _09381_);
  or (_21645_, _09083_, _08149_);
  and (_21646_, _21645_, _09397_);
  and (_21647_, _21646_, _21643_);
  nor (_21648_, _21647_, _09406_);
  and (_21649_, _21648_, _21642_);
  or (_21650_, _21649_, _21409_);
  nand (_21651_, _21650_, _07881_);
  nor (_21652_, _09083_, _07881_);
  nor (_21653_, _21652_, _02991_);
  and (_21654_, _21653_, _21651_);
  and (_21656_, _08892_, _02991_);
  or (_21657_, _21656_, _03094_);
  nor (_21658_, _21657_, _21654_);
  and (_21659_, _09084_, _03094_);
  or (_21660_, _21659_, _21658_);
  nand (_21661_, _21660_, _10353_);
  and (_21662_, _05612_, _02594_);
  nor (_21663_, _21662_, _08807_);
  nand (_21664_, _21663_, _21661_);
  nor (_21665_, _21434_, \oc8051_golden_model_1.PSW [7]);
  nor (_21667_, _09083_, _07294_);
  nor (_21668_, _21667_, _08808_);
  not (_21669_, _21668_);
  nor (_21670_, _21669_, _21665_);
  nor (_21671_, _21670_, _09418_);
  and (_21672_, _21671_, _21664_);
  or (_21673_, _21672_, _21408_);
  nand (_21674_, _21673_, _07900_);
  nor (_21675_, _09083_, _07900_);
  nor (_21676_, _21675_, _02994_);
  and (_21678_, _21676_, _21674_);
  and (_21679_, _08892_, _02994_);
  or (_21680_, _21679_, _03099_);
  nor (_21681_, _21680_, _21678_);
  and (_21682_, _09084_, _03099_);
  or (_21683_, _21682_, _21681_);
  nand (_21684_, _21683_, _02590_);
  and (_21685_, _05612_, _02589_);
  nor (_21686_, _21685_, _08799_);
  nand (_21687_, _21686_, _21684_);
  and (_21689_, _09083_, _07294_);
  and (_21690_, _21434_, \oc8051_golden_model_1.PSW [7]);
  or (_21691_, _21690_, _21689_);
  and (_21692_, _21691_, _08799_);
  nor (_21693_, _21692_, _09434_);
  and (_21694_, _21693_, _21687_);
  or (_21695_, _21694_, _21407_);
  nand (_21696_, _21695_, _07947_);
  nor (_21697_, _09083_, _07947_);
  nor (_21698_, _21697_, _08027_);
  nand (_21700_, _21698_, _21696_);
  and (_21701_, _21401_, _08027_);
  nor (_21702_, _21701_, _03113_);
  and (_21703_, _21702_, _21700_);
  and (_21704_, _06027_, _03113_);
  or (_21705_, _21704_, _21703_);
  nand (_21706_, _21705_, _05741_);
  and (_21707_, _05612_, _02592_);
  nor (_21708_, _21707_, _02993_);
  nand (_21709_, _21708_, _21706_);
  nor (_21711_, _09640_, _08892_);
  and (_21712_, _21422_, _09640_);
  or (_21713_, _21712_, _03549_);
  or (_21714_, _21713_, _21711_);
  and (_21715_, _21714_, _08795_);
  and (_21716_, _21715_, _21709_);
  or (_21717_, _21716_, _21406_);
  nand (_21718_, _21717_, _20297_);
  and (_21719_, _09084_, _08772_);
  nor (_21720_, _21719_, _07143_);
  nand (_21722_, _21720_, _21718_);
  and (_21723_, _21401_, _07143_);
  nor (_21724_, _21723_, _02854_);
  and (_21725_, _21724_, _21722_);
  or (_21726_, _21725_, _21405_);
  nand (_21727_, _21726_, _19640_);
  and (_21728_, _05612_, _02575_);
  nor (_21729_, _21728_, _02990_);
  nand (_21730_, _21729_, _21727_);
  nor (_21731_, _21421_, _09640_);
  and (_21733_, _09640_, _08893_);
  nor (_21734_, _21733_, _21731_);
  and (_21735_, _21734_, _02990_);
  nor (_21736_, _21735_, _09668_);
  nand (_21737_, _21736_, _21730_);
  nor (_21738_, _21401_, _09667_);
  nor (_21739_, _21738_, _03133_);
  and (_21740_, _21739_, _21737_);
  or (_21741_, _21740_, _21404_);
  nand (_21742_, _21741_, _09675_);
  nor (_21744_, _21415_, _09675_);
  nor (_21745_, _21744_, _04331_);
  nand (_21746_, _21745_, _21742_);
  and (_21747_, _05612_, _04331_);
  nor (_21748_, _21747_, _02778_);
  nand (_21749_, _21748_, _21746_);
  and (_21750_, _21734_, _02778_);
  nor (_21751_, _21750_, _09689_);
  nand (_21752_, _21751_, _21749_);
  nor (_21753_, _21401_, _09688_);
  nor (_21755_, _21753_, _02852_);
  nand (_21756_, _21755_, _21752_);
  and (_21757_, _09083_, _02852_);
  nor (_21758_, _21757_, _21033_);
  and (_21759_, _21758_, _21756_);
  or (_21760_, _21759_, _21403_);
  nand (_21761_, _21760_, _10310_);
  and (_21762_, _19634_, _05612_);
  nor (_21763_, _21762_, _09706_);
  and (_21764_, _21763_, _21761_);
  and (_21766_, _21401_, _09706_);
  or (_21767_, _21766_, _21764_);
  or (_21768_, _21767_, _34450_);
  or (_21769_, _34446_, \oc8051_golden_model_1.PC [5]);
  and (_21770_, _21769_, _35583_);
  and (_35629_[5], _21770_, _21768_);
  and (_21771_, _19634_, _05549_);
  and (_21772_, _05313_, _08774_);
  nor (_21773_, _21772_, \oc8051_golden_model_1.PC [6]);
  nor (_21774_, _21773_, _08775_);
  not (_21776_, _21774_);
  nor (_21777_, _21776_, _09696_);
  and (_21778_, _09077_, _02852_);
  or (_21779_, _21778_, _21033_);
  and (_21780_, _05549_, _04331_);
  and (_21781_, _21776_, _07143_);
  nor (_21782_, _09076_, _07900_);
  or (_21783_, _09076_, _05267_);
  nand (_21784_, _09077_, _02894_);
  or (_21785_, _21774_, _02499_);
  nand (_21787_, _21776_, _08827_);
  and (_21788_, _09252_, _08885_);
  nor (_21789_, _08929_, _08889_);
  nor (_21790_, _21789_, _08930_);
  not (_21791_, _21790_);
  nor (_21792_, _21791_, _09252_);
  or (_21793_, _21792_, _21788_);
  or (_21794_, _21793_, _09217_);
  nand (_21795_, _09077_, _02796_);
  or (_21796_, _21774_, _09199_);
  nand (_21798_, _21776_, _03806_);
  and (_21799_, _21798_, _06162_);
  and (_21800_, _09150_, _09076_);
  nor (_21801_, _09113_, _09080_);
  nor (_21802_, _21801_, _09114_);
  and (_21803_, _21802_, _09148_);
  or (_21804_, _21803_, _21800_);
  or (_21805_, _21804_, _05325_);
  nand (_21806_, _05549_, _02804_);
  and (_21807_, _09076_, _02837_);
  and (_21809_, _09168_, \oc8051_golden_model_1.PC [6]);
  or (_21810_, _21809_, _21807_);
  and (_21811_, _21810_, _09163_);
  nor (_21812_, _21776_, _09164_);
  or (_21813_, _21812_, _21811_);
  and (_21814_, _21813_, _09159_);
  or (_21815_, _21814_, _02804_);
  and (_21816_, _21815_, _21806_);
  nor (_21817_, _21776_, _09159_);
  or (_21818_, _21817_, _02934_);
  or (_21820_, _21818_, _21816_);
  and (_21821_, _09077_, _02934_);
  nor (_21822_, _21821_, _07428_);
  and (_21823_, _21822_, _21820_);
  and (_21824_, _21774_, _07428_);
  or (_21825_, _21824_, _09178_);
  or (_21826_, _21825_, _21823_);
  nand (_21827_, _05549_, _09178_);
  and (_21828_, _21827_, _21080_);
  and (_21829_, _21828_, _21826_);
  nand (_21831_, _21774_, _07425_);
  nand (_21832_, _21831_, _05325_);
  or (_21833_, _21832_, _21829_);
  and (_21834_, _21833_, _21805_);
  or (_21835_, _21834_, _03806_);
  and (_21836_, _21835_, _21799_);
  and (_21837_, _09025_, _08885_);
  and (_21838_, _21790_, _09023_);
  or (_21839_, _21838_, _21837_);
  and (_21840_, _21839_, _02932_);
  or (_21842_, _21840_, _21836_);
  and (_21843_, _21842_, _09018_);
  nor (_21844_, _21776_, _09018_);
  or (_21845_, _21844_, _02799_);
  or (_21846_, _21845_, _21843_);
  nand (_21847_, _09077_, _02799_);
  and (_21848_, _21847_, _02540_);
  and (_21849_, _21848_, _21846_);
  nor (_21850_, _05549_, _02540_);
  or (_21851_, _21850_, _02930_);
  or (_21853_, _21851_, _21849_);
  nand (_21854_, _09077_, _02930_);
  and (_21855_, _21854_, _21853_);
  or (_21856_, _21855_, _09200_);
  and (_21857_, _21856_, _21796_);
  or (_21858_, _21857_, _02928_);
  and (_21859_, _09077_, _02928_);
  nor (_21860_, _21859_, _09206_);
  and (_21861_, _21860_, _21858_);
  and (_21862_, _21774_, _09206_);
  or (_21864_, _21862_, _02796_);
  or (_21865_, _21864_, _21861_);
  and (_21866_, _21865_, _21795_);
  or (_21867_, _21866_, _09209_);
  nand (_21868_, _05549_, _09209_);
  and (_21869_, _21868_, _03932_);
  and (_21870_, _21869_, _21867_);
  nand (_21871_, _09076_, _02795_);
  nand (_21872_, _21871_, _09217_);
  or (_21873_, _21872_, _21870_);
  and (_21874_, _21873_, _21794_);
  or (_21875_, _21874_, _02972_);
  and (_21876_, _09000_, _08885_);
  nor (_21877_, _21791_, _09000_);
  or (_21878_, _21877_, _09858_);
  or (_21879_, _21878_, _21876_);
  and (_21880_, _21879_, _03397_);
  and (_21881_, _21880_, _21875_);
  nor (_21882_, _21791_, _09008_);
  and (_21883_, _09008_, _08885_);
  or (_21886_, _21883_, _21882_);
  and (_21887_, _21886_, _02944_);
  or (_21888_, _21887_, _21881_);
  and (_21889_, _21888_, _08969_);
  or (_21890_, _21790_, _08839_);
  nand (_21891_, _08886_, _08839_);
  and (_21892_, _21891_, _02979_);
  and (_21893_, _21892_, _21890_);
  or (_21894_, _21893_, _08827_);
  or (_21895_, _21894_, _21889_);
  and (_21897_, _21895_, _21787_);
  or (_21898_, _21897_, _02790_);
  nand (_21899_, _09077_, _02790_);
  and (_21900_, _21899_, _02533_);
  and (_21901_, _21900_, _21898_);
  nor (_21902_, _05549_, _02533_);
  or (_21903_, _21902_, _20432_);
  or (_21904_, _21903_, _21901_);
  or (_21905_, _20048_, _09076_);
  and (_21906_, _21905_, _21904_);
  or (_21908_, _21906_, _09281_);
  or (_21909_, _21774_, _09273_);
  and (_21910_, _21909_, _09276_);
  and (_21911_, _21910_, _21908_);
  and (_21912_, _09076_, _02902_);
  or (_21913_, _21912_, _09277_);
  or (_21914_, _21913_, _21911_);
  nand (_21915_, _05549_, _09277_);
  and (_21916_, _21915_, _09759_);
  and (_21917_, _21916_, _21914_);
  nand (_21919_, _09076_, _02901_);
  nand (_21920_, _21919_, _09285_);
  or (_21921_, _21920_, _21917_);
  or (_21922_, _21774_, _09285_);
  and (_21923_, _21922_, _09289_);
  and (_21924_, _21923_, _21921_);
  nor (_21925_, _09289_, _09077_);
  or (_21926_, _21925_, _07700_);
  or (_21927_, _21926_, _21924_);
  and (_21928_, _21927_, _21785_);
  or (_21930_, _21928_, _02785_);
  nand (_21931_, _09077_, _02785_);
  and (_21932_, _21931_, _04132_);
  and (_21933_, _21932_, _21930_);
  nor (_21934_, _05549_, _04132_);
  or (_21935_, _21934_, _02975_);
  or (_21936_, _21935_, _21933_);
  nand (_21937_, _08886_, _02975_);
  and (_21938_, _21937_, _09305_);
  and (_21939_, _21938_, _21936_);
  nor (_21941_, _09305_, _09077_);
  or (_21942_, _21941_, _02524_);
  or (_21943_, _21942_, _21939_);
  nor (_21944_, _08886_, _08824_);
  or (_21945_, _21944_, _10325_);
  and (_21946_, _21945_, _21943_);
  and (_21947_, _21774_, _08824_);
  or (_21948_, _21947_, _02894_);
  or (_21949_, _21948_, _21946_);
  and (_21950_, _21949_, _21784_);
  or (_21952_, _21950_, _02578_);
  nand (_21953_, _05549_, _02578_);
  and (_21954_, _21953_, _09319_);
  and (_21955_, _21954_, _21952_);
  and (_21956_, _21802_, _09318_);
  or (_21957_, _21956_, _05516_);
  or (_21958_, _21957_, _21955_);
  and (_21959_, _21958_, _21783_);
  or (_21960_, _21959_, _02974_);
  nand (_21961_, _08886_, _02974_);
  and (_21963_, _21961_, _07808_);
  and (_21964_, _21963_, _21960_);
  and (_21965_, _09076_, _07807_);
  or (_21966_, _21965_, _09334_);
  or (_21967_, _21966_, _21964_);
  nor (_21968_, _09355_, _09344_);
  nor (_21969_, _21968_, _09356_);
  or (_21970_, _21969_, _09335_);
  and (_21971_, _21970_, _10067_);
  and (_21972_, _21971_, _21967_);
  and (_21974_, _09076_, _02893_);
  or (_21975_, _21974_, _02585_);
  or (_21976_, _21975_, _21972_);
  nand (_21977_, _05549_, _02585_);
  and (_21978_, _21977_, _10350_);
  and (_21979_, _21978_, _21976_);
  or (_21980_, _21802_, _08149_);
  or (_21981_, _09076_, _09381_);
  and (_21982_, _21981_, _09375_);
  and (_21983_, _21982_, _21980_);
  nor (_21985_, _21776_, _08822_);
  or (_21986_, _21985_, _21983_);
  or (_21987_, _21986_, _21979_);
  and (_21988_, _21987_, _08814_);
  nor (_21989_, _08814_, _09077_);
  or (_21990_, _21989_, _02977_);
  or (_21991_, _21990_, _21988_);
  nand (_21992_, _08886_, _02977_);
  and (_21993_, _21992_, _07104_);
  and (_21994_, _21993_, _21991_);
  and (_21996_, _09076_, _03107_);
  or (_21997_, _21996_, _02582_);
  or (_21998_, _21997_, _21994_);
  nand (_21999_, _05549_, _02582_);
  and (_22000_, _21999_, _10355_);
  nand (_22001_, _22000_, _21998_);
  or (_22002_, _21802_, _09381_);
  or (_22003_, _09076_, _08149_);
  and (_22004_, _22003_, _09397_);
  and (_22005_, _22004_, _22002_);
  nor (_22007_, _21776_, _08812_);
  or (_22008_, _22007_, _07882_);
  nor (_22009_, _22008_, _22005_);
  and (_22010_, _22009_, _22001_);
  nor (_22011_, _09076_, _07881_);
  or (_22012_, _22011_, _22010_);
  and (_22013_, _22012_, _03881_);
  and (_22014_, _08886_, _02991_);
  or (_22015_, _22014_, _03094_);
  or (_22016_, _22015_, _22013_);
  nand (_22018_, _09076_, _03094_);
  and (_22019_, _22018_, _10353_);
  and (_22020_, _22019_, _22016_);
  nand (_22021_, _05549_, _02594_);
  nand (_22022_, _22021_, _10379_);
  or (_22023_, _22022_, _22020_);
  nor (_22024_, _21802_, \oc8051_golden_model_1.PSW [7]);
  or (_22025_, _09076_, _07294_);
  nand (_22026_, _22025_, _08807_);
  or (_22027_, _22026_, _22024_);
  or (_22029_, _21776_, _08805_);
  and (_22030_, _22029_, _07900_);
  and (_22031_, _22030_, _22027_);
  and (_22032_, _22031_, _22023_);
  or (_22033_, _22032_, _21782_);
  and (_22034_, _22033_, _07120_);
  and (_22035_, _08886_, _02994_);
  or (_22036_, _22035_, _03099_);
  or (_22037_, _22036_, _22034_);
  nand (_22038_, _09076_, _03099_);
  and (_22040_, _22038_, _02590_);
  and (_22041_, _22040_, _22037_);
  and (_22042_, _05549_, _02589_);
  or (_22043_, _22042_, _21308_);
  or (_22044_, _22043_, _22041_);
  nor (_22045_, _21802_, _07294_);
  or (_22046_, _09076_, \oc8051_golden_model_1.PSW [7]);
  nand (_22047_, _22046_, _08799_);
  or (_22048_, _22047_, _22045_);
  or (_22049_, _21776_, _08797_);
  and (_22051_, _22049_, _07947_);
  and (_22052_, _22051_, _22048_);
  and (_22053_, _22052_, _22044_);
  nor (_22054_, _09076_, _07947_);
  or (_22055_, _22054_, _08027_);
  or (_22056_, _22055_, _22053_);
  nand (_22057_, _21774_, _08027_);
  and (_22058_, _22057_, _22056_);
  or (_22059_, _22058_, _03113_);
  nand (_22060_, _05798_, _03113_);
  and (_22062_, _22060_, _05741_);
  and (_22063_, _22062_, _22059_);
  and (_22064_, _05549_, _02592_);
  or (_22065_, _22064_, _02993_);
  or (_22066_, _22065_, _22063_);
  nor (_22067_, _09640_, _08885_);
  and (_22068_, _21791_, _09640_);
  or (_22069_, _22068_, _03549_);
  or (_22070_, _22069_, _22067_);
  and (_22071_, _22070_, _08795_);
  and (_22073_, _22071_, _22066_);
  nor (_22074_, _21776_, _08772_);
  nor (_22075_, _22074_, _10297_);
  or (_22076_, _22075_, _22073_);
  nand (_22077_, _09076_, _08772_);
  and (_22078_, _22077_, _09650_);
  and (_22079_, _22078_, _22076_);
  or (_22080_, _22079_, _21781_);
  and (_22081_, _22080_, _02855_);
  nor (_22082_, _05798_, _02855_);
  or (_22084_, _22082_, _02575_);
  or (_22085_, _22084_, _22081_);
  or (_22086_, _05549_, _19640_);
  and (_22087_, _22086_, _03134_);
  and (_22088_, _22087_, _22085_);
  and (_22089_, _09640_, _08886_);
  nor (_22090_, _21790_, _09640_);
  or (_22091_, _22090_, _22089_);
  and (_22092_, _22091_, _02990_);
  or (_22093_, _22092_, _22088_);
  and (_22095_, _22093_, _09667_);
  nor (_22096_, _21774_, _09667_);
  or (_22097_, _22096_, _22095_);
  and (_22098_, _22097_, _03138_);
  nand (_22099_, _09077_, _03133_);
  nand (_22100_, _22099_, _09675_);
  or (_22101_, _22100_, _22098_);
  or (_22102_, _21776_, _09675_);
  and (_22103_, _22102_, _03907_);
  and (_22104_, _22103_, _22101_);
  or (_22106_, _22104_, _21780_);
  and (_22107_, _22106_, _03142_);
  and (_22108_, _22091_, _02778_);
  or (_22109_, _22108_, _09689_);
  nor (_22110_, _22109_, _22107_);
  nor (_22111_, _21776_, _09688_);
  nor (_22112_, _22111_, _02852_);
  not (_22113_, _22112_);
  nor (_22114_, _22113_, _22110_);
  nor (_22115_, _22114_, _21779_);
  or (_22117_, _22115_, _19634_);
  nor (_22118_, _22117_, _21777_);
  nor (_22119_, _22118_, _21771_);
  nor (_22120_, _22119_, _09706_);
  and (_22121_, _21776_, _09706_);
  nor (_22122_, _22121_, _22120_);
  or (_22123_, _22122_, _34450_);
  or (_22124_, _34446_, \oc8051_golden_model_1.PC [6]);
  and (_22125_, _22124_, _35583_);
  and (_35629_[6], _22125_, _22123_);
  and (_22127_, _05318_, _03133_);
  nor (_22128_, _08775_, \oc8051_golden_model_1.PC [7]);
  nor (_22129_, _22128_, _08776_);
  nor (_22130_, _22129_, _08795_);
  nor (_22131_, _22129_, _08797_);
  nor (_22132_, _22129_, _08805_);
  nor (_22133_, _22129_, _08812_);
  nor (_22134_, _22129_, _08822_);
  nor (_22135_, _05318_, _05267_);
  nor (_22136_, _22129_, _09285_);
  nor (_22137_, _20048_, _05318_);
  not (_22138_, _22129_);
  and (_22139_, _22138_, _08827_);
  and (_22140_, _08839_, _06098_);
  not (_22141_, _08839_);
  and (_22142_, _08931_, _08882_);
  nor (_22143_, _22142_, _08932_);
  and (_22144_, _22143_, _22141_);
  nor (_22145_, _22144_, _22140_);
  nor (_22146_, _22145_, _08969_);
  nor (_22149_, _22146_, _08827_);
  or (_22150_, _09023_, _06098_);
  or (_22151_, _22143_, _09025_);
  and (_22152_, _22151_, _22150_);
  or (_22153_, _22152_, _06162_);
  and (_22154_, _09115_, _09073_);
  nor (_22155_, _22154_, _09116_);
  and (_22156_, _22155_, _09148_);
  and (_22157_, _19690_, _05318_);
  nor (_22158_, _22157_, _22156_);
  nand (_22160_, _22158_, _05327_);
  and (_22161_, _22138_, _07428_);
  and (_22162_, _05318_, _02934_);
  nor (_22163_, _05256_, _02546_);
  and (_22164_, _09168_, \oc8051_golden_model_1.PC [7]);
  and (_22165_, _05318_, _02837_);
  nor (_22166_, _22165_, _22164_);
  nor (_22167_, _22166_, _20341_);
  nor (_22168_, _22138_, _09164_);
  nor (_22169_, _22168_, _22167_);
  nor (_22171_, _22169_, _02804_);
  nor (_22172_, _22171_, _20340_);
  not (_22173_, _22172_);
  nor (_22174_, _22173_, _22163_);
  nor (_22175_, _22129_, _09159_);
  nor (_22176_, _22175_, _02934_);
  not (_22177_, _22176_);
  nor (_22178_, _22177_, _22174_);
  or (_22179_, _22178_, _07428_);
  nor (_22180_, _22179_, _22162_);
  or (_22182_, _22180_, _09178_);
  nor (_22183_, _22182_, _22161_);
  nor (_22184_, _05256_, _02544_);
  nor (_22185_, _22184_, _22183_);
  nor (_22186_, _22185_, _07425_);
  and (_22187_, _22129_, _07425_);
  nor (_22188_, _22187_, _05327_);
  not (_22189_, _22188_);
  nor (_22190_, _22189_, _22186_);
  nor (_22191_, _22190_, _03806_);
  and (_22193_, _22191_, _22160_);
  and (_22194_, _22129_, _03806_);
  or (_22195_, _22194_, _02932_);
  or (_22196_, _22195_, _22193_);
  nand (_22197_, _22196_, _22153_);
  nand (_22198_, _22197_, _09018_);
  nor (_22199_, _22129_, _09018_);
  nor (_22200_, _22199_, _02799_);
  and (_22201_, _22200_, _22198_);
  and (_22202_, _05318_, _02799_);
  or (_22204_, _22202_, _04239_);
  or (_22205_, _22204_, _22201_);
  and (_22206_, _05256_, _04239_);
  nor (_22207_, _22206_, _02930_);
  nand (_22208_, _22207_, _22205_);
  and (_22209_, _05318_, _02930_);
  nor (_22210_, _22209_, _09200_);
  nand (_22211_, _22210_, _22208_);
  nor (_22212_, _22129_, _09199_);
  nor (_22213_, _22212_, _02928_);
  nand (_22215_, _22213_, _22211_);
  and (_22216_, _05318_, _02928_);
  nor (_22217_, _22216_, _09206_);
  nand (_22218_, _22217_, _22215_);
  and (_22219_, _22138_, _09206_);
  nor (_22220_, _22219_, _02796_);
  and (_22221_, _22220_, _22218_);
  and (_22222_, _05318_, _02796_);
  or (_22223_, _22222_, _09209_);
  or (_22224_, _22223_, _22221_);
  and (_22226_, _05256_, _09209_);
  nor (_22227_, _22226_, _02795_);
  nand (_22228_, _22227_, _22224_);
  and (_22229_, _05318_, _02795_);
  nor (_22230_, _22229_, _09906_);
  and (_22231_, _22230_, _22228_);
  and (_22232_, _09252_, _06098_);
  not (_22233_, _22143_);
  nor (_22234_, _22233_, _09252_);
  or (_22235_, _22234_, _22232_);
  nor (_22237_, _22235_, _09217_);
  or (_22238_, _22237_, _22231_);
  nand (_22239_, _22238_, _09858_);
  nand (_22240_, _09000_, _06098_);
  or (_22241_, _22233_, _09000_);
  and (_22242_, _22241_, _02972_);
  nand (_22243_, _22242_, _22240_);
  and (_22244_, _22243_, _03397_);
  nand (_22245_, _22244_, _22239_);
  nand (_22246_, _09008_, _06098_);
  or (_22248_, _22233_, _09008_);
  and (_22249_, _22248_, _22246_);
  or (_22250_, _22249_, _03397_);
  nand (_22251_, _22250_, _22245_);
  nand (_22252_, _22251_, _08969_);
  and (_22253_, _22252_, _22149_);
  or (_22254_, _22253_, _22139_);
  nand (_22255_, _22254_, _06189_);
  and (_22256_, _05476_, _02790_);
  nor (_22257_, _22256_, _04230_);
  nand (_22259_, _22257_, _22255_);
  nor (_22260_, _05256_, _02533_);
  nor (_22261_, _22260_, _20432_);
  and (_22262_, _22261_, _22259_);
  or (_22263_, _22262_, _22137_);
  nand (_22264_, _22263_, _09273_);
  nor (_22265_, _22129_, _09273_);
  nor (_22266_, _22265_, _02902_);
  nand (_22267_, _22266_, _22264_);
  and (_22268_, _05318_, _02902_);
  nor (_22270_, _22268_, _09277_);
  nand (_22271_, _22270_, _22267_);
  and (_22272_, _05256_, _09277_);
  nor (_22273_, _22272_, _02901_);
  nand (_22274_, _22273_, _22271_);
  and (_22275_, _05318_, _02901_);
  nor (_22276_, _22275_, _20447_);
  and (_22277_, _22276_, _22274_);
  or (_22278_, _22277_, _22136_);
  nand (_22279_, _22278_, _09289_);
  nor (_22281_, _09289_, _05318_);
  nor (_22282_, _22281_, _07700_);
  and (_22283_, _22282_, _22279_);
  nor (_22284_, _22138_, _02499_);
  or (_22285_, _22284_, _02785_);
  nor (_22286_, _22285_, _22283_);
  and (_22287_, _05476_, _02785_);
  or (_22288_, _22287_, _22286_);
  nand (_22289_, _22288_, _04132_);
  and (_22290_, _05256_, _02518_);
  nor (_22292_, _22290_, _02975_);
  nand (_22293_, _22292_, _22289_);
  and (_22294_, _06098_, _02975_);
  not (_22295_, _22294_);
  and (_22296_, _22295_, _09305_);
  nand (_22297_, _22296_, _22293_);
  nor (_22298_, _09305_, _05318_);
  nor (_22299_, _22298_, _02524_);
  and (_22300_, _22299_, _22297_);
  nor (_22301_, _08824_, _06098_);
  nor (_22303_, _22301_, _10325_);
  or (_22304_, _22303_, _22300_);
  and (_22305_, _22138_, _08824_);
  nor (_22306_, _22305_, _02894_);
  nand (_22307_, _22306_, _22304_);
  and (_22308_, _05318_, _02894_);
  nor (_22309_, _22308_, _02578_);
  nand (_22310_, _22309_, _22307_);
  and (_22311_, _05256_, _02578_);
  nor (_22312_, _22311_, _09318_);
  nand (_22314_, _22312_, _22310_);
  and (_22315_, _22155_, _09318_);
  nor (_22316_, _22315_, _05516_);
  and (_22317_, _22316_, _22314_);
  or (_22318_, _22317_, _22135_);
  nand (_22319_, _22318_, _05261_);
  and (_22320_, _08878_, _02974_);
  nor (_22321_, _22320_, _07807_);
  nand (_22322_, _22321_, _22319_);
  and (_22323_, _07807_, _05318_);
  nor (_22325_, _22323_, _09334_);
  nand (_22326_, _22325_, _22322_);
  and (_22327_, _09357_, _09341_);
  nor (_22328_, _22327_, _09358_);
  nor (_22329_, _22328_, _09335_);
  nor (_22330_, _22329_, _02893_);
  and (_22331_, _22330_, _22326_);
  and (_22332_, _05318_, _02893_);
  or (_22333_, _22332_, _02585_);
  or (_22334_, _22333_, _22331_);
  and (_22336_, _05256_, _02585_);
  nor (_22337_, _22336_, _09375_);
  nand (_22338_, _22337_, _22334_);
  and (_22339_, _08149_, _05318_);
  and (_22340_, _22155_, _09381_);
  or (_22341_, _22340_, _22339_);
  and (_22342_, _22341_, _09375_);
  nor (_22343_, _22342_, _09385_);
  and (_22344_, _22343_, _22338_);
  or (_22345_, _22344_, _22134_);
  nand (_22347_, _22345_, _08814_);
  nor (_22348_, _08814_, _05318_);
  nor (_22349_, _22348_, _02977_);
  and (_22350_, _22349_, _22347_);
  and (_22351_, _06098_, _02977_);
  or (_22352_, _22351_, _03107_);
  nor (_22353_, _22352_, _22350_);
  and (_22354_, _05476_, _03107_);
  or (_22355_, _22354_, _22353_);
  nand (_22356_, _22355_, _19652_);
  and (_22358_, _05256_, _02582_);
  nor (_22359_, _22358_, _09397_);
  nand (_22360_, _22359_, _22356_);
  or (_22361_, _22155_, _09381_);
  or (_22362_, _08149_, _05318_);
  and (_22363_, _22362_, _09397_);
  and (_22364_, _22363_, _22361_);
  nor (_22365_, _22364_, _09406_);
  and (_22366_, _22365_, _22360_);
  or (_22367_, _22366_, _22133_);
  nand (_22369_, _22367_, _07881_);
  nor (_22370_, _07881_, _05318_);
  nor (_22371_, _22370_, _02991_);
  and (_22372_, _22371_, _22369_);
  and (_22373_, _06098_, _02991_);
  or (_22374_, _22373_, _03094_);
  nor (_22375_, _22374_, _22372_);
  and (_22376_, _05476_, _03094_);
  or (_22377_, _22376_, _22375_);
  nand (_22378_, _22377_, _10353_);
  and (_22380_, _05256_, _02594_);
  nor (_22381_, _22380_, _08807_);
  nand (_22382_, _22381_, _22378_);
  nor (_22383_, _22155_, \oc8051_golden_model_1.PSW [7]);
  nor (_22384_, _05318_, _07294_);
  nor (_22385_, _22384_, _08808_);
  not (_22386_, _22385_);
  nor (_22387_, _22386_, _22383_);
  nor (_22388_, _22387_, _09418_);
  and (_22389_, _22388_, _22382_);
  or (_22391_, _22389_, _22132_);
  nand (_22392_, _22391_, _07900_);
  nor (_22393_, _07900_, _05318_);
  nor (_22394_, _22393_, _02994_);
  and (_22395_, _22394_, _22392_);
  and (_22396_, _06098_, _02994_);
  or (_22397_, _22396_, _03099_);
  nor (_22398_, _22397_, _22395_);
  and (_22399_, _05476_, _03099_);
  or (_22400_, _22399_, _22398_);
  nand (_22402_, _22400_, _02590_);
  and (_22403_, _05256_, _02589_);
  nor (_22404_, _22403_, _08799_);
  nand (_22405_, _22404_, _22402_);
  nor (_22406_, _22155_, _07294_);
  nor (_22407_, _05318_, \oc8051_golden_model_1.PSW [7]);
  nor (_22408_, _22407_, _08800_);
  not (_22409_, _22408_);
  nor (_22410_, _22409_, _22406_);
  nor (_22411_, _22410_, _09434_);
  and (_22413_, _22411_, _22405_);
  or (_22414_, _22413_, _22131_);
  nand (_22415_, _22414_, _07947_);
  nor (_22416_, _07947_, _05318_);
  nor (_22417_, _22416_, _08027_);
  and (_22418_, _22417_, _22415_);
  and (_22419_, _22129_, _08027_);
  or (_22420_, _22419_, _03113_);
  nor (_22421_, _22420_, _22418_);
  nor (_22422_, _05426_, _10159_);
  or (_22424_, _22422_, _22421_);
  nand (_22425_, _22424_, _05741_);
  and (_22426_, _05256_, _02592_);
  nor (_22427_, _22426_, _02993_);
  nand (_22428_, _22427_, _22425_);
  and (_22429_, _22233_, _09640_);
  nor (_22430_, _09640_, _06098_);
  or (_22431_, _22430_, _03549_);
  or (_22432_, _22431_, _22429_);
  and (_22433_, _22432_, _08795_);
  and (_22435_, _22433_, _22428_);
  or (_22436_, _22435_, _22130_);
  nand (_22437_, _22436_, _20297_);
  and (_22438_, _08772_, _05476_);
  nor (_22439_, _22438_, _07143_);
  nand (_22440_, _22439_, _22437_);
  and (_22441_, _22129_, _07143_);
  nor (_22442_, _22441_, _02854_);
  and (_22443_, _22442_, _22440_);
  nor (_22444_, _05426_, _02855_);
  or (_22446_, _22444_, _22443_);
  nand (_22447_, _22446_, _19640_);
  and (_22448_, _05256_, _02575_);
  nor (_22449_, _22448_, _02990_);
  nand (_22450_, _22449_, _22447_);
  nor (_22451_, _22143_, _09640_);
  and (_22452_, _09640_, _08878_);
  nor (_22453_, _22452_, _22451_);
  and (_22454_, _22453_, _02990_);
  nor (_22455_, _22454_, _09668_);
  nand (_22457_, _22455_, _22450_);
  nor (_22458_, _22129_, _09667_);
  nor (_22459_, _22458_, _03133_);
  and (_22460_, _22459_, _22457_);
  or (_22461_, _22460_, _22127_);
  nand (_22462_, _22461_, _09675_);
  nor (_22463_, _22138_, _09675_);
  nor (_22464_, _22463_, _04331_);
  nand (_22465_, _22464_, _22462_);
  and (_22466_, _05256_, _04331_);
  nor (_22468_, _22466_, _02778_);
  nand (_22469_, _22468_, _22465_);
  and (_22470_, _22453_, _02778_);
  nor (_22471_, _22470_, _09689_);
  nand (_22472_, _22471_, _22469_);
  nor (_22473_, _22129_, _09688_);
  nor (_22474_, _22473_, _02852_);
  and (_22475_, _22474_, _22472_);
  and (_22476_, _09696_, _05476_);
  nor (_22477_, _22476_, _10371_);
  nor (_22479_, _22477_, _22475_);
  nor (_22480_, _22129_, _09696_);
  or (_22481_, _22480_, _22479_);
  nand (_22482_, _22481_, _10310_);
  and (_22483_, _19634_, _05256_);
  nor (_22484_, _22483_, _09706_);
  and (_22485_, _22484_, _22482_);
  and (_22486_, _22129_, _09706_);
  or (_22487_, _22486_, _22485_);
  or (_22488_, _22487_, _34450_);
  or (_22490_, _34446_, \oc8051_golden_model_1.PC [7]);
  and (_22491_, _22490_, _35583_);
  and (_35629_[7], _22491_, _22488_);
  nor (_22492_, _09699_, _02835_);
  nor (_22493_, _05219_, _02835_);
  nor (_22494_, _08776_, \oc8051_golden_model_1.PC [8]);
  nor (_22495_, _22494_, _08783_);
  nor (_22496_, _22495_, _08795_);
  nor (_22497_, _22495_, _08797_);
  nor (_22498_, _22495_, _08805_);
  nor (_22500_, _22495_, _08812_);
  and (_22501_, _08935_, _02977_);
  nor (_22502_, _22495_, _08822_);
  nor (_22503_, _09067_, _05267_);
  nor (_22504_, _09318_, _02578_);
  nor (_22505_, _20048_, _09067_);
  and (_22506_, _08940_, _08933_);
  nor (_22507_, _22506_, _08941_);
  not (_22508_, _22507_);
  nor (_22509_, _22508_, _09000_);
  and (_22511_, _09000_, _08935_);
  or (_22512_, _22511_, _22509_);
  and (_22513_, _22512_, _02972_);
  and (_22514_, _09008_, _08935_);
  nor (_22515_, _22508_, _09008_);
  nor (_22516_, _22515_, _22514_);
  nor (_22517_, _22516_, _03397_);
  nor (_22518_, _02795_, _09209_);
  and (_22519_, _09067_, _02796_);
  nor (_22520_, _02930_, _04239_);
  and (_22522_, _09067_, _02799_);
  and (_22523_, _22508_, _09023_);
  and (_22524_, _09025_, _08936_);
  nor (_22525_, _22524_, _22523_);
  nor (_22526_, _22525_, _06162_);
  and (_22527_, _09120_, _09117_);
  nor (_22528_, _22527_, _09121_);
  and (_22529_, _22528_, _09148_);
  and (_22530_, _09150_, _09067_);
  or (_22531_, _22530_, _22529_);
  nor (_22533_, _22531_, _05325_);
  and (_22534_, _22495_, _07428_);
  and (_22535_, _09067_, _02934_);
  and (_22536_, _09067_, _02837_);
  and (_22537_, _09168_, \oc8051_golden_model_1.PC [8]);
  nor (_22538_, _22537_, _22536_);
  nor (_22539_, _22538_, _20341_);
  not (_22540_, _22539_);
  not (_22541_, _21085_);
  not (_22542_, _22495_);
  nor (_22544_, _22542_, _09164_);
  nor (_22545_, _22544_, _22541_);
  and (_22546_, _22545_, _22540_);
  nor (_22547_, _22495_, _09159_);
  nor (_22548_, _22547_, _02934_);
  not (_22549_, _22548_);
  nor (_22550_, _22549_, _22546_);
  nor (_22551_, _22550_, _22535_);
  nor (_22552_, _22551_, _07428_);
  or (_22553_, _22552_, _09178_);
  nor (_22555_, _22553_, _22534_);
  nor (_22556_, _22555_, _07425_);
  and (_22557_, _22495_, _07425_);
  nor (_22558_, _22557_, _05327_);
  not (_22559_, _22558_);
  nor (_22560_, _22559_, _22556_);
  or (_22561_, _22560_, _03806_);
  or (_22562_, _22561_, _22533_);
  nand (_22563_, _22495_, _03806_);
  and (_22564_, _22563_, _06162_);
  and (_22566_, _22564_, _22562_);
  or (_22567_, _22566_, _22526_);
  nand (_22568_, _22567_, _09018_);
  nor (_22569_, _22495_, _09018_);
  nor (_22570_, _22569_, _02799_);
  and (_22571_, _22570_, _22568_);
  or (_22572_, _22571_, _22522_);
  nand (_22573_, _22572_, _22520_);
  and (_22574_, _09067_, _02930_);
  nor (_22575_, _22574_, _09200_);
  nand (_22577_, _22575_, _22573_);
  nor (_22578_, _22495_, _09199_);
  nor (_22579_, _22578_, _02928_);
  nand (_22580_, _22579_, _22577_);
  and (_22581_, _09067_, _02928_);
  nor (_22582_, _22581_, _09206_);
  nand (_22583_, _22582_, _22580_);
  and (_22584_, _22542_, _09206_);
  nor (_22585_, _22584_, _02796_);
  and (_22586_, _22585_, _22583_);
  or (_22588_, _22586_, _22519_);
  nand (_22589_, _22588_, _22518_);
  and (_22590_, _09067_, _02795_);
  nor (_22591_, _22590_, _09906_);
  nand (_22592_, _22591_, _22589_);
  not (_22593_, _02973_);
  and (_22594_, _09252_, _08935_);
  nor (_22595_, _22508_, _09252_);
  or (_22596_, _22595_, _22594_);
  nor (_22597_, _22596_, _09217_);
  nor (_22599_, _22597_, _22593_);
  and (_22600_, _22599_, _22592_);
  or (_22601_, _22600_, _22517_);
  or (_22602_, _22601_, _22513_);
  nand (_22603_, _22602_, _08969_);
  and (_22604_, _08936_, _08839_);
  nor (_22605_, _22507_, _08839_);
  or (_22606_, _22605_, _08969_);
  nor (_22607_, _22606_, _22604_);
  nor (_22608_, _22607_, _08827_);
  nand (_22610_, _22608_, _22603_);
  and (_22611_, _22542_, _08827_);
  nor (_22612_, _22611_, _02790_);
  nand (_22613_, _22612_, _22610_);
  and (_22614_, _09067_, _02790_);
  not (_22615_, _22614_);
  and (_22616_, _20048_, _02533_);
  and (_22617_, _22616_, _22615_);
  and (_22618_, _22617_, _22613_);
  or (_22619_, _22618_, _22505_);
  nand (_22621_, _22619_, _09273_);
  nor (_22622_, _22495_, _09273_);
  nor (_22623_, _22622_, _02902_);
  nand (_22624_, _22623_, _22621_);
  and (_22625_, _09067_, _02902_);
  nor (_22626_, _22625_, _09277_);
  nand (_22627_, _22626_, _22624_);
  nand (_22628_, _22627_, _09759_);
  and (_22629_, _09067_, _02901_);
  nor (_22630_, _22629_, _20447_);
  and (_22632_, _22630_, _22628_);
  nor (_22633_, _22495_, _09285_);
  or (_22634_, _22633_, _22632_);
  nand (_22635_, _22634_, _09289_);
  nor (_22636_, _09289_, _09067_);
  nor (_22637_, _22636_, _07700_);
  nand (_22638_, _22637_, _22635_);
  nor (_22639_, _22542_, _02499_);
  nor (_22640_, _22639_, _02785_);
  nand (_22641_, _22640_, _22638_);
  and (_22643_, _09068_, _02785_);
  nor (_22644_, _02975_, _02518_);
  not (_22645_, _22644_);
  nor (_22646_, _22645_, _22643_);
  nand (_22647_, _22646_, _22641_);
  and (_22648_, _08935_, _02975_);
  not (_22649_, _22648_);
  and (_22650_, _22649_, _09305_);
  nand (_22651_, _22650_, _22647_);
  nor (_22652_, _09305_, _09067_);
  nor (_22654_, _22652_, _02524_);
  and (_22655_, _22654_, _22651_);
  nor (_22656_, _08935_, _08824_);
  nor (_22657_, _22656_, _10325_);
  or (_22658_, _22657_, _22655_);
  and (_22659_, _22542_, _08824_);
  nor (_22660_, _22659_, _02894_);
  and (_22661_, _22660_, _22658_);
  and (_22662_, _09067_, _02894_);
  or (_22663_, _22662_, _22661_);
  nand (_22665_, _22663_, _22504_);
  and (_22666_, _22528_, _09318_);
  nor (_22667_, _22666_, _05516_);
  and (_22668_, _22667_, _22665_);
  or (_22669_, _22668_, _22503_);
  nand (_22670_, _22669_, _05261_);
  and (_22671_, _08936_, _02974_);
  nor (_22672_, _22671_, _07807_);
  nand (_22673_, _22672_, _22670_);
  and (_22674_, _09067_, _07807_);
  nor (_22676_, _22674_, _09334_);
  nand (_22677_, _22676_, _22673_);
  and (_22678_, _09359_, _09337_);
  nor (_22679_, _22678_, _09360_);
  nor (_22680_, _22679_, _09335_);
  nor (_22681_, _22680_, _02893_);
  nand (_22682_, _22681_, _22677_);
  and (_22683_, _09067_, _02893_);
  nor (_22684_, _22683_, _02585_);
  nand (_22685_, _22684_, _22682_);
  nand (_22687_, _22685_, _09376_);
  nor (_22688_, _22528_, _08149_);
  nor (_22689_, _09067_, _09381_);
  nor (_22690_, _22689_, _09376_);
  not (_22691_, _22690_);
  nor (_22692_, _22691_, _22688_);
  nor (_22693_, _22692_, _09385_);
  and (_22694_, _22693_, _22687_);
  or (_22695_, _22694_, _22502_);
  nand (_22696_, _22695_, _08814_);
  nor (_22698_, _08814_, _09067_);
  nor (_22699_, _22698_, _02977_);
  and (_22700_, _22699_, _22696_);
  or (_22701_, _22700_, _22501_);
  nand (_22702_, _22701_, _07104_);
  and (_22703_, _09067_, _03107_);
  nor (_22704_, _22703_, _02582_);
  nand (_22705_, _22704_, _22702_);
  nand (_22706_, _22705_, _09398_);
  or (_22707_, _22528_, _09381_);
  or (_22709_, _09067_, _08149_);
  and (_22710_, _22709_, _09397_);
  and (_22711_, _22710_, _22707_);
  nor (_22712_, _22711_, _09406_);
  and (_22713_, _22712_, _22706_);
  or (_22714_, _22713_, _22500_);
  nand (_22715_, _22714_, _07881_);
  nor (_22716_, _09067_, _07881_);
  nor (_22717_, _22716_, _02991_);
  and (_22718_, _22717_, _22715_);
  and (_22720_, _08935_, _02991_);
  or (_22721_, _22720_, _03094_);
  or (_22722_, _22721_, _22718_);
  nor (_22723_, _08807_, _02594_);
  and (_22724_, _09068_, _03094_);
  not (_22725_, _22724_);
  and (_22726_, _22725_, _22723_);
  nand (_22727_, _22726_, _22722_);
  nor (_22728_, _22528_, \oc8051_golden_model_1.PSW [7]);
  nor (_22729_, _09067_, _07294_);
  nor (_22731_, _22729_, _08808_);
  not (_22732_, _22731_);
  nor (_22733_, _22732_, _22728_);
  nor (_22734_, _22733_, _09418_);
  and (_22735_, _22734_, _22727_);
  or (_22736_, _22735_, _22498_);
  nand (_22737_, _22736_, _07900_);
  nor (_22738_, _09067_, _07900_);
  nor (_22739_, _22738_, _02994_);
  and (_22740_, _22739_, _22737_);
  and (_22742_, _08935_, _02994_);
  or (_22743_, _22742_, _03099_);
  or (_22744_, _22743_, _22740_);
  nor (_22745_, _08799_, _02589_);
  and (_22746_, _09068_, _03099_);
  not (_22747_, _22746_);
  and (_22748_, _22747_, _22745_);
  nand (_22749_, _22748_, _22744_);
  nor (_22750_, _22528_, _07294_);
  nor (_22751_, _09067_, \oc8051_golden_model_1.PSW [7]);
  nor (_22753_, _22751_, _08800_);
  not (_22754_, _22753_);
  nor (_22755_, _22754_, _22750_);
  nor (_22756_, _22755_, _09434_);
  and (_22757_, _22756_, _22749_);
  or (_22758_, _22757_, _22497_);
  nand (_22759_, _22758_, _07947_);
  nor (_22760_, _09067_, _07947_);
  nor (_22761_, _22760_, _08027_);
  and (_22762_, _22761_, _22759_);
  and (_22764_, _22495_, _08027_);
  or (_22765_, _22764_, _22762_);
  nand (_22766_, _22765_, _10159_);
  and (_22767_, _03805_, _03113_);
  nor (_22768_, _22767_, _02592_);
  nand (_22769_, _22768_, _22766_);
  nand (_22770_, _22769_, _03549_);
  nor (_22771_, _09640_, _08935_);
  and (_22772_, _22508_, _09640_);
  or (_22773_, _22772_, _03549_);
  or (_22774_, _22773_, _22771_);
  and (_22775_, _22774_, _08795_);
  and (_22776_, _22775_, _22770_);
  or (_22777_, _22776_, _22496_);
  nand (_22778_, _22777_, _20297_);
  and (_22779_, _09068_, _08772_);
  nor (_22780_, _22779_, _07143_);
  and (_22781_, _22780_, _22778_);
  and (_22782_, _22495_, _07143_);
  or (_22783_, _22782_, _22781_);
  nand (_22785_, _22783_, _02855_);
  and (_22786_, _03805_, _02854_);
  nor (_22787_, _22786_, _02575_);
  nand (_22788_, _22787_, _22785_);
  nand (_22789_, _22788_, _03134_);
  nor (_22790_, _22507_, _09640_);
  and (_22791_, _09640_, _08936_);
  nor (_22792_, _22791_, _22790_);
  and (_22793_, _22792_, _02990_);
  nor (_22794_, _22793_, _09668_);
  nand (_22796_, _22794_, _22789_);
  nor (_22797_, _22495_, _09667_);
  nor (_22798_, _22797_, _03133_);
  nand (_22799_, _22798_, _22796_);
  and (_22800_, _09067_, _03133_);
  nor (_22801_, _22800_, _21371_);
  nand (_22802_, _22801_, _22799_);
  nor (_22803_, _22495_, _09675_);
  nor (_22804_, _22803_, _02988_);
  and (_22805_, _22804_, _22802_);
  or (_22806_, _22805_, _22493_);
  nor (_22807_, _02778_, _02572_);
  nand (_22808_, _22807_, _22806_);
  and (_22809_, _22792_, _02778_);
  nor (_22810_, _22809_, _09689_);
  nand (_22811_, _22810_, _22808_);
  nor (_22812_, _22495_, _09688_);
  nor (_22813_, _22812_, _02852_);
  nand (_22814_, _22813_, _22811_);
  and (_22815_, _09067_, _02852_);
  nor (_22816_, _22815_, _21033_);
  nand (_22817_, _22816_, _22814_);
  nor (_22818_, _22495_, _09696_);
  nor (_22819_, _22818_, _02982_);
  and (_22820_, _22819_, _22817_);
  or (_22821_, _22820_, _22492_);
  nor (_22822_, _09706_, _02568_);
  and (_22823_, _22822_, _22821_);
  and (_22824_, _22495_, _09706_);
  or (_22825_, _22824_, _22823_);
  or (_22826_, _22825_, _34450_);
  or (_22827_, _34446_, \oc8051_golden_model_1.PC [8]);
  and (_22828_, _22827_, _35583_);
  and (_35629_[8], _22828_, _22826_);
  nor (_22829_, _03742_, _05219_);
  nor (_22830_, _08783_, \oc8051_golden_model_1.PC [9]);
  nor (_22831_, _22830_, _08784_);
  nor (_22832_, _22831_, _08795_);
  nor (_22833_, _22831_, _08797_);
  and (_22834_, _08873_, _02994_);
  nor (_22835_, _22831_, _08805_);
  and (_22836_, _08873_, _02991_);
  nor (_22837_, _22831_, _08812_);
  and (_22838_, _08873_, _02977_);
  nor (_22839_, _22831_, _08822_);
  nor (_22840_, _09061_, _05267_);
  not (_22841_, _22831_);
  and (_22842_, _22841_, _08827_);
  and (_22843_, _09061_, _02795_);
  nand (_22844_, _09061_, _02934_);
  nand (_22845_, _09061_, _02837_);
  nand (_22846_, _09168_, \oc8051_golden_model_1.PC [9]);
  and (_22847_, _22846_, _22845_);
  or (_22848_, _22847_, _20341_);
  or (_22849_, _22841_, _09164_);
  and (_22850_, _22849_, _21085_);
  and (_22851_, _22850_, _22848_);
  nor (_22852_, _22831_, _09159_);
  or (_22853_, _22852_, _02934_);
  or (_22854_, _22853_, _22851_);
  and (_22856_, _22854_, _22844_);
  or (_22857_, _22856_, _07428_);
  nand (_22858_, _22831_, _07428_);
  and (_22859_, _22858_, _02544_);
  and (_22860_, _22859_, _22857_);
  or (_22861_, _22860_, _07425_);
  nand (_22862_, _22831_, _07425_);
  and (_22863_, _22862_, _05325_);
  and (_22864_, _22863_, _22861_);
  or (_22865_, _09063_, _09064_);
  and (_22867_, _22865_, _09122_);
  nor (_22868_, _22865_, _09122_);
  or (_22869_, _22868_, _22867_);
  or (_22870_, _22869_, _09150_);
  or (_22871_, _09148_, _09062_);
  and (_22872_, _22871_, _22870_);
  and (_22873_, _22872_, _05327_);
  or (_22874_, _22873_, _22864_);
  and (_22875_, _22874_, _05311_);
  and (_22876_, _22841_, _03806_);
  or (_22877_, _22876_, _02932_);
  or (_22878_, _22877_, _22875_);
  and (_22879_, _19708_, _08874_);
  nor (_22880_, _08941_, _08937_);
  and (_22881_, _22880_, _08877_);
  nor (_22882_, _22880_, _08877_);
  nor (_22883_, _22882_, _22881_);
  and (_22884_, _22883_, _09023_);
  or (_22885_, _22884_, _06162_);
  or (_22886_, _22885_, _22879_);
  and (_22888_, _22886_, _09018_);
  and (_22889_, _22888_, _22878_);
  nor (_22890_, _22831_, _09018_);
  or (_22891_, _22890_, _02799_);
  or (_22892_, _22891_, _22889_);
  nand (_22893_, _09061_, _02799_);
  and (_22894_, _22893_, _02540_);
  and (_22895_, _22894_, _22892_);
  nor (_22896_, _22895_, _02930_);
  and (_22897_, _09061_, _02930_);
  nor (_22899_, _22897_, _09200_);
  not (_22900_, _22899_);
  nor (_22901_, _22900_, _22896_);
  nor (_22902_, _22831_, _09199_);
  nor (_22903_, _22902_, _02928_);
  not (_22904_, _22903_);
  nor (_22905_, _22904_, _22901_);
  and (_22906_, _09061_, _02928_);
  nor (_22907_, _22906_, _09206_);
  not (_22908_, _22907_);
  nor (_22909_, _22908_, _22905_);
  and (_22910_, _22841_, _09206_);
  nor (_22911_, _22910_, _02796_);
  not (_22912_, _22911_);
  nor (_22913_, _22912_, _22909_);
  and (_22914_, _09062_, _02538_);
  nor (_22915_, _22914_, _09210_);
  or (_22916_, _22915_, _22913_);
  and (_22917_, _22916_, _03932_);
  or (_22918_, _22917_, _09906_);
  nor (_22921_, _22918_, _22843_);
  and (_22922_, _09252_, _08873_);
  nor (_22923_, _22883_, _09252_);
  or (_22924_, _22923_, _22922_);
  nor (_22925_, _22924_, _09217_);
  or (_22926_, _22925_, _22921_);
  nand (_22927_, _22926_, _09858_);
  and (_22928_, _09000_, _08873_);
  nor (_22929_, _22883_, _09000_);
  or (_22930_, _22929_, _22928_);
  nor (_22931_, _22930_, _09858_);
  nor (_22932_, _22931_, _02944_);
  nand (_22933_, _22932_, _22927_);
  and (_22934_, _09008_, _08874_);
  not (_22935_, _22883_);
  nor (_22936_, _22935_, _09008_);
  or (_22937_, _22936_, _03397_);
  or (_22938_, _22937_, _22934_);
  nand (_22939_, _22938_, _22933_);
  nand (_22940_, _22939_, _08969_);
  and (_22941_, _08874_, _08839_);
  and (_22942_, _22883_, _22141_);
  or (_22943_, _22942_, _08969_);
  nor (_22944_, _22943_, _22941_);
  nor (_22945_, _22944_, _08827_);
  and (_22946_, _22945_, _22940_);
  or (_22947_, _22946_, _22842_);
  nand (_22948_, _22947_, _06189_);
  and (_22949_, _09062_, _02790_);
  not (_22950_, _22949_);
  and (_22953_, _22950_, _22616_);
  nand (_22954_, _22953_, _22948_);
  nor (_22955_, _20048_, _09062_);
  nor (_22956_, _22955_, _09281_);
  nand (_22957_, _22956_, _22954_);
  nor (_22958_, _22831_, _09273_);
  nor (_22959_, _22958_, _02902_);
  and (_22960_, _22959_, _22957_);
  and (_22961_, _09061_, _02902_);
  or (_22962_, _22961_, _22960_);
  nand (_22964_, _22962_, _09278_);
  and (_22965_, _09061_, _02901_);
  nor (_22966_, _22965_, _20447_);
  and (_22967_, _22966_, _22964_);
  nor (_22968_, _22831_, _09285_);
  or (_22969_, _22968_, _22967_);
  nand (_22970_, _22969_, _09289_);
  nor (_22971_, _09289_, _09061_);
  nor (_22972_, _22971_, _07700_);
  nand (_22973_, _22972_, _22970_);
  nor (_22974_, _22841_, _02499_);
  nor (_22975_, _22974_, _02785_);
  nand (_22976_, _22975_, _22973_);
  and (_22977_, _09062_, _02785_);
  nor (_22978_, _22977_, _22645_);
  nand (_22979_, _22978_, _22976_);
  and (_22980_, _08873_, _02975_);
  not (_22981_, _22980_);
  and (_22982_, _22981_, _09305_);
  nand (_22983_, _22982_, _22979_);
  nor (_22986_, _09305_, _09061_);
  nor (_22987_, _22986_, _02524_);
  and (_22988_, _22987_, _22983_);
  nor (_22989_, _08873_, _08824_);
  nor (_22990_, _22989_, _10325_);
  or (_22991_, _22990_, _22988_);
  and (_22992_, _22841_, _08824_);
  nor (_22993_, _22992_, _02894_);
  and (_22994_, _22993_, _22991_);
  and (_22995_, _09061_, _02894_);
  or (_22996_, _22995_, _22994_);
  nand (_22997_, _22996_, _22504_);
  nor (_22998_, _22869_, _09319_);
  nor (_22999_, _22998_, _05516_);
  and (_23000_, _22999_, _22997_);
  or (_23001_, _23000_, _22840_);
  nand (_23002_, _23001_, _05261_);
  and (_23003_, _08874_, _02974_);
  nor (_23004_, _23003_, _07807_);
  nand (_23005_, _23004_, _23002_);
  and (_23006_, _09061_, _07807_);
  nor (_23007_, _23006_, _09334_);
  nand (_23008_, _23007_, _23005_);
  nor (_23009_, _09360_, \oc8051_golden_model_1.DPH [1]);
  nor (_23010_, _23009_, _09361_);
  nor (_23011_, _23010_, _09335_);
  nor (_23012_, _23011_, _02893_);
  nand (_23013_, _23012_, _23008_);
  and (_23014_, _09061_, _02893_);
  nor (_23015_, _23014_, _02585_);
  nand (_23018_, _23015_, _23013_);
  nand (_23019_, _23018_, _09376_);
  and (_23020_, _09061_, _08149_);
  nor (_23021_, _22869_, _08149_);
  or (_23022_, _23021_, _23020_);
  and (_23023_, _23022_, _09375_);
  nor (_23024_, _23023_, _09385_);
  and (_23025_, _23024_, _23019_);
  or (_23026_, _23025_, _22839_);
  nand (_23027_, _23026_, _08814_);
  nor (_23029_, _08814_, _09061_);
  nor (_23030_, _23029_, _02977_);
  and (_23031_, _23030_, _23027_);
  or (_23032_, _23031_, _22838_);
  nand (_23033_, _23032_, _07104_);
  and (_23034_, _09061_, _03107_);
  nor (_23035_, _23034_, _02582_);
  nand (_23036_, _23035_, _23033_);
  nand (_23037_, _23036_, _09398_);
  nand (_23038_, _22869_, _08149_);
  or (_23040_, _09061_, _08149_);
  and (_23041_, _23040_, _09397_);
  and (_23042_, _23041_, _23038_);
  nor (_23043_, _23042_, _09406_);
  and (_23044_, _23043_, _23037_);
  or (_23045_, _23044_, _22837_);
  nand (_23046_, _23045_, _07881_);
  nor (_23047_, _09061_, _07881_);
  nor (_23048_, _23047_, _02991_);
  and (_23049_, _23048_, _23046_);
  or (_23051_, _23049_, _22836_);
  nand (_23052_, _23051_, _06161_);
  and (_23053_, _09061_, _03094_);
  nor (_23054_, _23053_, _02594_);
  nand (_23055_, _23054_, _23052_);
  nand (_23056_, _23055_, _08808_);
  and (_23057_, _22869_, _07294_);
  nor (_23058_, _09061_, _07294_);
  nor (_23059_, _23058_, _08808_);
  not (_23060_, _23059_);
  nor (_23061_, _23060_, _23057_);
  nor (_23062_, _23061_, _09418_);
  and (_23063_, _23062_, _23056_);
  or (_23064_, _23063_, _22835_);
  nand (_23065_, _23064_, _07900_);
  nor (_23066_, _09061_, _07900_);
  nor (_23067_, _23066_, _02994_);
  and (_23068_, _23067_, _23065_);
  or (_23069_, _23068_, _22834_);
  nand (_23070_, _23069_, _07118_);
  and (_23072_, _09061_, _03099_);
  nor (_23073_, _23072_, _02589_);
  nand (_23074_, _23073_, _23070_);
  nand (_23075_, _23074_, _08800_);
  and (_23076_, _22869_, \oc8051_golden_model_1.PSW [7]);
  nor (_23077_, _09061_, \oc8051_golden_model_1.PSW [7]);
  nor (_23078_, _23077_, _08800_);
  not (_23079_, _23078_);
  nor (_23080_, _23079_, _23076_);
  nor (_23081_, _23080_, _09434_);
  and (_23083_, _23081_, _23075_);
  or (_23084_, _23083_, _22833_);
  nand (_23085_, _23084_, _07947_);
  nor (_23086_, _09061_, _07947_);
  nor (_23087_, _23086_, _08027_);
  nand (_23088_, _23087_, _23085_);
  and (_23089_, _22831_, _08027_);
  nor (_23090_, _23089_, _03113_);
  nand (_23091_, _23090_, _23088_);
  nor (_23092_, _02993_, _02592_);
  not (_23094_, _23092_);
  and (_23095_, _03989_, _03113_);
  nor (_23096_, _23095_, _23094_);
  nand (_23097_, _23096_, _23091_);
  and (_23098_, _22883_, _09640_);
  nor (_23099_, _09640_, _08873_);
  or (_23100_, _23099_, _03549_);
  or (_23101_, _23100_, _23098_);
  and (_23102_, _23101_, _08795_);
  and (_23103_, _23102_, _23097_);
  or (_23105_, _23103_, _22832_);
  nand (_23106_, _23105_, _20297_);
  and (_23107_, _09062_, _08772_);
  nor (_23108_, _23107_, _07143_);
  nand (_23109_, _23108_, _23106_);
  and (_23110_, _22831_, _07143_);
  nor (_23111_, _23110_, _02854_);
  nand (_23112_, _23111_, _23109_);
  nor (_23113_, _02990_, _02575_);
  not (_23114_, _23113_);
  and (_23116_, _03989_, _02854_);
  nor (_23117_, _23116_, _23114_);
  nand (_23118_, _23117_, _23112_);
  and (_23119_, _09640_, _08874_);
  nor (_23120_, _22935_, _09640_);
  nor (_23121_, _23120_, _23119_);
  and (_23122_, _23121_, _02990_);
  nor (_23123_, _23122_, _09668_);
  nand (_23124_, _23123_, _23118_);
  nor (_23125_, _22831_, _09667_);
  nor (_23126_, _23125_, _03133_);
  nand (_23127_, _23126_, _23124_);
  and (_23128_, _09061_, _03133_);
  nor (_23129_, _23128_, _21371_);
  nand (_23130_, _23129_, _23127_);
  nor (_23131_, _22831_, _09675_);
  nor (_23132_, _23131_, _02988_);
  and (_23133_, _23132_, _23130_);
  or (_23134_, _23133_, _22829_);
  nand (_23135_, _23134_, _22807_);
  and (_23137_, _23121_, _02778_);
  nor (_23138_, _23137_, _09689_);
  nand (_23139_, _23138_, _23135_);
  nor (_23140_, _22831_, _09688_);
  nor (_23141_, _23140_, _02852_);
  and (_23142_, _23141_, _23139_);
  and (_23143_, _09696_, _09062_);
  nor (_23144_, _23143_, _10371_);
  or (_23145_, _23144_, _23142_);
  nor (_23146_, _22831_, _09696_);
  nor (_23148_, _23146_, _02982_);
  and (_23149_, _23148_, _23145_);
  nor (_23150_, _03742_, _09699_);
  or (_23151_, _23150_, _23149_);
  and (_23152_, _23151_, _22822_);
  and (_23153_, _22831_, _09706_);
  or (_23154_, _23153_, _23152_);
  or (_23155_, _23154_, _34450_);
  or (_23156_, _34446_, \oc8051_golden_model_1.PC [9]);
  and (_23157_, _23156_, _35583_);
  and (_35629_[9], _23157_, _23155_);
  nor (_23159_, _08784_, \oc8051_golden_model_1.PC [10]);
  nor (_23160_, _23159_, _08777_);
  not (_23161_, _23160_);
  nand (_23162_, _23161_, _07143_);
  nand (_23163_, _23161_, _08027_);
  nand (_23164_, _08866_, _02994_);
  nand (_23165_, _08866_, _02991_);
  nand (_23166_, _08866_, _02977_);
  nor (_23167_, _09055_, _05267_);
  or (_23169_, _23167_, _02974_);
  and (_23170_, _08866_, _02524_);
  nor (_23171_, _23170_, _08824_);
  nand (_23172_, _09055_, _02901_);
  nand (_23173_, _09055_, _02930_);
  and (_23174_, _09054_, _02799_);
  nor (_23175_, _08945_, _08942_);
  not (_23176_, _23175_);
  and (_23177_, _23176_, _08869_);
  nor (_23178_, _23176_, _08869_);
  nor (_23180_, _23178_, _23177_);
  or (_23181_, _23180_, _09025_);
  or (_23182_, _09023_, _08865_);
  and (_23183_, _23182_, _23181_);
  or (_23184_, _23183_, _06162_);
  nor (_23185_, _09125_, _09058_);
  nor (_23186_, _23185_, _09126_);
  and (_23187_, _23186_, _09148_);
  and (_23188_, _09150_, _09054_);
  or (_23189_, _23188_, _23187_);
  or (_23190_, _23189_, _05325_);
  or (_23191_, _23160_, _09159_);
  or (_23192_, _23160_, _09163_);
  nor (_23193_, _23161_, _09164_);
  and (_23194_, _09054_, _02837_);
  and (_23195_, _09168_, \oc8051_golden_model_1.PC [10]);
  or (_23196_, _23195_, _23194_);
  or (_23197_, _23196_, _23193_);
  and (_23198_, _23197_, _23192_);
  or (_23199_, _23198_, _22541_);
  and (_23201_, _23199_, _23191_);
  or (_23202_, _23201_, _02934_);
  and (_23203_, _09055_, _02934_);
  nor (_23204_, _23203_, _07428_);
  and (_23205_, _23204_, _23202_);
  and (_23206_, _23160_, _07428_);
  or (_23207_, _23206_, _09178_);
  or (_23208_, _23207_, _23205_);
  and (_23209_, _23208_, _21080_);
  nand (_23210_, _23160_, _07425_);
  nand (_23212_, _23210_, _05325_);
  or (_23213_, _23212_, _23209_);
  and (_23214_, _23213_, _05311_);
  and (_23215_, _23214_, _23190_);
  and (_23216_, _23160_, _03806_);
  or (_23217_, _23216_, _02932_);
  or (_23218_, _23217_, _23215_);
  nand (_23219_, _23218_, _23184_);
  nand (_23220_, _23219_, _09018_);
  or (_23221_, _23160_, _09018_);
  and (_23223_, _23221_, _03186_);
  and (_23224_, _23223_, _23220_);
  nor (_23225_, _23224_, _23174_);
  nand (_23226_, _23225_, _22520_);
  and (_23227_, _23226_, _23173_);
  and (_23228_, _23227_, _09199_);
  nor (_23229_, _23161_, _09199_);
  or (_23230_, _23229_, _02928_);
  or (_23231_, _23230_, _23228_);
  nand (_23232_, _09055_, _02928_);
  and (_23234_, _23232_, _23231_);
  or (_23235_, _23234_, _09206_);
  nand (_23236_, _23161_, _09206_);
  and (_23237_, _23236_, _02927_);
  and (_23238_, _23237_, _23235_);
  and (_23239_, _09054_, _02796_);
  or (_23240_, _23239_, _09209_);
  or (_23241_, _23240_, _23238_);
  and (_23242_, _23241_, _03932_);
  nand (_23243_, _09054_, _02795_);
  nand (_23245_, _23243_, _09217_);
  or (_23246_, _23245_, _23242_);
  or (_23247_, _23180_, _09252_);
  nand (_23248_, _09252_, _08866_);
  and (_23249_, _23248_, _23247_);
  or (_23250_, _23249_, _09217_);
  and (_23251_, _23250_, _23246_);
  or (_23252_, _23251_, _02972_);
  and (_23253_, _09000_, _08865_);
  not (_23254_, _09000_);
  and (_23255_, _23180_, _23254_);
  or (_23256_, _23255_, _09858_);
  or (_23257_, _23256_, _23253_);
  and (_23258_, _23257_, _03397_);
  and (_23259_, _23258_, _23252_);
  and (_23260_, _23180_, _09009_);
  and (_23261_, _09008_, _08865_);
  or (_23262_, _23261_, _23260_);
  and (_23263_, _23262_, _02944_);
  or (_23264_, _23263_, _23259_);
  and (_23266_, _23264_, _08969_);
  or (_23267_, _23180_, _08839_);
  nand (_23268_, _08866_, _08839_);
  and (_23269_, _23268_, _02979_);
  and (_23270_, _23269_, _23267_);
  or (_23271_, _23270_, _08827_);
  or (_23272_, _23271_, _23266_);
  nand (_23273_, _23161_, _08827_);
  and (_23274_, _20048_, _06189_);
  and (_23275_, _23274_, _23273_);
  and (_23277_, _23275_, _23272_);
  nor (_23278_, _23274_, _09055_);
  nand (_23279_, _09273_, _02533_);
  or (_23280_, _23279_, _23278_);
  or (_23281_, _23280_, _23277_);
  or (_23282_, _23160_, _09273_);
  and (_23283_, _23282_, _09276_);
  and (_23284_, _23283_, _23281_);
  and (_23285_, _09054_, _02902_);
  nor (_23286_, _23285_, _23284_);
  nand (_23288_, _23286_, _09278_);
  and (_23289_, _23288_, _23172_);
  or (_23290_, _23289_, _20447_);
  or (_23291_, _23160_, _09285_);
  and (_23292_, _23291_, _09289_);
  and (_23293_, _23292_, _23290_);
  nor (_23294_, _09289_, _09055_);
  or (_23295_, _23294_, _07700_);
  or (_23296_, _23295_, _23293_);
  nor (_23297_, _23160_, _02499_);
  nor (_23299_, _23297_, _02785_);
  and (_23300_, _23299_, _23296_);
  nand (_23301_, _09054_, _02785_);
  nand (_23302_, _23301_, _22644_);
  or (_23303_, _23302_, _23300_);
  nand (_23304_, _08866_, _02975_);
  and (_23305_, _23304_, _09305_);
  and (_23306_, _23305_, _23303_);
  nor (_23307_, _09305_, _09055_);
  or (_23308_, _23307_, _02524_);
  or (_23310_, _23308_, _23306_);
  and (_23311_, _23310_, _23171_);
  and (_23312_, _23160_, _08824_);
  or (_23313_, _23312_, _23311_);
  and (_23314_, _23313_, _03474_);
  nand (_23315_, _09054_, _02894_);
  nand (_23316_, _23315_, _22504_);
  or (_23317_, _23316_, _23314_);
  or (_23318_, _23186_, _09319_);
  and (_23319_, _23318_, _05267_);
  and (_23320_, _23319_, _23317_);
  or (_23321_, _23320_, _23169_);
  nand (_23322_, _08866_, _02974_);
  and (_23323_, _23322_, _23321_);
  or (_23324_, _23323_, _07807_);
  and (_23325_, _09055_, _07807_);
  nor (_23326_, _23325_, _09334_);
  and (_23327_, _23326_, _23324_);
  nor (_23328_, _09361_, \oc8051_golden_model_1.DPH [2]);
  nor (_23329_, _23328_, _09362_);
  and (_23331_, _23329_, _09334_);
  or (_23332_, _23331_, _02893_);
  or (_23333_, _23332_, _23327_);
  nor (_23334_, _09375_, _02585_);
  nand (_23335_, _09055_, _02893_);
  and (_23336_, _23335_, _23334_);
  and (_23337_, _23336_, _23333_);
  or (_23338_, _23186_, _08149_);
  or (_23339_, _09054_, _09381_);
  and (_23340_, _23339_, _09375_);
  and (_23342_, _23340_, _23338_);
  or (_23343_, _23342_, _09385_);
  or (_23344_, _23343_, _23337_);
  or (_23345_, _23160_, _08822_);
  and (_23346_, _23345_, _08814_);
  and (_23347_, _23346_, _23344_);
  nor (_23348_, _08814_, _09055_);
  or (_23349_, _23348_, _02977_);
  or (_23350_, _23349_, _23347_);
  and (_23351_, _23350_, _23166_);
  or (_23353_, _23351_, _03107_);
  nand (_23354_, _09055_, _03107_);
  nor (_23355_, _09397_, _02582_);
  and (_23356_, _23355_, _23354_);
  and (_23357_, _23356_, _23353_);
  or (_23358_, _23186_, _09381_);
  or (_23359_, _09054_, _08149_);
  and (_23360_, _23359_, _09397_);
  and (_23361_, _23360_, _23358_);
  or (_23362_, _23361_, _09406_);
  or (_23364_, _23362_, _23357_);
  or (_23365_, _23160_, _08812_);
  and (_23366_, _23365_, _07881_);
  and (_23367_, _23366_, _23364_);
  nor (_23368_, _09055_, _07881_);
  or (_23369_, _23368_, _02991_);
  or (_23370_, _23369_, _23367_);
  and (_23371_, _23370_, _23165_);
  or (_23372_, _23371_, _03094_);
  nand (_23373_, _09055_, _03094_);
  and (_23375_, _23373_, _22723_);
  and (_23376_, _23375_, _23372_);
  or (_23377_, _23186_, \oc8051_golden_model_1.PSW [7]);
  or (_23378_, _09054_, _07294_);
  and (_23379_, _23378_, _08807_);
  and (_23380_, _23379_, _23377_);
  or (_23381_, _23380_, _09418_);
  or (_23382_, _23381_, _23376_);
  or (_23383_, _23160_, _08805_);
  and (_23384_, _23383_, _07900_);
  and (_23386_, _23384_, _23382_);
  nor (_23387_, _09055_, _07900_);
  or (_23388_, _23387_, _02994_);
  or (_23389_, _23388_, _23386_);
  and (_23390_, _23389_, _23164_);
  or (_23391_, _23390_, _03099_);
  nand (_23392_, _09055_, _03099_);
  and (_23393_, _23392_, _22745_);
  and (_23394_, _23393_, _23391_);
  or (_23395_, _23186_, _07294_);
  or (_23397_, _09054_, \oc8051_golden_model_1.PSW [7]);
  and (_23398_, _23397_, _08799_);
  and (_23399_, _23398_, _23395_);
  or (_23400_, _23399_, _09434_);
  or (_23401_, _23400_, _23394_);
  or (_23402_, _23160_, _08797_);
  and (_23403_, _23402_, _07947_);
  and (_23404_, _23403_, _23401_);
  nor (_23405_, _09055_, _07947_);
  or (_23406_, _23405_, _08027_);
  or (_23408_, _23406_, _23404_);
  and (_23409_, _23408_, _23163_);
  or (_23410_, _23409_, _03113_);
  nand (_23411_, _04413_, _03113_);
  and (_23412_, _23411_, _23092_);
  and (_23413_, _23412_, _23410_);
  or (_23414_, _23180_, _09641_);
  or (_23415_, _09640_, _08865_);
  and (_23416_, _23415_, _02993_);
  and (_23417_, _23416_, _23414_);
  or (_23419_, _23417_, _09455_);
  or (_23420_, _23419_, _23413_);
  nor (_23421_, _23161_, _08772_);
  or (_23422_, _23421_, _10297_);
  and (_23423_, _23422_, _23420_);
  and (_23424_, _09054_, _08772_);
  or (_23425_, _23424_, _07143_);
  or (_23426_, _23425_, _23423_);
  and (_23427_, _23426_, _23162_);
  or (_23428_, _23427_, _02854_);
  nand (_23430_, _04413_, _02854_);
  and (_23431_, _23430_, _23113_);
  and (_23432_, _23431_, _23428_);
  nand (_23433_, _09640_, _08866_);
  or (_23434_, _23180_, _09640_);
  and (_23435_, _23434_, _23433_);
  and (_23436_, _23435_, _02990_);
  or (_23437_, _23436_, _09668_);
  or (_23438_, _23437_, _23432_);
  or (_23439_, _23160_, _09667_);
  and (_23441_, _23439_, _23438_);
  or (_23442_, _23441_, _03133_);
  nand (_23443_, _09055_, _03133_);
  and (_23444_, _23443_, _09675_);
  and (_23445_, _23444_, _23442_);
  nor (_23446_, _23161_, _09675_);
  or (_23447_, _23446_, _02988_);
  or (_23448_, _23447_, _23445_);
  nand (_23449_, _03320_, _02988_);
  and (_23450_, _23449_, _22807_);
  and (_23452_, _23450_, _23448_);
  and (_23453_, _23435_, _02778_);
  or (_23454_, _23453_, _09689_);
  or (_23455_, _23454_, _23452_);
  or (_23456_, _23160_, _09688_);
  and (_23457_, _23456_, _23455_);
  or (_23458_, _23457_, _02852_);
  nand (_23459_, _09055_, _02852_);
  and (_23460_, _23459_, _09696_);
  and (_23461_, _23460_, _23458_);
  nor (_23463_, _23161_, _09696_);
  or (_23464_, _23463_, _02982_);
  or (_23465_, _23464_, _23461_);
  nand (_23466_, _03320_, _02982_);
  and (_23467_, _23466_, _22822_);
  and (_23468_, _23467_, _23465_);
  and (_23469_, _23160_, _09706_);
  or (_23470_, _23469_, _23468_);
  or (_23471_, _23470_, _34450_);
  or (_23472_, _34446_, \oc8051_golden_model_1.PC [10]);
  and (_23474_, _23472_, _35583_);
  and (_35629_[10], _23474_, _23471_);
  not (_23475_, \oc8051_golden_model_1.PC [11]);
  nor (_23476_, _08777_, _23475_);
  and (_23477_, _08777_, _23475_);
  or (_23478_, _23477_, _23476_);
  and (_23479_, _23478_, _09706_);
  or (_23480_, _23478_, _08795_);
  or (_23481_, _23478_, _08797_);
  or (_23482_, _09048_, _08801_);
  and (_23484_, _23482_, _08800_);
  or (_23485_, _23478_, _08805_);
  or (_23486_, _09048_, _08809_);
  and (_23487_, _23486_, _08808_);
  or (_23488_, _23478_, _08822_);
  or (_23489_, _09048_, _05267_);
  nor (_23490_, _23177_, _08867_);
  and (_23491_, _23490_, _08862_);
  nor (_23492_, _23490_, _08862_);
  or (_23493_, _23492_, _23491_);
  and (_23495_, _23493_, _23254_);
  and (_23496_, _09000_, _08858_);
  or (_23497_, _23496_, _23495_);
  and (_23498_, _23497_, _02972_);
  and (_23499_, _09008_, _08858_);
  and (_23500_, _23493_, _09009_);
  or (_23501_, _23500_, _23499_);
  and (_23502_, _23501_, _02944_);
  or (_23503_, _09015_, _09048_);
  or (_23504_, _09023_, _08858_);
  or (_23506_, _23493_, _09025_);
  and (_23507_, _23506_, _02932_);
  and (_23508_, _23507_, _23504_);
  and (_23509_, _09150_, _09048_);
  or (_23510_, _09050_, _09051_);
  nand (_23511_, _23510_, _09127_);
  or (_23512_, _23510_, _09127_);
  and (_23513_, _23512_, _23511_);
  and (_23514_, _23513_, _09148_);
  or (_23515_, _23514_, _23509_);
  or (_23517_, _23515_, _05325_);
  and (_23518_, _09048_, _09178_);
  or (_23519_, _23478_, _09159_);
  and (_23520_, _23519_, _07406_);
  and (_23521_, _09179_, _09048_);
  not (_23522_, _23478_);
  nor (_23523_, _23522_, _09165_);
  and (_23524_, _09163_, \oc8051_golden_model_1.PC [11]);
  and (_23525_, _23524_, _09168_);
  or (_23526_, _23525_, _23523_);
  and (_23528_, _23526_, _02546_);
  or (_23529_, _23528_, _23521_);
  and (_23530_, _23529_, _23520_);
  and (_23531_, _09048_, _02934_);
  or (_23532_, _23531_, _07428_);
  or (_23533_, _23532_, _23530_);
  nand (_23534_, _23522_, _07428_);
  and (_23535_, _23534_, _02544_);
  and (_23536_, _23535_, _23533_);
  or (_23537_, _23536_, _23518_);
  and (_23539_, _23537_, _21080_);
  nand (_23540_, _23478_, _07425_);
  nand (_23541_, _23540_, _05325_);
  or (_23542_, _23541_, _23539_);
  and (_23543_, _23542_, _09188_);
  and (_23544_, _23543_, _23517_);
  or (_23545_, _23544_, _23508_);
  and (_23546_, _23545_, _09018_);
  and (_23547_, _23478_, _09194_);
  or (_23548_, _23547_, _09193_);
  or (_23550_, _23548_, _23546_);
  and (_23551_, _23550_, _23503_);
  or (_23552_, _23551_, _09200_);
  or (_23553_, _23478_, _09199_);
  and (_23554_, _23553_, _02943_);
  and (_23555_, _23554_, _23552_);
  and (_23556_, _09048_, _02928_);
  or (_23557_, _23556_, _09206_);
  or (_23558_, _23557_, _23555_);
  nand (_23559_, _23522_, _09206_);
  and (_23561_, _23559_, _09211_);
  and (_23562_, _23561_, _23558_);
  or (_23563_, _09211_, _09049_);
  nand (_23564_, _23563_, _09217_);
  or (_23565_, _23564_, _23562_);
  or (_23566_, _23493_, _09252_);
  nand (_23567_, _09252_, _08859_);
  and (_23568_, _23567_, _23566_);
  or (_23569_, _23568_, _09217_);
  and (_23570_, _23569_, _02973_);
  and (_23572_, _23570_, _23565_);
  or (_23573_, _23572_, _23502_);
  or (_23574_, _23573_, _23498_);
  and (_23575_, _23574_, _08969_);
  or (_23576_, _23493_, _08839_);
  nand (_23577_, _08859_, _08839_);
  and (_23578_, _23577_, _02979_);
  and (_23579_, _23578_, _23576_);
  or (_23580_, _23579_, _23575_);
  and (_23581_, _23580_, _08828_);
  nand (_23583_, _23478_, _08827_);
  nand (_23584_, _23583_, _09267_);
  or (_23585_, _23584_, _23581_);
  or (_23586_, _09267_, _09048_);
  and (_23587_, _23586_, _09273_);
  and (_23588_, _23587_, _23585_);
  nor (_23589_, _23522_, _09273_);
  or (_23590_, _23589_, _09280_);
  or (_23591_, _23590_, _23588_);
  or (_23592_, _09279_, _09048_);
  and (_23594_, _23592_, _09285_);
  and (_23595_, _23594_, _23591_);
  nor (_23596_, _23522_, _09285_);
  or (_23597_, _23596_, _09290_);
  or (_23598_, _23597_, _23595_);
  or (_23599_, _09289_, _09048_);
  and (_23600_, _23599_, _02499_);
  and (_23601_, _23600_, _23598_);
  and (_23602_, _23522_, _09298_);
  nor (_23603_, _23602_, _10331_);
  or (_23605_, _23603_, _23601_);
  or (_23606_, _09298_, _09048_);
  and (_23607_, _23606_, _08194_);
  and (_23608_, _23607_, _23605_);
  nand (_23609_, _08858_, _02975_);
  nand (_23610_, _23609_, _09305_);
  or (_23611_, _23610_, _23608_);
  or (_23612_, _09305_, _09048_);
  and (_23613_, _23612_, _02970_);
  and (_23614_, _23613_, _23611_);
  nor (_23616_, _08858_, _08824_);
  nor (_23617_, _23616_, _10325_);
  or (_23618_, _23617_, _23614_);
  nand (_23619_, _23522_, _08824_);
  and (_23620_, _23619_, _23618_);
  or (_23621_, _23620_, _09316_);
  or (_23622_, _09315_, _09048_);
  and (_23623_, _23622_, _09319_);
  and (_23624_, _23623_, _23621_);
  and (_23625_, _23513_, _09318_);
  or (_23627_, _23625_, _05516_);
  or (_23628_, _23627_, _23624_);
  and (_23629_, _23628_, _23489_);
  or (_23630_, _23629_, _02974_);
  nand (_23631_, _08859_, _02974_);
  and (_23632_, _23631_, _07808_);
  and (_23633_, _23632_, _23630_);
  and (_23634_, _09048_, _07807_);
  or (_23635_, _23634_, _23633_);
  and (_23636_, _23635_, _09335_);
  nor (_23638_, _09362_, \oc8051_golden_model_1.DPH [3]);
  nor (_23639_, _23638_, _09363_);
  and (_23640_, _23639_, _09334_);
  or (_23641_, _23640_, _09372_);
  or (_23642_, _23641_, _23636_);
  or (_23643_, _09371_, _09048_);
  and (_23644_, _23643_, _09376_);
  and (_23645_, _23644_, _23642_);
  or (_23646_, _23513_, _08149_);
  or (_23647_, _09048_, _09381_);
  and (_23649_, _23647_, _09375_);
  and (_23650_, _23649_, _23646_);
  or (_23651_, _23650_, _09385_);
  or (_23652_, _23651_, _23645_);
  and (_23653_, _23652_, _23488_);
  or (_23654_, _23653_, _08815_);
  or (_23655_, _08814_, _09048_);
  and (_23656_, _23655_, _07092_);
  and (_23657_, _23656_, _23654_);
  nand (_23658_, _08858_, _02977_);
  nand (_23660_, _23658_, _09394_);
  or (_23661_, _23660_, _23657_);
  or (_23662_, _09394_, _09048_);
  and (_23663_, _23662_, _09398_);
  and (_23664_, _23663_, _23661_);
  or (_23665_, _23513_, _09381_);
  or (_23666_, _09048_, _08149_);
  and (_23667_, _23666_, _09397_);
  and (_23668_, _23667_, _23665_);
  or (_23669_, _23668_, _23664_);
  and (_23671_, _23669_, _08812_);
  nor (_23672_, _23522_, _08812_);
  or (_23673_, _23672_, _07882_);
  or (_23674_, _23673_, _23671_);
  or (_23675_, _09048_, _07881_);
  and (_23676_, _23675_, _03881_);
  and (_23677_, _23676_, _23674_);
  nand (_23678_, _08858_, _02991_);
  nand (_23679_, _23678_, _08809_);
  or (_23680_, _23679_, _23677_);
  and (_23682_, _23680_, _23487_);
  or (_23683_, _23513_, \oc8051_golden_model_1.PSW [7]);
  or (_23684_, _09048_, _07294_);
  and (_23685_, _23684_, _08807_);
  and (_23686_, _23685_, _23683_);
  or (_23687_, _23686_, _09418_);
  or (_23688_, _23687_, _23682_);
  and (_23689_, _23688_, _23485_);
  or (_23690_, _23689_, _07901_);
  or (_23691_, _09048_, _07900_);
  and (_23693_, _23691_, _07120_);
  and (_23694_, _23693_, _23690_);
  nand (_23695_, _08858_, _02994_);
  nand (_23696_, _23695_, _08801_);
  or (_23697_, _23696_, _23694_);
  and (_23698_, _23697_, _23484_);
  or (_23699_, _23513_, _07294_);
  or (_23700_, _09048_, \oc8051_golden_model_1.PSW [7]);
  and (_23701_, _23700_, _08799_);
  and (_23702_, _23701_, _23699_);
  or (_23704_, _23702_, _09434_);
  or (_23705_, _23704_, _23698_);
  and (_23706_, _23705_, _23481_);
  or (_23707_, _23706_, _07948_);
  or (_23708_, _09048_, _07947_);
  and (_23709_, _23708_, _08028_);
  and (_23710_, _23709_, _23707_);
  and (_23711_, _23478_, _08027_);
  or (_23712_, _23711_, _03113_);
  or (_23713_, _23712_, _23710_);
  nand (_23715_, _04226_, _03113_);
  and (_23716_, _23715_, _23713_);
  or (_23717_, _23716_, _02592_);
  nand (_23718_, _09049_, _02592_);
  and (_23719_, _23718_, _03549_);
  and (_23720_, _23719_, _23717_);
  or (_23721_, _23493_, _09641_);
  or (_23722_, _09640_, _08858_);
  and (_23723_, _23722_, _02993_);
  and (_23724_, _23723_, _23721_);
  or (_23726_, _23724_, _09455_);
  or (_23727_, _23726_, _23720_);
  and (_23728_, _23727_, _23480_);
  or (_23729_, _23728_, _08772_);
  nand (_23730_, _09049_, _08772_);
  and (_23731_, _23730_, _09650_);
  and (_23732_, _23731_, _23729_);
  and (_23733_, _23478_, _07143_);
  or (_23734_, _23733_, _02854_);
  or (_23735_, _23734_, _23732_);
  nand (_23737_, _04226_, _02854_);
  and (_23738_, _23737_, _23735_);
  or (_23739_, _23738_, _02575_);
  nand (_23740_, _09049_, _02575_);
  and (_23741_, _23740_, _03134_);
  and (_23742_, _23741_, _23739_);
  or (_23743_, _23493_, _09640_);
  nand (_23744_, _09640_, _08859_);
  and (_23745_, _23744_, _23743_);
  and (_23746_, _23745_, _02990_);
  or (_23748_, _23746_, _09668_);
  or (_23749_, _23748_, _23742_);
  or (_23750_, _23478_, _09667_);
  and (_23751_, _23750_, _03138_);
  and (_23752_, _23751_, _23749_);
  nand (_23753_, _09048_, _03133_);
  nand (_23754_, _23753_, _09675_);
  or (_23755_, _23754_, _23752_);
  or (_23756_, _23478_, _09675_);
  and (_23757_, _23756_, _05219_);
  and (_23759_, _23757_, _23755_);
  and (_23760_, _02988_, _02774_);
  or (_23761_, _23760_, _02572_);
  or (_23762_, _23761_, _23759_);
  nand (_23763_, _09049_, _02572_);
  and (_23764_, _23763_, _03142_);
  and (_23765_, _23764_, _23762_);
  and (_23766_, _23745_, _02778_);
  or (_23767_, _23766_, _09689_);
  or (_23768_, _23767_, _23765_);
  or (_23770_, _23478_, _09688_);
  and (_23771_, _23770_, _02853_);
  and (_23772_, _23771_, _23768_);
  nand (_23773_, _09048_, _02852_);
  nand (_23774_, _23773_, _09696_);
  or (_23775_, _23774_, _23772_);
  or (_23776_, _23478_, _09696_);
  and (_23777_, _23776_, _09699_);
  and (_23778_, _23777_, _23775_);
  and (_23779_, _02982_, _02774_);
  or (_23781_, _23779_, _02568_);
  or (_23782_, _23781_, _23778_);
  nand (_23783_, _09049_, _02568_);
  and (_23784_, _23783_, _09707_);
  and (_23785_, _23784_, _23782_);
  or (_23786_, _23785_, _23479_);
  or (_23787_, _23786_, _34450_);
  or (_23788_, _34446_, \oc8051_golden_model_1.PC [11]);
  and (_23789_, _23788_, _35583_);
  and (_35629_[11], _23789_, _23787_);
  nand (_23791_, _09044_, _02852_);
  nor (_23792_, _08778_, \oc8051_golden_model_1.PC [12]);
  nor (_23793_, _23792_, _08779_);
  not (_23794_, _23793_);
  and (_23795_, _23794_, _07143_);
  nor (_23796_, _09371_, _09044_);
  and (_23797_, _08952_, _08949_);
  nor (_23798_, _23797_, _08953_);
  not (_23799_, _23798_);
  or (_23800_, _23799_, _09000_);
  nand (_23802_, _09000_, _08853_);
  and (_23803_, _23802_, _23800_);
  or (_23804_, _23803_, _09858_);
  and (_23805_, _09044_, _02928_);
  or (_23806_, _09148_, _09044_);
  nor (_23807_, _09131_, _09129_);
  nor (_23808_, _23807_, _09132_);
  nand (_23809_, _23808_, _09148_);
  and (_23810_, _23809_, _23806_);
  and (_23811_, _23810_, _05327_);
  or (_23813_, _23794_, _09165_);
  or (_23814_, _09044_, _02546_);
  nand (_23815_, _09043_, _02837_);
  nand (_23816_, _09168_, \oc8051_golden_model_1.PC [12]);
  and (_23817_, _23816_, _23815_);
  nand (_23818_, _09163_, _02546_);
  or (_23819_, _23818_, _23817_);
  and (_23820_, _23819_, _23814_);
  or (_23821_, _23820_, _20340_);
  and (_23822_, _23821_, _07406_);
  and (_23824_, _23822_, _23813_);
  and (_23825_, _09044_, _02934_);
  or (_23826_, _23825_, _07428_);
  or (_23827_, _23826_, _23824_);
  nand (_23828_, _23793_, _07428_);
  and (_23829_, _23828_, _02544_);
  and (_23830_, _23829_, _23827_);
  and (_23831_, _09044_, _09178_);
  or (_23832_, _23831_, _07425_);
  or (_23833_, _23832_, _23830_);
  nand (_23835_, _23793_, _07425_);
  and (_23836_, _23835_, _05325_);
  and (_23837_, _23836_, _23833_);
  or (_23838_, _23837_, _23811_);
  and (_23839_, _23838_, _05311_);
  and (_23840_, _23794_, _03806_);
  or (_23841_, _23840_, _02932_);
  or (_23842_, _23841_, _23839_);
  and (_23843_, _23799_, _09023_);
  or (_23844_, _23843_, _06162_);
  and (_23846_, _19708_, _08854_);
  or (_23847_, _23846_, _23844_);
  and (_23848_, _23847_, _09018_);
  and (_23849_, _23848_, _23842_);
  nor (_23850_, _23793_, _09018_);
  or (_23851_, _23850_, _23849_);
  and (_23852_, _23851_, _09015_);
  or (_23853_, _09015_, _09043_);
  nand (_23854_, _23853_, _09199_);
  or (_23855_, _23854_, _23852_);
  or (_23857_, _23794_, _09199_);
  and (_23858_, _23857_, _02943_);
  and (_23859_, _23858_, _23855_);
  or (_23860_, _23859_, _23805_);
  and (_23861_, _23860_, _09212_);
  nand (_23862_, _23794_, _09206_);
  nand (_23863_, _23862_, _09211_);
  or (_23864_, _23863_, _23861_);
  or (_23865_, _09211_, _09044_);
  and (_23866_, _23865_, _09217_);
  and (_23868_, _23866_, _23864_);
  nand (_23869_, _09252_, _08853_);
  or (_23870_, _23799_, _09252_);
  and (_23871_, _23870_, _23869_);
  and (_23872_, _23871_, _09906_);
  or (_23873_, _23872_, _02972_);
  or (_23874_, _23873_, _23868_);
  and (_23875_, _23874_, _03397_);
  and (_23876_, _23875_, _23804_);
  or (_23877_, _23799_, _09008_);
  nand (_23879_, _09008_, _08853_);
  and (_23880_, _23879_, _02944_);
  and (_23881_, _23880_, _23877_);
  or (_23882_, _23881_, _02979_);
  or (_23883_, _23882_, _23876_);
  nor (_23884_, _23798_, _08839_);
  and (_23885_, _08854_, _08839_);
  or (_23886_, _23885_, _08969_);
  or (_23887_, _23886_, _23884_);
  and (_23888_, _23887_, _08828_);
  and (_23890_, _23888_, _23883_);
  and (_23891_, _23793_, _09267_);
  nor (_23892_, _23891_, _10341_);
  or (_23893_, _23892_, _23890_);
  or (_23894_, _09267_, _09044_);
  and (_23895_, _23894_, _09273_);
  and (_23896_, _23895_, _23893_);
  nor (_23897_, _23793_, _09273_);
  or (_23898_, _23897_, _09280_);
  or (_23899_, _23898_, _23896_);
  or (_23901_, _09279_, _09044_);
  and (_23902_, _23901_, _09285_);
  and (_23903_, _23902_, _23899_);
  nor (_23904_, _23793_, _09285_);
  or (_23905_, _23904_, _09290_);
  or (_23906_, _23905_, _23903_);
  or (_23907_, _09289_, _09044_);
  and (_23908_, _23907_, _02499_);
  and (_23909_, _23908_, _23906_);
  and (_23910_, _23793_, _09298_);
  nor (_23912_, _23910_, _10331_);
  or (_23913_, _23912_, _23909_);
  or (_23914_, _09298_, _09044_);
  and (_23915_, _23914_, _08194_);
  and (_23916_, _23915_, _23913_);
  and (_23917_, _09305_, _08853_);
  nor (_23918_, _23917_, _10308_);
  or (_23919_, _23918_, _23916_);
  or (_23920_, _09305_, _09044_);
  and (_23921_, _23920_, _02970_);
  and (_23923_, _23921_, _23919_);
  nor (_23924_, _08854_, _08824_);
  nor (_23925_, _23924_, _10325_);
  nor (_23926_, _23925_, _23923_);
  nand (_23927_, _23793_, _08824_);
  nand (_23928_, _23927_, _09315_);
  or (_23929_, _23928_, _23926_);
  or (_23930_, _09315_, _09043_);
  and (_23931_, _23930_, _09319_);
  and (_23932_, _23931_, _23929_);
  and (_23934_, _23808_, _09318_);
  or (_23935_, _23934_, _23932_);
  and (_23936_, _23935_, _05267_);
  nor (_23937_, _09044_, _05267_);
  or (_23938_, _23937_, _02974_);
  or (_23939_, _23938_, _23936_);
  nand (_23940_, _08854_, _02974_);
  and (_23941_, _23940_, _07808_);
  and (_23942_, _23941_, _23939_);
  and (_23943_, _09043_, _07807_);
  or (_23945_, _23943_, _09334_);
  or (_23946_, _23945_, _23942_);
  nor (_23947_, _09363_, \oc8051_golden_model_1.DPH [4]);
  nor (_23948_, _23947_, _09364_);
  or (_23949_, _23948_, _09335_);
  and (_23950_, _23949_, _09371_);
  and (_23951_, _23950_, _23946_);
  or (_23952_, _23951_, _23796_);
  and (_23953_, _23952_, _10350_);
  or (_23954_, _23808_, _08149_);
  or (_23956_, _09043_, _09381_);
  and (_23957_, _23956_, _09375_);
  and (_23958_, _23957_, _23954_);
  nor (_23959_, _23794_, _08822_);
  or (_23960_, _23959_, _23958_);
  or (_23961_, _23960_, _23953_);
  and (_23962_, _23961_, _08814_);
  nor (_23963_, _08814_, _09044_);
  or (_23964_, _23963_, _02977_);
  or (_23965_, _23964_, _23962_);
  nand (_23967_, _08854_, _02977_);
  and (_23968_, _23967_, _09394_);
  and (_23969_, _23968_, _23965_);
  nor (_23970_, _09394_, _09044_);
  or (_23971_, _23970_, _23969_);
  and (_23972_, _23971_, _10355_);
  nor (_23973_, _23794_, _08812_);
  or (_23974_, _23808_, _09381_);
  or (_23975_, _09043_, _08149_);
  and (_23976_, _23975_, _09397_);
  and (_23978_, _23976_, _23974_);
  or (_23979_, _23978_, _23973_);
  or (_23980_, _23979_, _23972_);
  and (_23981_, _23980_, _07881_);
  nor (_23982_, _09044_, _07881_);
  or (_23983_, _23982_, _02991_);
  or (_23984_, _23983_, _23981_);
  nand (_23985_, _08854_, _02991_);
  and (_23986_, _23985_, _08809_);
  and (_23987_, _23986_, _23984_);
  nor (_23989_, _09044_, _08809_);
  or (_23990_, _23989_, _23987_);
  and (_23991_, _23990_, _10379_);
  nor (_23992_, _23794_, _08805_);
  or (_23993_, _23808_, \oc8051_golden_model_1.PSW [7]);
  or (_23994_, _09043_, _07294_);
  and (_23995_, _23994_, _08807_);
  and (_23996_, _23995_, _23993_);
  or (_23997_, _23996_, _23992_);
  or (_23998_, _23997_, _23991_);
  and (_23999_, _23998_, _07900_);
  nor (_24000_, _09044_, _07900_);
  or (_24001_, _24000_, _02994_);
  or (_24002_, _24001_, _23999_);
  nand (_24003_, _08854_, _02994_);
  and (_24004_, _24003_, _08801_);
  and (_24005_, _24004_, _24002_);
  nor (_24006_, _09044_, _08801_);
  or (_24007_, _24006_, _24005_);
  nand (_24008_, _24007_, _10376_);
  or (_24010_, _23808_, _07294_);
  or (_24011_, _09043_, \oc8051_golden_model_1.PSW [7]);
  and (_24012_, _24011_, _08799_);
  and (_24013_, _24012_, _24010_);
  nor (_24014_, _23794_, _08797_);
  or (_24015_, _24014_, _07948_);
  nor (_24016_, _24015_, _24013_);
  and (_24017_, _24016_, _24008_);
  nor (_24018_, _09043_, _07947_);
  or (_24019_, _24018_, _08027_);
  or (_24021_, _24019_, _24017_);
  nand (_24022_, _23793_, _08027_);
  and (_24023_, _24022_, _24021_);
  or (_24024_, _24023_, _03113_);
  or (_24025_, _05143_, _10159_);
  and (_24026_, _24025_, _05741_);
  and (_24027_, _24026_, _24024_);
  and (_24028_, _09044_, _02592_);
  or (_24029_, _24028_, _02993_);
  or (_24030_, _24029_, _24027_);
  nor (_24032_, _09640_, _08853_);
  and (_24033_, _23799_, _09640_);
  or (_24034_, _24033_, _03549_);
  or (_24035_, _24034_, _24032_);
  and (_24036_, _24035_, _08795_);
  and (_24037_, _24036_, _24030_);
  nor (_24038_, _23794_, _08772_);
  nor (_24039_, _24038_, _10297_);
  or (_24040_, _24039_, _24037_);
  nand (_24041_, _09043_, _08772_);
  and (_24043_, _24041_, _09650_);
  and (_24044_, _24043_, _24040_);
  or (_24045_, _24044_, _23795_);
  and (_24046_, _24045_, _02855_);
  and (_24047_, _05143_, _02854_);
  or (_24048_, _24047_, _02575_);
  or (_24049_, _24048_, _24046_);
  nand (_24050_, _09043_, _02575_);
  and (_24051_, _24050_, _03134_);
  and (_24052_, _24051_, _24049_);
  and (_24054_, _09640_, _08854_);
  nor (_24055_, _23798_, _09640_);
  nor (_24056_, _24055_, _24054_);
  nor (_24057_, _24056_, _03134_);
  or (_24058_, _24057_, _24052_);
  nand (_24059_, _24058_, _09667_);
  or (_24060_, _23793_, _09667_);
  and (_24061_, _24060_, _24059_);
  or (_24062_, _24061_, _03133_);
  nand (_24063_, _09044_, _03133_);
  and (_24065_, _24063_, _09675_);
  and (_24066_, _24065_, _24062_);
  or (_24067_, _23794_, _09675_);
  nand (_24068_, _24067_, _05219_);
  or (_24069_, _24068_, _24066_);
  nand (_24070_, _03620_, _02988_);
  and (_24071_, _24070_, _05218_);
  and (_24072_, _24071_, _24069_);
  and (_24073_, _09043_, _02572_);
  or (_24074_, _24073_, _02778_);
  or (_24077_, _24074_, _24072_);
  or (_24078_, _24056_, _03142_);
  and (_24079_, _24078_, _09688_);
  and (_24080_, _24079_, _24077_);
  nor (_24081_, _23794_, _09688_);
  or (_24082_, _24081_, _02852_);
  or (_24083_, _24082_, _24080_);
  and (_24084_, _24083_, _23791_);
  nor (_24085_, _24084_, _21033_);
  nor (_24086_, _23793_, _09696_);
  nor (_24088_, _24086_, _02982_);
  not (_24089_, _24088_);
  nor (_24090_, _24089_, _24085_);
  nor (_24091_, _03620_, _09699_);
  or (_24092_, _24091_, _02568_);
  nor (_24093_, _24092_, _24090_);
  and (_24094_, _09044_, _02568_);
  nor (_24095_, _24094_, _24093_);
  and (_24096_, _24095_, _09707_);
  and (_24097_, _23793_, _09706_);
  or (_24099_, _24097_, _24096_);
  or (_24100_, _24099_, _34450_);
  or (_24101_, _34446_, \oc8051_golden_model_1.PC [12]);
  and (_24102_, _24101_, _35583_);
  and (_35629_[12], _24102_, _24100_);
  not (_24103_, \oc8051_golden_model_1.PC [13]);
  and (_24104_, _08776_, _06138_);
  and (_24105_, _24104_, \oc8051_golden_model_1.PC [12]);
  nor (_24106_, _24105_, _24103_);
  and (_24107_, _24105_, _24103_);
  or (_24109_, _24107_, _24106_);
  or (_24110_, _24109_, _08795_);
  or (_24111_, _24109_, _08797_);
  or (_24112_, _09037_, _08801_);
  and (_24113_, _24112_, _08800_);
  or (_24114_, _24109_, _08805_);
  or (_24115_, _09037_, _08809_);
  and (_24116_, _24115_, _08808_);
  or (_24117_, _09039_, _09040_);
  nand (_24118_, _24117_, _09133_);
  or (_24120_, _24117_, _09133_);
  and (_24121_, _24120_, _24118_);
  or (_24122_, _24121_, _09381_);
  or (_24123_, _09037_, _08149_);
  and (_24124_, _24123_, _09397_);
  and (_24125_, _24124_, _24122_);
  or (_24126_, _24109_, _08822_);
  or (_24127_, _09037_, _05267_);
  and (_24128_, _09000_, _08848_);
  or (_24129_, _08851_, _08850_);
  nand (_24131_, _24129_, _08954_);
  or (_24132_, _24129_, _08954_);
  and (_24133_, _24132_, _24131_);
  and (_24134_, _24133_, _23254_);
  or (_24135_, _24134_, _09858_);
  or (_24136_, _24135_, _24128_);
  or (_24137_, _24133_, _09252_);
  nand (_24138_, _09252_, _08849_);
  and (_24139_, _24138_, _24137_);
  or (_24140_, _24139_, _09217_);
  or (_24142_, _09015_, _09037_);
  or (_24143_, _09023_, _08848_);
  or (_24144_, _24133_, _09025_);
  and (_24145_, _24144_, _02932_);
  and (_24146_, _24145_, _24143_);
  and (_24147_, _09150_, _09037_);
  and (_24148_, _24121_, _09148_);
  or (_24149_, _24148_, _24147_);
  or (_24150_, _24149_, _05325_);
  and (_24151_, _09037_, _09178_);
  or (_24153_, _24109_, _09159_);
  and (_24154_, _24153_, _07406_);
  and (_24155_, _09179_, _09037_);
  not (_24156_, _24109_);
  nor (_24157_, _24156_, _09165_);
  and (_24158_, _09163_, \oc8051_golden_model_1.PC [13]);
  and (_24159_, _24158_, _09168_);
  or (_24160_, _24159_, _24157_);
  and (_24161_, _24160_, _02546_);
  or (_24162_, _24161_, _24155_);
  and (_24164_, _24162_, _24154_);
  and (_24165_, _09037_, _02934_);
  or (_24166_, _24165_, _07428_);
  or (_24167_, _24166_, _24164_);
  nand (_24168_, _24156_, _07428_);
  and (_24169_, _24168_, _02544_);
  and (_24170_, _24169_, _24167_);
  or (_24171_, _24170_, _24151_);
  and (_24172_, _24171_, _21080_);
  nand (_24173_, _24109_, _07425_);
  nand (_24175_, _24173_, _05325_);
  or (_24176_, _24175_, _24172_);
  and (_24177_, _24176_, _09188_);
  and (_24178_, _24177_, _24150_);
  or (_24179_, _24178_, _24146_);
  and (_24180_, _24179_, _09018_);
  and (_24181_, _24109_, _09194_);
  or (_24182_, _24181_, _09193_);
  or (_24183_, _24182_, _24180_);
  and (_24184_, _24183_, _24142_);
  or (_24186_, _24184_, _09200_);
  or (_24187_, _24109_, _09199_);
  and (_24188_, _24187_, _02943_);
  and (_24189_, _24188_, _24186_);
  and (_24190_, _09037_, _02928_);
  or (_24191_, _24190_, _09206_);
  or (_24192_, _24191_, _24189_);
  nand (_24193_, _24156_, _09206_);
  and (_24194_, _24193_, _09211_);
  and (_24195_, _24194_, _24192_);
  or (_24197_, _09211_, _09038_);
  nand (_24198_, _24197_, _09217_);
  or (_24199_, _24198_, _24195_);
  and (_24200_, _24199_, _24140_);
  or (_24201_, _24200_, _02972_);
  and (_24202_, _24201_, _09927_);
  and (_24203_, _24202_, _24136_);
  or (_24204_, _24133_, _08839_);
  nand (_24205_, _08849_, _08839_);
  and (_24206_, _24205_, _02979_);
  and (_24208_, _24206_, _24204_);
  and (_24209_, _24133_, _09009_);
  and (_24210_, _09008_, _08848_);
  or (_24211_, _24210_, _24209_);
  and (_24212_, _24211_, _02944_);
  or (_24213_, _24212_, _24208_);
  or (_24214_, _24213_, _24203_);
  and (_24215_, _24214_, _08828_);
  nand (_24216_, _24109_, _08827_);
  nand (_24217_, _24216_, _09267_);
  or (_24219_, _24217_, _24215_);
  or (_24220_, _09267_, _09037_);
  and (_24221_, _24220_, _09273_);
  and (_24222_, _24221_, _24219_);
  nor (_24223_, _24156_, _09273_);
  or (_24224_, _24223_, _09280_);
  or (_24225_, _24224_, _24222_);
  or (_24226_, _09279_, _09037_);
  and (_24227_, _24226_, _09285_);
  and (_24228_, _24227_, _24225_);
  nor (_24230_, _24156_, _09285_);
  or (_24231_, _24230_, _09290_);
  or (_24232_, _24231_, _24228_);
  or (_24233_, _09289_, _09037_);
  and (_24234_, _24233_, _02499_);
  and (_24235_, _24234_, _24232_);
  and (_24236_, _24156_, _09298_);
  nor (_24237_, _24236_, _10331_);
  or (_24238_, _24237_, _24235_);
  or (_24239_, _09298_, _09037_);
  and (_24241_, _24239_, _08194_);
  and (_24242_, _24241_, _24238_);
  nand (_24243_, _08848_, _02975_);
  nand (_24244_, _24243_, _09305_);
  or (_24245_, _24244_, _24242_);
  or (_24246_, _09305_, _09037_);
  and (_24247_, _24246_, _02970_);
  and (_24248_, _24247_, _24245_);
  nor (_24249_, _08848_, _08824_);
  nor (_24250_, _24249_, _10325_);
  or (_24252_, _24250_, _24248_);
  nand (_24253_, _24156_, _08824_);
  and (_24254_, _24253_, _24252_);
  or (_24255_, _24254_, _09316_);
  or (_24256_, _09315_, _09037_);
  and (_24257_, _24256_, _09319_);
  and (_24258_, _24257_, _24255_);
  and (_24259_, _24121_, _09318_);
  or (_24260_, _24259_, _05516_);
  or (_24261_, _24260_, _24258_);
  and (_24263_, _24261_, _24127_);
  or (_24264_, _24263_, _02974_);
  nand (_24265_, _08849_, _02974_);
  and (_24266_, _24265_, _07808_);
  and (_24267_, _24266_, _24264_);
  and (_24268_, _09037_, _07807_);
  or (_24269_, _24268_, _24267_);
  and (_24270_, _24269_, _09335_);
  nor (_24271_, _09364_, \oc8051_golden_model_1.DPH [5]);
  nor (_24272_, _24271_, _09365_);
  and (_24274_, _24272_, _09334_);
  or (_24275_, _24274_, _09372_);
  or (_24276_, _24275_, _24270_);
  or (_24277_, _09371_, _09037_);
  and (_24278_, _24277_, _09376_);
  and (_24279_, _24278_, _24276_);
  or (_24280_, _24121_, _08149_);
  or (_24281_, _09037_, _09381_);
  and (_24282_, _24281_, _09375_);
  and (_24283_, _24282_, _24280_);
  or (_24285_, _24283_, _09385_);
  or (_24286_, _24285_, _24279_);
  and (_24287_, _24286_, _24126_);
  or (_24288_, _24287_, _08815_);
  or (_24289_, _08814_, _09037_);
  and (_24290_, _24289_, _07092_);
  and (_24291_, _24290_, _24288_);
  nand (_24292_, _08848_, _02977_);
  nand (_24293_, _24292_, _09394_);
  or (_24294_, _24293_, _24291_);
  or (_24296_, _09394_, _09037_);
  and (_24297_, _24296_, _09398_);
  and (_24298_, _24297_, _24294_);
  or (_24299_, _24298_, _24125_);
  and (_24300_, _24299_, _08812_);
  nor (_24301_, _24156_, _08812_);
  or (_24302_, _24301_, _07882_);
  or (_24303_, _24302_, _24300_);
  or (_24304_, _09037_, _07881_);
  and (_24305_, _24304_, _03881_);
  and (_24307_, _24305_, _24303_);
  nand (_24308_, _08848_, _02991_);
  nand (_24309_, _24308_, _08809_);
  or (_24310_, _24309_, _24307_);
  and (_24311_, _24310_, _24116_);
  or (_24312_, _24121_, \oc8051_golden_model_1.PSW [7]);
  or (_24313_, _09037_, _07294_);
  and (_24314_, _24313_, _08807_);
  and (_24315_, _24314_, _24312_);
  or (_24316_, _24315_, _09418_);
  or (_24318_, _24316_, _24311_);
  and (_24319_, _24318_, _24114_);
  or (_24320_, _24319_, _07901_);
  or (_24321_, _09037_, _07900_);
  and (_24322_, _24321_, _07120_);
  and (_24323_, _24322_, _24320_);
  nand (_24324_, _08848_, _02994_);
  nand (_24325_, _24324_, _08801_);
  or (_24326_, _24325_, _24323_);
  and (_24327_, _24326_, _24113_);
  or (_24329_, _24121_, _07294_);
  or (_24330_, _09037_, \oc8051_golden_model_1.PSW [7]);
  and (_24331_, _24330_, _08799_);
  and (_24332_, _24331_, _24329_);
  or (_24333_, _24332_, _09434_);
  or (_24334_, _24333_, _24327_);
  and (_24335_, _24334_, _24111_);
  or (_24336_, _24335_, _07948_);
  or (_24337_, _09037_, _07947_);
  and (_24338_, _24337_, _08028_);
  and (_24340_, _24338_, _24336_);
  and (_24341_, _24109_, _08027_);
  or (_24342_, _24341_, _03113_);
  or (_24343_, _24342_, _24340_);
  nand (_24344_, _04839_, _03113_);
  and (_24345_, _24344_, _24343_);
  or (_24346_, _24345_, _02592_);
  nand (_24347_, _09038_, _02592_);
  and (_24348_, _24347_, _03549_);
  and (_24349_, _24348_, _24346_);
  or (_24351_, _24133_, _09641_);
  or (_24352_, _09640_, _08848_);
  and (_24353_, _24352_, _02993_);
  and (_24354_, _24353_, _24351_);
  or (_24355_, _24354_, _09455_);
  or (_24356_, _24355_, _24349_);
  and (_24357_, _24356_, _24110_);
  or (_24358_, _24357_, _08772_);
  nand (_24359_, _09038_, _08772_);
  and (_24360_, _24359_, _09650_);
  and (_24362_, _24360_, _24358_);
  and (_24363_, _24109_, _07143_);
  or (_24364_, _24363_, _02854_);
  or (_24365_, _24364_, _24362_);
  nand (_24366_, _04839_, _02854_);
  and (_24367_, _24366_, _24365_);
  or (_24368_, _24367_, _02575_);
  nand (_24369_, _09038_, _02575_);
  and (_24370_, _24369_, _03134_);
  and (_24371_, _24370_, _24368_);
  or (_24373_, _24133_, _09640_);
  nand (_24374_, _09640_, _08849_);
  and (_24375_, _24374_, _24373_);
  and (_24376_, _24375_, _02990_);
  or (_24377_, _24376_, _09668_);
  or (_24378_, _24377_, _24371_);
  or (_24379_, _24109_, _09667_);
  and (_24380_, _24379_, _03138_);
  and (_24381_, _24380_, _24378_);
  nand (_24382_, _09037_, _03133_);
  nand (_24384_, _24382_, _09675_);
  or (_24385_, _24384_, _24381_);
  or (_24386_, _24109_, _09675_);
  and (_24387_, _24386_, _05219_);
  and (_24388_, _24387_, _24385_);
  nor (_24389_, _03179_, _05219_);
  or (_24390_, _24389_, _02572_);
  or (_24391_, _24390_, _24388_);
  nand (_24392_, _09038_, _02572_);
  and (_24393_, _24392_, _03142_);
  and (_24395_, _24393_, _24391_);
  and (_24396_, _24375_, _02778_);
  or (_24397_, _24396_, _09689_);
  or (_24398_, _24397_, _24395_);
  or (_24399_, _24109_, _09688_);
  and (_24400_, _24399_, _02853_);
  and (_24401_, _24400_, _24398_);
  nand (_24402_, _09037_, _02852_);
  nand (_24403_, _24402_, _09696_);
  or (_24404_, _24403_, _24401_);
  or (_24406_, _24109_, _09696_);
  and (_24407_, _24406_, _09699_);
  and (_24408_, _24407_, _24404_);
  nand (_24409_, _03179_, _02569_);
  and (_24410_, _24409_, _19634_);
  or (_24411_, _24410_, _24408_);
  nand (_24412_, _09038_, _02568_);
  and (_24413_, _24412_, _09707_);
  and (_24414_, _24413_, _24411_);
  and (_24415_, _24109_, _09706_);
  or (_24417_, _24415_, _24414_);
  or (_24418_, _24417_, _34450_);
  or (_24419_, _34446_, \oc8051_golden_model_1.PC [13]);
  and (_24420_, _24419_, _35583_);
  and (_35629_[13], _24420_, _24418_);
  nand (_24421_, _09031_, _02852_);
  nor (_24422_, _08780_, \oc8051_golden_model_1.PC [14]);
  nor (_24423_, _24422_, _08781_);
  not (_24424_, _24423_);
  and (_24425_, _24424_, _07143_);
  nor (_24427_, _09371_, _09031_);
  or (_24428_, _09030_, _05267_);
  nor (_24429_, _09289_, _09030_);
  nor (_24430_, _24423_, _09273_);
  and (_24431_, _08956_, _08846_);
  nor (_24432_, _24431_, _08957_);
  not (_24433_, _24432_);
  or (_24434_, _24433_, _09000_);
  nand (_24435_, _09000_, _08841_);
  and (_24436_, _24435_, _24434_);
  or (_24438_, _24436_, _09858_);
  nand (_24439_, _24423_, _09206_);
  nor (_24440_, _24423_, _09199_);
  and (_24441_, _09025_, _08842_);
  and (_24442_, _24433_, _09023_);
  or (_24443_, _24442_, _24441_);
  and (_24444_, _24443_, _02932_);
  nand (_24445_, _09165_, _19664_);
  and (_24446_, _24445_, _24423_);
  and (_24447_, _09030_, _02934_);
  and (_24449_, _09179_, _09030_);
  and (_24450_, _02546_, \oc8051_golden_model_1.PC [14]);
  and (_24451_, _24450_, _07406_);
  and (_24452_, _24451_, _09163_);
  and (_24453_, _24452_, _09168_);
  or (_24454_, _24453_, _24449_);
  and (_24455_, _24454_, _09159_);
  or (_24456_, _24455_, _24447_);
  and (_24457_, _24456_, _19664_);
  or (_24458_, _24457_, _09178_);
  nor (_24460_, _24458_, _24446_);
  and (_24461_, _09031_, _09178_);
  or (_24462_, _24461_, _07425_);
  or (_24463_, _24462_, _24460_);
  nand (_24464_, _24423_, _07425_);
  and (_24465_, _24464_, _05325_);
  and (_24466_, _24465_, _24463_);
  and (_24467_, _09135_, _09035_);
  nor (_24468_, _24467_, _09136_);
  nand (_24469_, _24468_, _09148_);
  or (_24471_, _09148_, _09031_);
  and (_24472_, _24471_, _24469_);
  and (_24473_, _24472_, _05327_);
  or (_24474_, _24473_, _24466_);
  and (_24475_, _24474_, _09188_);
  or (_24476_, _24475_, _24444_);
  and (_24477_, _24476_, _09018_);
  and (_24478_, _24424_, _09194_);
  or (_24479_, _24478_, _09193_);
  or (_24480_, _24479_, _24477_);
  or (_24482_, _09015_, _09031_);
  and (_24483_, _24482_, _09199_);
  and (_24484_, _24483_, _24480_);
  or (_24485_, _24484_, _24440_);
  and (_24486_, _24485_, _02943_);
  and (_24487_, _09031_, _02928_);
  or (_24488_, _24487_, _09206_);
  or (_24489_, _24488_, _24486_);
  nand (_24490_, _24489_, _24439_);
  nand (_24491_, _24490_, _09211_);
  or (_24493_, _09211_, _09031_);
  and (_24494_, _24493_, _09217_);
  and (_24495_, _24494_, _24491_);
  nand (_24496_, _09252_, _08841_);
  or (_24497_, _24433_, _09252_);
  and (_24498_, _24497_, _24496_);
  and (_24499_, _24498_, _09906_);
  or (_24500_, _24499_, _02972_);
  or (_24501_, _24500_, _24495_);
  and (_24502_, _24501_, _03397_);
  and (_24504_, _24502_, _24438_);
  or (_24505_, _24433_, _09008_);
  nand (_24506_, _09008_, _08841_);
  and (_24507_, _24506_, _02944_);
  and (_24508_, _24507_, _24505_);
  or (_24509_, _24508_, _02979_);
  or (_24510_, _24509_, _24504_);
  nor (_24511_, _24432_, _08839_);
  and (_24512_, _08842_, _08839_);
  or (_24513_, _24512_, _08969_);
  or (_24515_, _24513_, _24511_);
  and (_24516_, _24515_, _08828_);
  and (_24517_, _24516_, _24510_);
  and (_24518_, _24423_, _09267_);
  nor (_24519_, _24518_, _10341_);
  or (_24520_, _24519_, _24517_);
  or (_24521_, _09267_, _09031_);
  and (_24522_, _24521_, _09273_);
  and (_24523_, _24522_, _24520_);
  or (_24524_, _24523_, _24430_);
  and (_24526_, _24524_, _09279_);
  or (_24527_, _09279_, _09030_);
  nand (_24528_, _24527_, _09285_);
  or (_24529_, _24528_, _24526_);
  or (_24530_, _24424_, _09285_);
  and (_24531_, _24530_, _09289_);
  and (_24532_, _24531_, _24529_);
  or (_24533_, _24532_, _24429_);
  and (_24534_, _24533_, _02499_);
  or (_24535_, _24423_, _02499_);
  nand (_24537_, _24535_, _09298_);
  or (_24538_, _24537_, _24534_);
  or (_24539_, _09298_, _09031_);
  and (_24540_, _24539_, _08194_);
  and (_24541_, _24540_, _24538_);
  and (_24542_, _09305_, _08841_);
  nor (_24543_, _24542_, _10308_);
  or (_24544_, _24543_, _24541_);
  or (_24545_, _09305_, _09031_);
  and (_24546_, _24545_, _02970_);
  and (_24548_, _24546_, _24544_);
  nor (_24549_, _08842_, _08824_);
  nor (_24550_, _24549_, _10325_);
  nor (_24551_, _24550_, _24548_);
  nand (_24552_, _24423_, _08824_);
  nand (_24553_, _24552_, _09315_);
  or (_24554_, _24553_, _24551_);
  or (_24555_, _09315_, _09030_);
  and (_24556_, _24555_, _09319_);
  and (_24557_, _24556_, _24554_);
  and (_24559_, _24468_, _09318_);
  or (_24560_, _24559_, _05516_);
  or (_24561_, _24560_, _24557_);
  and (_24562_, _24561_, _24428_);
  or (_24563_, _24562_, _02974_);
  nand (_24564_, _08842_, _02974_);
  and (_24565_, _24564_, _07808_);
  and (_24566_, _24565_, _24563_);
  and (_24567_, _09030_, _07807_);
  or (_24568_, _24567_, _09334_);
  or (_24570_, _24568_, _24566_);
  nor (_24571_, _09365_, \oc8051_golden_model_1.DPH [6]);
  nor (_24572_, _24571_, _09366_);
  or (_24573_, _24572_, _09335_);
  and (_24574_, _24573_, _09371_);
  and (_24575_, _24574_, _24570_);
  or (_24576_, _24575_, _24427_);
  and (_24577_, _24576_, _10350_);
  or (_24578_, _24468_, _08149_);
  or (_24579_, _09030_, _09381_);
  and (_24581_, _24579_, _09375_);
  and (_24582_, _24581_, _24578_);
  nor (_24583_, _24424_, _08822_);
  or (_24584_, _24583_, _08815_);
  or (_24585_, _24584_, _24582_);
  or (_24586_, _24585_, _24577_);
  or (_24587_, _08814_, _09030_);
  and (_24588_, _24587_, _24586_);
  or (_24589_, _24588_, _02977_);
  nand (_24590_, _08842_, _02977_);
  and (_24592_, _24590_, _09394_);
  and (_24593_, _24592_, _24589_);
  nor (_24594_, _09394_, _09031_);
  or (_24595_, _24594_, _24593_);
  and (_24596_, _24595_, _10355_);
  or (_24597_, _24468_, _09381_);
  or (_24598_, _09030_, _08149_);
  and (_24599_, _24598_, _09397_);
  and (_24600_, _24599_, _24597_);
  nor (_24601_, _24424_, _08812_);
  or (_24603_, _24601_, _24600_);
  or (_24604_, _24603_, _24596_);
  and (_24605_, _24604_, _07881_);
  nor (_24606_, _09031_, _07881_);
  or (_24607_, _24606_, _02991_);
  or (_24608_, _24607_, _24605_);
  nand (_24609_, _08842_, _02991_);
  and (_24610_, _24609_, _08809_);
  and (_24611_, _24610_, _24608_);
  nor (_24612_, _09031_, _08809_);
  or (_24614_, _24612_, _24611_);
  and (_24615_, _24614_, _10379_);
  nor (_24616_, _24424_, _08805_);
  or (_24617_, _24468_, \oc8051_golden_model_1.PSW [7]);
  or (_24618_, _09030_, _07294_);
  and (_24619_, _24618_, _08807_);
  and (_24620_, _24619_, _24617_);
  or (_24621_, _24620_, _24616_);
  or (_24622_, _24621_, _24615_);
  and (_24623_, _24622_, _07900_);
  nor (_24625_, _09031_, _07900_);
  or (_24626_, _24625_, _02994_);
  or (_24627_, _24626_, _24623_);
  nand (_24628_, _08842_, _02994_);
  and (_24629_, _24628_, _08801_);
  and (_24630_, _24629_, _24627_);
  nor (_24631_, _09031_, _08801_);
  or (_24632_, _24631_, _24630_);
  nand (_24633_, _24632_, _10376_);
  or (_24634_, _24468_, _07294_);
  or (_24636_, _09030_, \oc8051_golden_model_1.PSW [7]);
  and (_24637_, _24636_, _08799_);
  and (_24638_, _24637_, _24634_);
  nor (_24639_, _24424_, _08797_);
  or (_24640_, _24639_, _07948_);
  nor (_24641_, _24640_, _24638_);
  and (_24642_, _24641_, _24633_);
  nor (_24643_, _09030_, _07947_);
  or (_24644_, _24643_, _08027_);
  or (_24645_, _24644_, _24642_);
  nand (_24647_, _24423_, _08027_);
  and (_24648_, _24647_, _24645_);
  or (_24649_, _24648_, _03113_);
  or (_24650_, _04735_, _10159_);
  and (_24651_, _24650_, _05741_);
  and (_24652_, _24651_, _24649_);
  and (_24653_, _09031_, _02592_);
  or (_24654_, _24653_, _02993_);
  or (_24655_, _24654_, _24652_);
  nor (_24656_, _09640_, _08841_);
  and (_24658_, _24433_, _09640_);
  or (_24659_, _24658_, _03549_);
  or (_24660_, _24659_, _24656_);
  and (_24661_, _24660_, _08795_);
  and (_24662_, _24661_, _24655_);
  nor (_24663_, _24424_, _08772_);
  nor (_24664_, _24663_, _10297_);
  or (_24665_, _24664_, _24662_);
  nand (_24666_, _09030_, _08772_);
  and (_24667_, _24666_, _09650_);
  and (_24669_, _24667_, _24665_);
  or (_24670_, _24669_, _24425_);
  and (_24671_, _24670_, _02855_);
  and (_24672_, _04735_, _02854_);
  or (_24673_, _24672_, _02575_);
  or (_24674_, _24673_, _24671_);
  nand (_24675_, _09030_, _02575_);
  and (_24676_, _24675_, _03134_);
  and (_24677_, _24676_, _24674_);
  and (_24678_, _09640_, _08842_);
  nor (_24680_, _24432_, _09640_);
  nor (_24681_, _24680_, _24678_);
  nor (_24682_, _24681_, _03134_);
  or (_24683_, _24682_, _24677_);
  nand (_24684_, _24683_, _09667_);
  or (_24685_, _24423_, _09667_);
  and (_24686_, _24685_, _24684_);
  or (_24687_, _24686_, _03133_);
  nand (_24688_, _09031_, _03133_);
  and (_24689_, _24688_, _09675_);
  and (_24691_, _24689_, _24687_);
  nor (_24692_, _24424_, _09675_);
  or (_24693_, _24692_, _02988_);
  or (_24694_, _24693_, _24691_);
  nand (_24695_, _02988_, _02889_);
  and (_24696_, _24695_, _05218_);
  and (_24697_, _24696_, _24694_);
  and (_24698_, _09030_, _02572_);
  or (_24699_, _24698_, _02778_);
  or (_24700_, _24699_, _24697_);
  or (_24702_, _24681_, _03142_);
  and (_24703_, _24702_, _09688_);
  and (_24704_, _24703_, _24700_);
  nor (_24705_, _24424_, _09688_);
  or (_24706_, _24705_, _02852_);
  or (_24707_, _24706_, _24704_);
  and (_24708_, _24707_, _24421_);
  nor (_24709_, _24708_, _21033_);
  nor (_24710_, _24423_, _09696_);
  nor (_24711_, _24710_, _02982_);
  not (_24713_, _24711_);
  nor (_24714_, _24713_, _24709_);
  nor (_24715_, _09699_, _02889_);
  nor (_24716_, _24715_, _24714_);
  or (_24717_, _24716_, _02568_);
  nand (_24718_, _09030_, _02568_);
  and (_24719_, _24718_, _24717_);
  nor (_24720_, _24719_, _09706_);
  and (_24721_, _24423_, _09706_);
  nor (_24722_, _24721_, _24720_);
  nand (_24724_, _24722_, _34446_);
  or (_24725_, _34446_, \oc8051_golden_model_1.PC [14]);
  and (_24726_, _24725_, _35583_);
  and (_35629_[14], _24726_, _24724_);
  and (_24727_, _34450_, \oc8051_golden_model_1.PSW [0]);
  nor (_24728_, _06856_, _06855_);
  nor (_24729_, _24728_, _06762_);
  and (_24730_, _24728_, _06762_);
  nor (_24731_, _24730_, _24729_);
  nor (_24732_, _06779_, _06778_);
  nor (_24734_, _24732_, _13770_);
  and (_24735_, _24732_, _13770_);
  nor (_24736_, _24735_, _24734_);
  and (_24737_, _24736_, _24731_);
  nor (_24738_, _24736_, _24731_);
  nor (_24739_, _24738_, _24737_);
  or (_24740_, _24739_, _05719_);
  nand (_24741_, _24739_, _05719_);
  and (_24742_, _24741_, _24740_);
  and (_24743_, _10316_, _19640_);
  nor (_24745_, _04108_, _02990_);
  and (_24746_, _24745_, _24743_);
  and (_24747_, _24746_, _05746_);
  or (_24748_, _24747_, _24742_);
  and (_24749_, _08809_, _08808_);
  or (_24750_, _24742_, _23355_);
  and (_24751_, _14105_, _07213_);
  nor (_24752_, _14105_, _07213_);
  nor (_24753_, _24752_, _24751_);
  and (_24754_, _13287_, _07217_);
  nor (_24756_, _24754_, _13885_);
  nor (_24757_, _24756_, _24753_);
  and (_24758_, _24756_, _24753_);
  nor (_24759_, _24758_, _24757_);
  and (_24760_, _07206_, _07202_);
  nor (_24761_, _07206_, _07202_);
  nor (_24762_, _24761_, _24760_);
  nor (_24763_, _24762_, _24759_);
  and (_24764_, _24762_, _24759_);
  nor (_24765_, _24764_, _24763_);
  nand (_24767_, _07199_, _07196_);
  or (_24768_, _07199_, _07196_);
  and (_24769_, _24768_, _24767_);
  nand (_24770_, _24769_, _24765_);
  or (_24771_, _24769_, _24765_);
  and (_24772_, _24771_, _24770_);
  or (_24773_, _24772_, _08821_);
  nor (_24774_, _14268_, _13967_);
  and (_24775_, _14268_, _13967_);
  nor (_24776_, _24775_, _24774_);
  nor (_24778_, _13659_, _13406_);
  and (_24779_, _13659_, _13406_);
  or (_24780_, _24779_, _24778_);
  nor (_24781_, _24780_, _24776_);
  and (_24782_, _24780_, _24776_);
  nor (_24783_, _24782_, _24781_);
  not (_24784_, _15168_);
  nor (_24785_, _14863_, _14563_);
  and (_24786_, _14863_, _14563_);
  nor (_24787_, _24786_, _24785_);
  nor (_24789_, _24787_, _24784_);
  and (_24790_, _24787_, _24784_);
  nor (_24791_, _24790_, _24789_);
  nor (_24792_, _24791_, _24783_);
  and (_24793_, _24791_, _24783_);
  or (_24794_, _24793_, _24792_);
  or (_24795_, _24794_, _07810_);
  nand (_24796_, _24794_, _07810_);
  and (_24797_, _24796_, _02974_);
  and (_24798_, _24797_, _24795_);
  and (_24800_, _03359_, _02794_);
  or (_24801_, _24742_, _02540_);
  or (_24802_, _24742_, _05325_);
  or (_24803_, _06118_, _05981_);
  nand (_24804_, _24803_, _10788_);
  or (_24805_, _24803_, _10788_);
  nand (_24806_, _24805_, _24804_);
  nor (_24807_, _06122_, _06073_);
  nand (_24808_, _24807_, _05798_);
  or (_24809_, _24807_, _05798_);
  nand (_24811_, _24809_, _24808_);
  nand (_24812_, _24811_, _24806_);
  or (_24813_, _24811_, _24806_);
  and (_24814_, _24813_, _24812_);
  nor (_24815_, _24814_, _05426_);
  and (_24816_, _24814_, _05426_);
  or (_24817_, _24816_, _24815_);
  and (_24818_, _24817_, _03343_);
  and (_24819_, _24742_, _02803_);
  and (_24820_, _02545_, \oc8051_golden_model_1.PSW [0]);
  or (_24822_, _24820_, _24819_);
  and (_24823_, _24822_, _07413_);
  nor (_24824_, _05330_, _05202_);
  nor (_24825_, _10606_, _05200_);
  and (_24826_, _10606_, _05200_);
  nor (_24827_, _24826_, _24825_);
  nor (_24828_, _24827_, _24824_);
  and (_24829_, _24827_, _24824_);
  nor (_24830_, _24829_, _24828_);
  not (_24831_, _24830_);
  and (_24833_, _05209_, _04839_);
  nor (_24834_, _05209_, _04839_);
  nor (_24835_, _24834_, _24833_);
  nand (_24836_, _24835_, _24831_);
  or (_24837_, _24835_, _24831_);
  and (_24838_, _24837_, _24836_);
  and (_24839_, _24838_, _14759_);
  or (_24840_, _24839_, _24823_);
  and (_24841_, _24840_, _07408_);
  or (_24842_, _24841_, _02934_);
  or (_24844_, _24842_, _24818_);
  and (_24845_, _07593_, _07572_);
  nor (_24846_, _24845_, _07957_);
  and (_24847_, _24846_, _07611_);
  nor (_24848_, _24846_, _07611_);
  nor (_24849_, _24848_, _24847_);
  nor (_24850_, _07651_, _07556_);
  and (_24851_, _07651_, _07556_);
  nor (_24852_, _24851_, _24850_);
  not (_24853_, _24852_);
  and (_24855_, _07952_, _07625_);
  and (_24856_, _07638_, _07951_);
  nor (_24857_, _24856_, _24855_);
  and (_24858_, _24857_, _24853_);
  nor (_24859_, _24857_, _24853_);
  nor (_24860_, _24859_, _24858_);
  nor (_24861_, _24860_, _24849_);
  and (_24862_, _24860_, _24849_);
  nor (_24863_, _24862_, _24861_);
  nor (_24864_, _24863_, _10031_);
  and (_24866_, _24863_, _10031_);
  or (_24867_, _24866_, _24864_);
  or (_24868_, _24867_, _07406_);
  and (_24869_, _24868_, _19664_);
  and (_24870_, _24869_, _24844_);
  and (_24871_, \oc8051_golden_model_1.XRAM_DATA_IN [0], \oc8051_golden_model_1.XRAM_DATA_IN [1]);
  nor (_24872_, \oc8051_golden_model_1.XRAM_DATA_IN [0], \oc8051_golden_model_1.XRAM_DATA_IN [1]);
  nor (_24873_, _24872_, _24871_);
  nor (_24874_, _24873_, _14770_);
  and (_24875_, _24873_, _14770_);
  or (_24877_, _24875_, _24874_);
  and (_24878_, \oc8051_golden_model_1.XRAM_DATA_IN [3], \oc8051_golden_model_1.XRAM_DATA_IN [2]);
  nor (_24879_, \oc8051_golden_model_1.XRAM_DATA_IN [3], \oc8051_golden_model_1.XRAM_DATA_IN [2]);
  or (_24880_, _24879_, _24878_);
  and (_24881_, _24880_, \oc8051_golden_model_1.XRAM_DATA_IN [4]);
  nor (_24882_, _24880_, \oc8051_golden_model_1.XRAM_DATA_IN [4]);
  nor (_24883_, _24882_, _24881_);
  and (_24884_, \oc8051_golden_model_1.XRAM_DATA_IN [7], \oc8051_golden_model_1.XRAM_DATA_IN [6]);
  nor (_24885_, \oc8051_golden_model_1.XRAM_DATA_IN [7], \oc8051_golden_model_1.XRAM_DATA_IN [6]);
  or (_24886_, _24885_, _24884_);
  and (_24888_, _24886_, _24883_);
  nor (_24889_, _24886_, _24883_);
  or (_24890_, _24889_, _24888_);
  and (_24891_, _24890_, _24877_);
  nor (_24892_, _24890_, _24877_);
  or (_24893_, _24892_, _24891_);
  and (_24894_, _24893_, _07432_);
  or (_24895_, _24894_, _09178_);
  or (_24896_, _24895_, _24870_);
  or (_24897_, _24742_, _02544_);
  and (_24899_, _24897_, _21080_);
  and (_24900_, _24899_, _24896_);
  nand (_24901_, _24893_, _07425_);
  nand (_24902_, _24901_, _05325_);
  or (_24903_, _24902_, _24900_);
  and (_24904_, _24903_, _24802_);
  or (_24905_, _24904_, _03806_);
  nor (_24906_, _24732_, \oc8051_golden_model_1.ACC [6]);
  and (_24907_, _24732_, \oc8051_golden_model_1.ACC [6]);
  nor (_24908_, _24907_, _24906_);
  nor (_24910_, _24908_, \oc8051_golden_model_1.ACC [7]);
  and (_24911_, _24908_, \oc8051_golden_model_1.ACC [7]);
  nor (_24912_, _24911_, _24910_);
  or (_24913_, _24912_, _24806_);
  nand (_24914_, _24912_, _24806_);
  and (_24915_, _24914_, _24913_);
  or (_24916_, _24915_, _05311_);
  and (_24917_, _24916_, _24905_);
  or (_24918_, _24917_, _02932_);
  not (_24919_, _13330_);
  nor (_24920_, _13564_, _24919_);
  and (_24921_, _13564_, _24919_);
  nor (_24922_, _24921_, _24920_);
  and (_24923_, _24922_, _13832_);
  nor (_24924_, _24922_, _13832_);
  nor (_24925_, _24924_, _24923_);
  and (_24926_, _24925_, _14755_);
  nor (_24927_, _24925_, _14755_);
  or (_24928_, _24927_, _24926_);
  not (_24929_, _14426_);
  and (_24932_, _24929_, _14149_);
  nor (_24933_, _24929_, _14149_);
  nor (_24934_, _24933_, _24932_);
  and (_24935_, _24934_, _24928_);
  nor (_24936_, _24934_, _24928_);
  nor (_24937_, _24936_, _24935_);
  and (_24938_, _24937_, _15039_);
  nor (_24939_, _24937_, _15039_);
  or (_24940_, _24939_, _24938_);
  and (_24941_, _24940_, _07404_);
  nor (_24943_, _24940_, _07404_);
  or (_24944_, _24943_, _24941_);
  or (_24945_, _24944_, _06162_);
  and (_24946_, _24945_, _09879_);
  and (_24947_, _24946_, _24918_);
  and (_24948_, _13568_, _06908_);
  or (_24949_, _24948_, _13839_);
  and (_24950_, _24949_, _14448_);
  nor (_24951_, _24949_, _14448_);
  nor (_24952_, _24951_, _24950_);
  nor (_24954_, _14156_, _13771_);
  and (_24955_, _14156_, _13771_);
  nor (_24956_, _24955_, _24954_);
  not (_24957_, _24956_);
  and (_24958_, _24957_, _24952_);
  nor (_24959_, _24957_, _24952_);
  nor (_24960_, _24959_, _24958_);
  and (_24961_, _24960_, _14778_);
  nor (_24962_, _24960_, _14778_);
  nor (_24963_, _24962_, _24961_);
  nor (_24964_, _15062_, _07459_);
  and (_24965_, _15062_, _07459_);
  nor (_24966_, _24965_, _24964_);
  not (_24967_, _24966_);
  nand (_24968_, _24967_, _24963_);
  or (_24969_, _24967_, _24963_);
  and (_24970_, _24969_, _07402_);
  and (_24971_, _24970_, _24968_);
  or (_24972_, _24971_, _09017_);
  or (_24973_, _24972_, _24947_);
  not (_24976_, _09017_);
  or (_24977_, _24742_, _24976_);
  and (_24978_, _24977_, _03186_);
  and (_24979_, _24978_, _24973_);
  and (_24980_, _13577_, _13308_);
  nor (_24981_, _13577_, _13308_);
  or (_24982_, _24981_, _24980_);
  nor (_24983_, _14160_, _13846_);
  and (_24984_, _14160_, _13846_);
  nor (_24985_, _24984_, _24983_);
  not (_24987_, _24985_);
  and (_24988_, _24987_, _24982_);
  nor (_24989_, _24987_, _24982_);
  nor (_24990_, _24989_, _24988_);
  not (_24991_, _15068_);
  nor (_24992_, _14782_, _14454_);
  and (_24993_, _14782_, _14454_);
  nor (_24994_, _24993_, _24992_);
  nor (_24995_, _24994_, _24991_);
  and (_24996_, _24994_, _24991_);
  nor (_24997_, _24996_, _24995_);
  and (_24998_, _24997_, _24990_);
  nor (_24999_, _24997_, _24990_);
  nor (_25000_, _24999_, _24998_);
  and (_25001_, _25000_, _07465_);
  nor (_25002_, _25000_, _07465_);
  or (_25003_, _25002_, _25001_);
  and (_25004_, _25003_, _02799_);
  or (_25005_, _25004_, _04239_);
  or (_25006_, _25005_, _24979_);
  and (_25009_, _25006_, _24801_);
  or (_25010_, _25009_, _02930_);
  and (_25011_, _13534_, _13299_);
  nor (_25012_, _13534_, _13299_);
  nor (_25013_, _25012_, _25011_);
  not (_25014_, _14121_);
  and (_25015_, _25014_, _13809_);
  nor (_25016_, _25014_, _13809_);
  nor (_25017_, _25016_, _25015_);
  nor (_25018_, _25017_, _25013_);
  and (_25020_, _25017_, _25013_);
  or (_25021_, _25020_, _25018_);
  nor (_25022_, _14718_, _14418_);
  and (_25023_, _14718_, _14418_);
  nor (_25024_, _25023_, _25022_);
  and (_25025_, _25024_, _15018_);
  nor (_25026_, _25024_, _15018_);
  nor (_25027_, _25026_, _25025_);
  nor (_25028_, _25027_, _25021_);
  and (_25029_, _25027_, _25021_);
  nor (_25031_, _25029_, _25028_);
  nand (_25032_, _25031_, _07327_);
  or (_25033_, _25031_, _07327_);
  and (_25034_, _25033_, _25032_);
  or (_25035_, _25034_, _03693_);
  and (_25036_, _25035_, _07475_);
  and (_25037_, _25036_, _25010_);
  and (_25038_, _10346_, _02794_);
  and (_25039_, _24838_, _07476_);
  or (_25040_, _25039_, _25038_);
  or (_25042_, _25040_, _25037_);
  not (_25043_, _25038_);
  or (_25044_, _24817_, _25043_);
  and (_25045_, _25044_, _25042_);
  or (_25046_, _25045_, _24800_);
  not (_25047_, _24800_);
  or (_25048_, _24817_, _25047_);
  and (_25049_, _25048_, _02943_);
  and (_25050_, _25049_, _25046_);
  and (_25051_, _24867_, _02928_);
  or (_25052_, _25051_, _09206_);
  or (_25053_, _25052_, _25050_);
  or (_25054_, _24742_, _09212_);
  and (_25055_, _25054_, _02927_);
  and (_25056_, _25055_, _25053_);
  and (_25057_, _13596_, _13293_);
  nor (_25058_, _13596_, _13293_);
  or (_25059_, _25058_, _25057_);
  not (_25060_, _14178_);
  and (_25061_, _25060_, _13864_);
  nor (_25064_, _25060_, _13864_);
  nor (_25065_, _25064_, _25061_);
  nor (_25066_, _25065_, _25059_);
  and (_25067_, _25065_, _25059_);
  or (_25068_, _25067_, _25066_);
  nor (_25069_, _14800_, _14472_);
  and (_25070_, _14800_, _14472_);
  nor (_25071_, _25070_, _25069_);
  nor (_25072_, _25071_, _15087_);
  and (_25073_, _25071_, _15087_);
  nor (_25075_, _25073_, _25072_);
  nor (_25076_, _25075_, _25068_);
  and (_25077_, _25075_, _25068_);
  nor (_25078_, _25077_, _25076_);
  nand (_25079_, _25078_, _07494_);
  or (_25080_, _25078_, _07494_);
  and (_25081_, _25080_, _25079_);
  nand (_25082_, _25081_, _02796_);
  and (_25083_, _10299_, _09927_);
  nor (_25084_, _08827_, _09209_);
  and (_25086_, _25084_, _25083_);
  nand (_25087_, _25086_, _25082_);
  or (_25088_, _25087_, _25056_);
  or (_25089_, _25086_, _24742_);
  and (_25090_, _25089_, _06189_);
  and (_25091_, _25090_, _25088_);
  not (_25092_, _14751_);
  nor (_25093_, _13869_, _13601_);
  and (_25094_, _13869_, _13601_);
  nor (_25095_, _25094_, _25093_);
  nor (_25097_, _25095_, _25092_);
  and (_25098_, _25095_, _25092_);
  nor (_25099_, _25098_, _25097_);
  nor (_25100_, _14126_, _24919_);
  and (_25101_, _14126_, _24919_);
  nor (_25102_, _25101_, _25100_);
  nor (_25103_, _25102_, _14477_);
  and (_25104_, _25102_, _14477_);
  or (_25105_, _25104_, _25103_);
  nor (_25106_, _15092_, _07499_);
  and (_25108_, _15092_, _07499_);
  nor (_25109_, _25108_, _25106_);
  nor (_25110_, _25109_, _25105_);
  and (_25111_, _25109_, _25105_);
  or (_25112_, _25111_, _25110_);
  nand (_25113_, _25112_, _25099_);
  or (_25114_, _25112_, _25099_);
  and (_25115_, _25114_, _02790_);
  nand (_25116_, _25115_, _25113_);
  not (_25117_, _09271_);
  and (_25119_, _22616_, _25117_);
  nand (_25120_, _25119_, _25116_);
  or (_25121_, _25120_, _25091_);
  or (_25122_, _25119_, _24742_);
  and (_25123_, _25122_, _06201_);
  and (_25124_, _25123_, _25121_);
  and (_25125_, _10342_, _08210_);
  nor (_25126_, _13607_, _13355_);
  and (_25127_, _13607_, _13355_);
  or (_25128_, _25127_, _25126_);
  nor (_25130_, _25128_, _13874_);
  and (_25131_, _25128_, _13874_);
  nor (_25132_, _25131_, _25130_);
  nor (_25133_, _25132_, _14185_);
  and (_25134_, _25132_, _14185_);
  or (_25135_, _25134_, _25133_);
  nor (_25136_, _25135_, _14482_);
  and (_25137_, _25135_, _14482_);
  or (_25138_, _25137_, _25136_);
  nor (_25139_, _25138_, _14807_);
  and (_25141_, _25138_, _14807_);
  or (_25142_, _25141_, _25139_);
  nor (_25143_, _25142_, _15098_);
  and (_25144_, _25142_, _15098_);
  or (_25145_, _25144_, _25143_);
  or (_25146_, _25145_, _07504_);
  nand (_25147_, _25145_, _07504_);
  and (_25148_, _25147_, _06195_);
  nand (_25149_, _25148_, _25146_);
  nand (_25150_, _25149_, _25125_);
  or (_25152_, _25150_, _25124_);
  or (_25153_, _24742_, _25125_);
  and (_25154_, _25153_, _09759_);
  and (_25155_, _25154_, _25152_);
  and (_25156_, _24742_, _02901_);
  or (_25157_, _25156_, _07399_);
  or (_25158_, _25157_, _25155_);
  not (_25159_, _07399_);
  and (_25160_, _13616_, _13359_);
  nor (_25161_, _25160_, _07525_);
  and (_25163_, _25161_, _13892_);
  nor (_25164_, _25161_, _13892_);
  or (_25165_, _25164_, _25163_);
  nor (_25166_, _25165_, _14199_);
  and (_25167_, _25165_, _14199_);
  nor (_25168_, _25167_, _25166_);
  or (_25169_, _25168_, _14499_);
  nand (_25170_, _25168_, _14499_);
  and (_25171_, _25170_, _25169_);
  nor (_25172_, _25171_, _14823_);
  and (_25174_, _25171_, _14823_);
  or (_25175_, _25174_, _25172_);
  nor (_25176_, _25175_, _15114_);
  and (_25177_, _25175_, _15114_);
  or (_25178_, _25177_, _25176_);
  nor (_25179_, _25178_, _07534_);
  and (_25180_, _25178_, _07534_);
  or (_25181_, _25180_, _25179_);
  or (_25182_, _25181_, _25159_);
  and (_25183_, _25182_, _25158_);
  or (_25184_, _25183_, _07398_);
  not (_25185_, _07398_);
  or (_25186_, _25181_, _25185_);
  and (_25187_, _25186_, _07330_);
  and (_25188_, _25187_, _25184_);
  or (_25189_, _13624_, _13367_);
  nand (_25190_, _13624_, _13367_);
  and (_25191_, _25190_, _25189_);
  nor (_25192_, _25191_, _13910_);
  and (_25193_, _25191_, _13910_);
  nor (_25196_, _25193_, _25192_);
  and (_25197_, _25196_, _14214_);
  nor (_25198_, _25196_, _14214_);
  or (_25199_, _25198_, _25197_);
  and (_25200_, _14746_, _14516_);
  nor (_25201_, _14746_, _14516_);
  or (_25202_, _25201_, _25200_);
  and (_25203_, _25202_, _25199_);
  nor (_25204_, _25202_, _25199_);
  nor (_25205_, _25204_, _25203_);
  nor (_25207_, _25205_, _15035_);
  and (_25208_, _25205_, _15035_);
  or (_25209_, _25208_, _25207_);
  and (_25210_, _25209_, _07396_);
  nor (_25211_, _25209_, _07396_);
  or (_25212_, _25211_, _25210_);
  and (_25213_, _25212_, _07329_);
  or (_25214_, _25213_, _02898_);
  or (_25215_, _25214_, _25188_);
  not (_25216_, _07696_);
  not (_25218_, _14223_);
  nand (_25219_, _13540_, _13372_);
  or (_25220_, _13540_, _13372_);
  and (_25221_, _25220_, _25219_);
  nor (_25222_, _25221_, _13920_);
  and (_25223_, _25221_, _13920_);
  nor (_25224_, _25223_, _25222_);
  and (_25225_, _25224_, _25218_);
  nor (_25226_, _25224_, _25218_);
  nor (_25227_, _25226_, _25225_);
  nor (_25229_, _25227_, _14421_);
  and (_25230_, _25227_, _14421_);
  or (_25231_, _25230_, _25229_);
  nor (_25232_, _25231_, _14830_);
  and (_25233_, _25231_, _14830_);
  or (_25234_, _25233_, _25232_);
  nor (_25235_, _25234_, _15021_);
  and (_25236_, _25234_, _15021_);
  or (_25237_, _25236_, _25235_);
  nor (_25238_, _25237_, _25216_);
  and (_25240_, _25237_, _25216_);
  or (_25241_, _25240_, _25238_);
  or (_25242_, _25241_, _02899_);
  and (_25243_, _25242_, _07541_);
  and (_25244_, _25243_, _25215_);
  or (_25245_, _07769_, _07759_);
  and (_25246_, _25245_, _07770_);
  nand (_25247_, _25246_, _13936_);
  or (_25248_, _25246_, _13936_);
  and (_25249_, _25248_, _25247_);
  nor (_25251_, _25249_, _14237_);
  and (_25252_, _25249_, _14237_);
  or (_25253_, _25252_, _25251_);
  and (_25254_, _14732_, _14532_);
  nor (_25255_, _14732_, _14532_);
  or (_25256_, _25255_, _25254_);
  and (_25257_, _25256_, _25253_);
  nor (_25258_, _25256_, _25253_);
  nor (_25259_, _25258_, _25257_);
  and (_25260_, _25259_, _15132_);
  nor (_25262_, _25259_, _15132_);
  nor (_25263_, _25262_, _25260_);
  nor (_25264_, _25263_, _07779_);
  and (_25265_, _25263_, _07779_);
  or (_25266_, _25265_, _25264_);
  and (_25267_, _25266_, _07540_);
  or (_25268_, _25267_, _07700_);
  or (_25269_, _25268_, _25244_);
  nor (_25270_, _04587_, _02890_);
  nor (_25271_, _04622_, _04598_);
  nor (_25273_, _04614_, _04603_);
  not (_25274_, _25273_);
  nor (_25275_, _04650_, _04591_);
  and (_25276_, _25275_, _25274_);
  nor (_25277_, _25275_, _25274_);
  nor (_25278_, _25277_, _25276_);
  nor (_25279_, _25278_, _25271_);
  and (_25280_, _25278_, _25271_);
  nor (_25281_, _25280_, _25279_);
  nor (_25282_, _25281_, _25270_);
  and (_25284_, _25281_, _25270_);
  or (_25285_, _25284_, _25282_);
  or (_25286_, _25285_, _02499_);
  and (_25287_, _25286_, _02966_);
  and (_25288_, _25287_, _25269_);
  not (_25289_, _07788_);
  nor (_25290_, _13636_, _13383_);
  and (_25291_, _13636_, _13383_);
  nor (_25292_, _25291_, _25290_);
  not (_25293_, _25292_);
  nor (_25295_, _14840_, _14540_);
  and (_25296_, _14840_, _14540_);
  nor (_25297_, _25296_, _25295_);
  and (_25298_, _25297_, _25293_);
  nor (_25299_, _25297_, _25293_);
  nor (_25300_, _25299_, _25298_);
  not (_25301_, _15141_);
  not (_25302_, _14245_);
  and (_25303_, _25302_, _13944_);
  nor (_25304_, _25302_, _13944_);
  nor (_25306_, _25304_, _25303_);
  nor (_25307_, _25306_, _25301_);
  and (_25308_, _25306_, _25301_);
  nor (_25309_, _25308_, _25307_);
  and (_25310_, _25309_, _25300_);
  nor (_25311_, _25309_, _25300_);
  nor (_25312_, _25311_, _25310_);
  nand (_25313_, _25312_, _25289_);
  or (_25314_, _25312_, _25289_);
  and (_25315_, _25314_, _02785_);
  and (_25317_, _25315_, _25313_);
  or (_25318_, _25317_, _22645_);
  or (_25319_, _25318_, _25288_);
  or (_25320_, _24742_, _22644_);
  and (_25321_, _25320_, _03856_);
  and (_25322_, _25321_, _25319_);
  and (_25323_, _25034_, _20307_);
  or (_25324_, _25323_, _25322_);
  and (_25325_, _25324_, _03859_);
  and (_25326_, _25034_, _03858_);
  or (_25328_, _25326_, _03850_);
  or (_25329_, _25328_, _25325_);
  and (_25330_, _13643_, _13390_);
  nor (_25331_, _13643_, _13390_);
  nor (_25332_, _25331_, _25330_);
  and (_25333_, _25332_, _13951_);
  nor (_25334_, _25332_, _13951_);
  or (_25335_, _25334_, _25333_);
  and (_25336_, _25335_, _14252_);
  nor (_25337_, _25335_, _14252_);
  or (_25339_, _25337_, _25336_);
  not (_25340_, _14847_);
  and (_25341_, _25340_, _14547_);
  nor (_25342_, _25340_, _14547_);
  nor (_25343_, _25342_, _25341_);
  nand (_25344_, _25343_, _15149_);
  or (_25345_, _25343_, _15149_);
  and (_25346_, _25345_, _25344_);
  or (_25347_, _25346_, _25339_);
  nand (_25348_, _25346_, _25339_);
  and (_25350_, _25348_, _25347_);
  and (_25351_, _07322_, _02970_);
  and (_25352_, _25351_, _25350_);
  nand (_25353_, _25350_, _03850_);
  and (_25354_, _25353_, _07324_);
  or (_25355_, _25354_, _25352_);
  and (_25356_, _25355_, _25329_);
  and (_25357_, _13648_, _13395_);
  nor (_25358_, _13648_, _13395_);
  nor (_25359_, _25358_, _25357_);
  and (_25360_, _25359_, _13956_);
  nor (_25361_, _25359_, _13956_);
  or (_25362_, _25361_, _25360_);
  nand (_25363_, _25362_, _14257_);
  or (_25364_, _25362_, _14257_);
  and (_25365_, _25364_, _25363_);
  nor (_25366_, _15154_, _14852_);
  and (_25367_, _15154_, _14852_);
  nor (_25368_, _25367_, _25366_);
  not (_25369_, _07796_);
  nor (_25372_, _14552_, _25369_);
  and (_25373_, _14552_, _25369_);
  nor (_25374_, _25373_, _25372_);
  nor (_25375_, _25374_, _25368_);
  and (_25376_, _25374_, _25368_);
  nor (_25377_, _25376_, _25375_);
  nand (_25378_, _25377_, _25365_);
  or (_25379_, _25377_, _25365_);
  and (_25380_, _25379_, _02524_);
  and (_25381_, _25380_, _25378_);
  or (_25383_, _25381_, _06731_);
  or (_25384_, _25383_, _25356_);
  nor (_25385_, _06928_, _06873_);
  and (_25386_, _06928_, _06873_);
  nor (_25387_, _25386_, _25385_);
  nor (_25388_, _25387_, _06823_);
  and (_25389_, _25387_, _06823_);
  nor (_25390_, _25389_, _25388_);
  and (_25391_, _25390_, _15160_);
  nor (_25392_, _25390_, _15160_);
  nor (_25394_, _25392_, _25391_);
  nor (_25395_, _06793_, _07800_);
  and (_25396_, _06793_, _07800_);
  nor (_25397_, _25396_, _25395_);
  and (_25398_, _25397_, _25394_);
  nor (_25399_, _25397_, _25394_);
  or (_25400_, _25399_, _25398_);
  nor (_25401_, _25400_, _06992_);
  and (_25402_, _25400_, _06992_);
  nor (_25403_, _25402_, _25401_);
  and (_25405_, _25403_, _07086_);
  nor (_25406_, _25403_, _07086_);
  or (_25407_, _25406_, _06737_);
  or (_25408_, _25407_, _25405_);
  and (_25409_, _25408_, _02552_);
  and (_25410_, _25409_, _25384_);
  nand (_25411_, _25285_, _02476_);
  nor (_25412_, _09318_, _04094_);
  and (_25413_, _25412_, _09315_);
  nand (_25414_, _25413_, _25411_);
  or (_25416_, _25414_, _25410_);
  or (_25417_, _25413_, _24742_);
  nand (_25418_, _25417_, _25416_);
  nor (_25419_, _04100_, _03870_);
  and (_25420_, _25419_, _04107_);
  and (_25421_, _25420_, _05263_);
  nand (_25422_, _25421_, _25418_);
  or (_25423_, _25421_, _24742_);
  and (_25424_, _25423_, _05261_);
  and (_25425_, _25424_, _25422_);
  or (_25427_, _25425_, _24798_);
  and (_25428_, _25427_, _07808_);
  nand (_25429_, _25285_, _07807_);
  nand (_25430_, _25429_, _10332_);
  or (_25431_, _25430_, _25428_);
  or (_25432_, _24742_, _10332_);
  and (_25433_, _25432_, _09376_);
  and (_25434_, _25433_, _25431_);
  nand (_25435_, _24742_, _09375_);
  nand (_25436_, _25435_, _08821_);
  or (_25438_, _25436_, _25434_);
  and (_25439_, _25438_, _24773_);
  or (_25440_, _25439_, _07832_);
  and (_25441_, _13423_, _07166_);
  nor (_25442_, _25441_, _13903_);
  and (_25443_, _14203_, _07162_);
  nor (_25444_, _14203_, _07162_);
  nor (_25445_, _25444_, _25443_);
  nor (_25446_, _25445_, _25442_);
  and (_25447_, _25445_, _25442_);
  nor (_25449_, _25447_, _25446_);
  and (_25450_, _07157_, _07153_);
  nor (_25451_, _07157_, _07153_);
  nor (_25452_, _25451_, _25450_);
  nor (_25453_, _25452_, _25449_);
  and (_25454_, _25452_, _25449_);
  or (_25455_, _25454_, _25453_);
  and (_25456_, _25455_, _07150_);
  nor (_25457_, _25455_, _07150_);
  nor (_25458_, _25457_, _25456_);
  nor (_25460_, _25458_, _07147_);
  and (_25461_, _25458_, _07147_);
  or (_25462_, _25461_, _25460_);
  or (_25463_, _25462_, _07833_);
  and (_25464_, _25463_, _03106_);
  and (_25465_, _25464_, _25440_);
  nor (_25466_, _10610_, _10546_);
  and (_25467_, _10610_, _10546_);
  nor (_25468_, _25467_, _25466_);
  not (_25469_, _25468_);
  nor (_25471_, _11134_, _10942_);
  and (_25472_, _11134_, _10942_);
  nor (_25473_, _25472_, _25471_);
  and (_25474_, _25473_, _25469_);
  nor (_25475_, _25473_, _25469_);
  nor (_25476_, _25475_, _25474_);
  or (_25477_, _25476_, _11333_);
  nand (_25478_, _25476_, _11333_);
  and (_25479_, _25478_, _25477_);
  nor (_25480_, _25479_, _11531_);
  and (_25482_, _25479_, _11531_);
  or (_25483_, _25482_, _25480_);
  nor (_25484_, _25483_, _11601_);
  and (_25485_, _25483_, _11601_);
  nor (_25486_, _25485_, _25484_);
  not (_25487_, _25486_);
  nor (_25488_, _25487_, _05722_);
  and (_25489_, _25487_, _05722_);
  or (_25490_, _25489_, _25488_);
  and (_25491_, _25490_, _03105_);
  or (_25493_, _25491_, _07319_);
  or (_25494_, _25493_, _25465_);
  and (_25495_, _08105_, _07845_);
  nor (_25496_, _25495_, _08836_);
  nor (_25497_, _14964_, _08110_);
  and (_25498_, _14964_, _08110_);
  or (_25499_, _25498_, _25497_);
  not (_25500_, _25499_);
  and (_25501_, _08832_, _08115_);
  nor (_25502_, _25501_, _08833_);
  not (_25504_, _25502_);
  and (_25505_, _08830_, _07762_);
  nor (_25506_, _25505_, _08831_);
  and (_25507_, _25506_, _25504_);
  nor (_25508_, _25506_, _25504_);
  nor (_25509_, _25508_, _25507_);
  nor (_25510_, _25509_, _25500_);
  and (_25511_, _25509_, _25500_);
  nor (_25512_, _25511_, _25510_);
  not (_25513_, _25512_);
  nor (_25515_, _25513_, _25496_);
  and (_25516_, _25513_, _25496_);
  or (_25517_, _25516_, _25515_);
  or (_25518_, _25517_, _07846_);
  and (_25519_, _25518_, _07092_);
  and (_25520_, _25519_, _25494_);
  not (_25521_, _15014_);
  nor (_25522_, _13530_, _13295_);
  and (_25523_, _13530_, _13295_);
  nor (_25524_, _25523_, _25522_);
  not (_25526_, _14115_);
  and (_25527_, _25526_, _13806_);
  nor (_25528_, _25526_, _13806_);
  nor (_25529_, _25528_, _25527_);
  nor (_25530_, _25529_, _25524_);
  and (_25531_, _25529_, _25524_);
  or (_25532_, _25531_, _25530_);
  not (_25533_, _14713_);
  and (_25534_, _25533_, _14415_);
  nor (_25535_, _25533_, _14415_);
  nor (_25537_, _25535_, _25534_);
  and (_25538_, _25537_, _25532_);
  nor (_25539_, _25537_, _25532_);
  nor (_25540_, _25539_, _25538_);
  nor (_25541_, _25540_, _25521_);
  and (_25542_, _25540_, _25521_);
  or (_25543_, _25542_, _25541_);
  and (_25544_, _25543_, _07851_);
  nor (_25545_, _25543_, _07851_);
  or (_25546_, _25545_, _25544_);
  and (_25548_, _25546_, _02977_);
  or (_25549_, _25548_, _25520_);
  and (_25550_, _25549_, _07104_);
  nand (_25551_, _24742_, _03107_);
  or (_25552_, _25551_, _04654_);
  nand (_25553_, _25552_, _23355_);
  or (_25554_, _25553_, _25550_);
  and (_25555_, _25554_, _24750_);
  or (_25556_, _25555_, _07860_);
  not (_25557_, _03225_);
  or (_25558_, _07218_, _07215_);
  nand (_25559_, _07218_, _07215_);
  and (_25560_, _25559_, _25558_);
  nor (_25561_, _07211_, _07209_);
  and (_25562_, _07211_, _07209_);
  nor (_25563_, _25562_, _25561_);
  not (_25564_, _25563_);
  and (_25565_, _25564_, _25560_);
  nor (_25566_, _25564_, _25560_);
  nor (_25567_, _25566_, _25565_);
  nor (_25570_, _07204_, _07200_);
  and (_25571_, _07204_, _07200_);
  nor (_25572_, _25571_, _25570_);
  and (_25573_, _07197_, _07195_);
  nor (_25574_, _25573_, _10116_);
  nor (_25575_, _25574_, _25572_);
  and (_25576_, _25574_, _25572_);
  nor (_25577_, _25576_, _25575_);
  or (_25578_, _25577_, _25567_);
  nand (_25579_, _25577_, _25567_);
  and (_25581_, _25579_, _25578_);
  and (_25582_, _25581_, _25557_);
  or (_25583_, _25582_, _07865_);
  and (_25584_, _25583_, _07867_);
  and (_25585_, _25584_, _25556_);
  or (_25586_, _07866_, _03225_);
  and (_25587_, _25581_, _25586_);
  or (_25588_, _25587_, _03499_);
  or (_25589_, _25588_, _25585_);
  not (_25590_, _07146_);
  not (_25592_, _07160_);
  or (_25593_, _07167_, _07164_);
  nand (_25594_, _07167_, _07164_);
  and (_25595_, _25594_, _25593_);
  nand (_25596_, _25595_, _25592_);
  or (_25597_, _25595_, _25592_);
  and (_25598_, _25597_, _25596_);
  nor (_25599_, _25598_, _07158_);
  and (_25600_, _25598_, _07158_);
  or (_25601_, _25600_, _25599_);
  not (_25603_, _07151_);
  nor (_25604_, _07155_, _07148_);
  and (_25605_, _07155_, _07148_);
  nor (_25606_, _25605_, _25604_);
  nor (_25607_, _25606_, _25603_);
  and (_25608_, _25606_, _25603_);
  nor (_25609_, _25608_, _25607_);
  not (_25610_, _25609_);
  nor (_25611_, _25610_, _25601_);
  and (_25612_, _25610_, _25601_);
  nor (_25614_, _25612_, _25611_);
  and (_25615_, _25614_, _25590_);
  nor (_25616_, _25614_, _25590_);
  or (_25617_, _25616_, _07876_);
  or (_25618_, _25617_, _25615_);
  and (_25619_, _25618_, _07881_);
  and (_25620_, _25619_, _25589_);
  not (_25621_, _08108_);
  or (_25622_, _08117_, _07761_);
  nand (_25623_, _08117_, _07761_);
  and (_25625_, _25623_, _25622_);
  not (_25626_, _08111_);
  and (_25627_, _25626_, _08113_);
  nor (_25628_, _25626_, _08113_);
  nor (_25629_, _25628_, _25627_);
  not (_25630_, _25629_);
  and (_25631_, _25630_, _25625_);
  nor (_25632_, _25630_, _25625_);
  nor (_25633_, _25632_, _25631_);
  nand (_25634_, _25633_, _25621_);
  or (_25636_, _25633_, _25621_);
  and (_25637_, _25636_, _25634_);
  or (_25638_, _25637_, _08106_);
  nand (_25639_, _25637_, _08106_);
  and (_25640_, _25639_, _25638_);
  nor (_25641_, _25640_, _08103_);
  and (_25642_, _25640_, _08103_);
  or (_25643_, _25642_, _25641_);
  nor (_25644_, _25643_, _09717_);
  and (_25645_, _25643_, _09717_);
  or (_25647_, _25645_, _25644_);
  and (_25648_, _25647_, _07880_);
  not (_25649_, _05720_);
  nor (_25650_, _10608_, _10545_);
  and (_25651_, _10608_, _10545_);
  nor (_25652_, _25651_, _25650_);
  not (_25653_, _25652_);
  not (_25654_, _11132_);
  and (_25655_, _25654_, _10940_);
  nor (_25656_, _25654_, _10940_);
  nor (_25658_, _25656_, _25655_);
  nor (_25659_, _25658_, _25653_);
  and (_25660_, _25658_, _25653_);
  nor (_25661_, _25660_, _25659_);
  not (_25662_, _11599_);
  nor (_25663_, _11529_, _11331_);
  and (_25664_, _11529_, _11331_);
  nor (_25665_, _25664_, _25663_);
  nor (_25666_, _25665_, _25662_);
  and (_25667_, _25665_, _25662_);
  nor (_25669_, _25667_, _25666_);
  not (_25670_, _25669_);
  nor (_25671_, _25670_, _25661_);
  and (_25672_, _25670_, _25661_);
  nor (_25673_, _25672_, _25671_);
  nor (_25674_, _25673_, _25649_);
  and (_25675_, _25673_, _25649_);
  or (_25676_, _25675_, _25674_);
  and (_25677_, _25676_, _03092_);
  or (_25678_, _25677_, _25648_);
  or (_25680_, _25678_, _25620_);
  and (_25681_, _25680_, _03881_);
  nor (_25682_, _14011_, _13452_);
  and (_25683_, _14011_, _13452_);
  nor (_25684_, _25683_, _25682_);
  nor (_25685_, _15218_, _14604_);
  and (_25686_, _15218_, _14604_);
  nor (_25687_, _25686_, _25685_);
  and (_25688_, _25687_, _25684_);
  nor (_25689_, _25687_, _25684_);
  nor (_25691_, _25689_, _25688_);
  not (_25692_, _14311_);
  and (_25693_, _25692_, _13699_);
  nor (_25694_, _25692_, _13699_);
  nor (_25695_, _25694_, _25693_);
  nor (_25696_, _14903_, _07890_);
  and (_25697_, _14903_, _07890_);
  nor (_25698_, _25697_, _25696_);
  and (_25699_, _25698_, _25695_);
  nor (_25700_, _25698_, _25695_);
  nor (_25702_, _25700_, _25699_);
  nand (_25703_, _25702_, _25691_);
  or (_25704_, _25702_, _25691_);
  and (_25705_, _25704_, _02991_);
  and (_25706_, _25705_, _25703_);
  or (_25707_, _25706_, _25681_);
  and (_25708_, _25707_, _24749_);
  nor (_25709_, _14410_, _14310_);
  not (_25710_, _24749_);
  nand (_25711_, _24742_, _25710_);
  nand (_25713_, _25711_, _25709_);
  or (_25714_, _25713_, _25708_);
  nor (_25715_, _13286_, _07216_);
  and (_25716_, _13286_, _07216_);
  nor (_25717_, _25716_, _25715_);
  not (_25718_, _25717_);
  nor (_25719_, _07212_, _14319_);
  and (_25720_, _07212_, _14319_);
  nor (_25721_, _25720_, _25719_);
  nor (_25722_, _25721_, _25718_);
  and (_25724_, _25721_, _25718_);
  nor (_25725_, _25724_, _25722_);
  not (_25726_, _07201_);
  nor (_25727_, _07205_, _07198_);
  and (_25728_, _07205_, _07198_);
  nor (_25729_, _25728_, _25727_);
  nor (_25730_, _25729_, _25726_);
  and (_25731_, _25729_, _25726_);
  nor (_25732_, _25731_, _25730_);
  not (_25733_, _25732_);
  nor (_25735_, _25733_, _25725_);
  and (_25736_, _25733_, _25725_);
  nor (_25737_, _25736_, _25735_);
  nand (_25738_, _25737_, _07194_);
  or (_25739_, _25737_, _07194_);
  and (_25740_, _25739_, _25738_);
  or (_25741_, _25740_, _25709_);
  and (_25742_, _25741_, _03525_);
  and (_25743_, _25742_, _25714_);
  and (_25744_, _25740_, _03524_);
  or (_25746_, _25744_, _07315_);
  or (_25747_, _25746_, _25743_);
  nor (_25748_, _13422_, _07165_);
  and (_25749_, _13422_, _07165_);
  nor (_25750_, _25749_, _25748_);
  and (_25751_, _25750_, _07161_);
  nor (_25752_, _25750_, _07161_);
  or (_25753_, _25752_, _25751_);
  and (_25754_, _25753_, _07159_);
  nor (_25755_, _25753_, _07159_);
  or (_25757_, _25755_, _25754_);
  not (_25758_, _07152_);
  nor (_25759_, _07156_, _07149_);
  and (_25760_, _07156_, _07149_);
  nor (_25761_, _25760_, _25759_);
  nor (_25762_, _25761_, _25758_);
  and (_25763_, _25761_, _25758_);
  nor (_25764_, _25763_, _25762_);
  not (_25765_, _25764_);
  nor (_25766_, _25765_, _25757_);
  and (_25768_, _25765_, _25757_);
  nor (_25769_, _25768_, _25766_);
  nand (_25770_, _25769_, _07145_);
  or (_25771_, _25769_, _07145_);
  and (_25772_, _25771_, _25770_);
  or (_25773_, _25772_, _08804_);
  and (_25774_, _25773_, _03098_);
  and (_25775_, _25774_, _25747_);
  nor (_25776_, _10609_, _10423_);
  and (_25777_, _10609_, _10423_);
  nor (_25779_, _25777_, _25776_);
  and (_25780_, _25779_, _10941_);
  nor (_25781_, _25779_, _10941_);
  or (_25782_, _25781_, _25780_);
  nand (_25783_, _25782_, _11133_);
  or (_25784_, _25782_, _11133_);
  and (_25785_, _25784_, _25783_);
  nor (_25786_, _11530_, _11332_);
  and (_25787_, _11530_, _11332_);
  nor (_25788_, _25787_, _25786_);
  nor (_25790_, _25788_, _11600_);
  and (_25791_, _25788_, _11600_);
  nor (_25792_, _25791_, _25790_);
  and (_25793_, _25792_, _25785_);
  nor (_25794_, _25792_, _25785_);
  nor (_25795_, _25794_, _25793_);
  and (_25796_, _25795_, _05721_);
  nor (_25797_, _25795_, _05721_);
  or (_25798_, _25797_, _25796_);
  and (_25799_, _25798_, _03097_);
  or (_25801_, _25799_, _07899_);
  or (_25802_, _25801_, _25775_);
  nor (_25803_, _08829_, _07760_);
  and (_25804_, _08829_, _07760_);
  nor (_25805_, _25804_, _25803_);
  not (_25806_, _25805_);
  not (_25807_, _08112_);
  and (_25808_, _25807_, _08114_);
  nor (_25809_, _25807_, _08114_);
  nor (_25810_, _25809_, _25808_);
  nor (_25812_, _25810_, _25806_);
  and (_25813_, _25810_, _25806_);
  nor (_25814_, _25813_, _25812_);
  and (_25815_, _25814_, _08109_);
  nor (_25816_, _25814_, _08109_);
  or (_25817_, _25816_, _25815_);
  and (_25818_, _25817_, _08107_);
  nor (_25819_, _25817_, _08107_);
  or (_25820_, _25819_, _25818_);
  and (_25821_, _25820_, _08104_);
  nor (_25823_, _25820_, _08104_);
  or (_25824_, _25823_, _25821_);
  nor (_25825_, _25824_, _07843_);
  and (_25826_, _25824_, _07843_);
  or (_25827_, _25826_, _25825_);
  or (_25828_, _25827_, _07902_);
  and (_25829_, _25828_, _07120_);
  and (_25830_, _25829_, _25802_);
  and (_25831_, _08801_, _08800_);
  nor (_25832_, _13721_, _13467_);
  and (_25834_, _13721_, _13467_);
  or (_25835_, _25834_, _25832_);
  nor (_25836_, _14333_, _14032_);
  and (_25837_, _14333_, _14032_);
  nor (_25838_, _25837_, _25836_);
  nor (_25839_, _25838_, _25835_);
  and (_25840_, _25838_, _25835_);
  nor (_25841_, _25840_, _25839_);
  not (_25842_, _25841_);
  nor (_25843_, _15234_, _14709_);
  and (_25845_, _15234_, _14709_);
  nor (_25846_, _25845_, _25843_);
  not (_25847_, _14625_);
  and (_25848_, _25847_, _07910_);
  nor (_25849_, _25847_, _07910_);
  nor (_25850_, _25849_, _25848_);
  nor (_25851_, _25850_, _25846_);
  and (_25852_, _25850_, _25846_);
  nor (_25853_, _25852_, _25851_);
  nand (_25854_, _25853_, _25842_);
  or (_25856_, _25853_, _25842_);
  and (_25857_, _25856_, _02994_);
  nand (_25858_, _25857_, _25854_);
  nand (_25859_, _25858_, _25831_);
  or (_25860_, _25859_, _25830_);
  or (_25861_, _24742_, _25831_);
  and (_25862_, _25861_, _07241_);
  and (_25863_, _25862_, _25860_);
  nor (_25864_, _07524_, _07293_);
  nor (_25865_, _13726_, _13359_);
  nor (_25867_, _25865_, _25864_);
  nor (_25868_, _25867_, _14037_);
  and (_25869_, _25867_, _14037_);
  nor (_25870_, _25869_, _25868_);
  nor (_25871_, _25870_, _14111_);
  and (_25872_, _25870_, _14111_);
  or (_25873_, _25872_, _25871_);
  nor (_25874_, _25873_, _14630_);
  and (_25875_, _25873_, _14630_);
  or (_25876_, _25875_, _25874_);
  nor (_25878_, _25876_, _14927_);
  and (_25879_, _25876_, _14927_);
  or (_25880_, _25879_, _25878_);
  and (_25881_, _25880_, _15240_);
  nor (_25882_, _25880_, _15240_);
  or (_25883_, _25882_, _25881_);
  nand (_25884_, _25883_, _07313_);
  or (_25885_, _25883_, _07313_);
  and (_25886_, _25885_, _25884_);
  and (_25887_, _25886_, _07912_);
  or (_25889_, _25887_, _07236_);
  or (_25890_, _25889_, _25863_);
  nor (_25891_, _13523_, _13367_);
  and (_25892_, _13523_, _13367_);
  or (_25893_, _25892_, _25891_);
  nor (_25894_, _25893_, _13799_);
  and (_25895_, _25893_, _13799_);
  nor (_25896_, _25895_, _25894_);
  nor (_25897_, _25896_, _14340_);
  and (_25898_, _25896_, _14340_);
  or (_25900_, _25898_, _25897_);
  nor (_25901_, _25900_, _14635_);
  and (_25902_, _25900_, _14635_);
  or (_25903_, _25902_, _25901_);
  nor (_25904_, _25903_, _14932_);
  and (_25905_, _25903_, _14932_);
  or (_25906_, _25905_, _25904_);
  nor (_25907_, _25906_, _15245_);
  and (_25908_, _25906_, _15245_);
  or (_25909_, _25908_, _25907_);
  not (_25910_, _25909_);
  nor (_25911_, _25910_, _07942_);
  and (_25912_, _25910_, _07942_);
  or (_25913_, _25912_, _25911_);
  or (_25914_, _25913_, _07917_);
  and (_25915_, _25914_, _03104_);
  and (_25916_, _25915_, _25890_);
  and (_25917_, _13733_, _13372_);
  nor (_25918_, _13733_, _13372_);
  nor (_25919_, _25918_, _25917_);
  nor (_25922_, _25919_, _14044_);
  and (_25923_, _25919_, _14044_);
  nor (_25924_, _25923_, _25922_);
  and (_25925_, _25924_, _14345_);
  nor (_25926_, _25924_, _14345_);
  or (_25927_, _25926_, _25925_);
  nor (_25928_, _25927_, _14640_);
  and (_25929_, _25927_, _14640_);
  or (_25930_, _25929_, _25928_);
  nor (_25931_, _25930_, _14937_);
  and (_25933_, _25930_, _14937_);
  or (_25934_, _25933_, _25931_);
  and (_25935_, _25934_, _15251_);
  nor (_25936_, _25934_, _15251_);
  nor (_25937_, _25936_, _25935_);
  or (_25938_, _25937_, _08023_);
  nand (_25939_, _25937_, _08023_);
  and (_25940_, _25939_, _03103_);
  and (_25941_, _25940_, _25938_);
  or (_25942_, _25941_, _07946_);
  or (_25944_, _25942_, _25916_);
  not (_25945_, _14049_);
  nor (_25946_, _13738_, _07759_);
  and (_25947_, _13738_, _07759_);
  or (_25948_, _25947_, _25946_);
  nor (_25949_, _25948_, _25945_);
  and (_25950_, _25948_, _25945_);
  nor (_25951_, _25950_, _25949_);
  and (_25952_, _25951_, _14350_);
  nor (_25953_, _25951_, _14350_);
  or (_25955_, _25953_, _25952_);
  nor (_25956_, _25955_, _14645_);
  and (_25957_, _25955_, _14645_);
  or (_25958_, _25957_, _25956_);
  nor (_25959_, _25958_, _14942_);
  and (_25960_, _25958_, _14942_);
  or (_25961_, _25960_, _25959_);
  nor (_25962_, _25961_, _15256_);
  and (_25963_, _25961_, _15256_);
  or (_25964_, _25963_, _25962_);
  and (_25966_, _25964_, _08054_);
  nor (_25967_, _25964_, _08054_);
  or (_25968_, _25967_, _25966_);
  or (_25969_, _25968_, _08029_);
  and (_25970_, _25969_, _08028_);
  and (_25971_, _25970_, _25944_);
  nor (_25972_, _07764_, _07763_);
  nor (_25973_, _13838_, \oc8051_golden_model_1.ACC [3]);
  and (_25974_, _13838_, \oc8051_golden_model_1.ACC [3]);
  nor (_25975_, _25974_, _25973_);
  and (_25977_, _25975_, _24908_);
  nor (_25978_, _25975_, _24908_);
  nor (_25979_, _25978_, _25977_);
  not (_25980_, _25979_);
  nand (_25981_, _25980_, _25972_);
  or (_25982_, _25980_, _25972_);
  and (_25983_, _25982_, _25981_);
  nand (_25984_, _25983_, _08027_);
  and (_25985_, _10309_, _03549_);
  nand (_25986_, _25985_, _25984_);
  or (_25988_, _25986_, _25971_);
  or (_25989_, _25985_, _24742_);
  and (_25990_, _25989_, _07193_);
  and (_25991_, _25990_, _25988_);
  nor (_25992_, _13286_, _07217_);
  and (_25993_, _13286_, _07217_);
  nor (_25994_, _25993_, _25992_);
  and (_25995_, _25994_, _13795_);
  nor (_25996_, _25994_, _13795_);
  nor (_25997_, _25996_, _25995_);
  and (_25999_, _25997_, _14108_);
  nor (_26000_, _25997_, _14108_);
  or (_26001_, _26000_, _25999_);
  nor (_26002_, _26001_, _14654_);
  and (_26003_, _26001_, _14654_);
  or (_26004_, _26003_, _26002_);
  nor (_26005_, _26004_, _14954_);
  and (_26006_, _26004_, _14954_);
  or (_26007_, _26006_, _26005_);
  and (_26008_, _26007_, _15267_);
  nor (_26010_, _26007_, _15267_);
  nor (_26011_, _26010_, _26008_);
  or (_26012_, _26011_, _07233_);
  nand (_26013_, _26011_, _07233_);
  and (_26014_, _26013_, _26012_);
  and (_26015_, _26014_, _13285_);
  or (_26016_, _26015_, _07183_);
  or (_26017_, _26016_, _25991_);
  not (_26018_, _07182_);
  not (_26019_, _13422_);
  and (_26020_, _26019_, _07166_);
  nor (_26021_, _26019_, _07166_);
  nor (_26022_, _26021_, _26020_);
  and (_26023_, _26022_, _14058_);
  nor (_26024_, _26022_, _14058_);
  nor (_26025_, _26024_, _26023_);
  and (_26026_, _26025_, _14361_);
  nor (_26027_, _26025_, _14361_);
  or (_26028_, _26027_, _26026_);
  and (_26029_, _26028_, _14659_);
  nor (_26032_, _26028_, _14659_);
  nor (_26033_, _26032_, _26029_);
  and (_26034_, _26033_, _14951_);
  nor (_26035_, _26033_, _14951_);
  or (_26036_, _26035_, _26034_);
  and (_26037_, _26036_, _15264_);
  nor (_26038_, _26036_, _15264_);
  nor (_26039_, _26038_, _26037_);
  and (_26040_, _26039_, _26018_);
  nor (_26041_, _26039_, _26018_);
  or (_26043_, _26041_, _08792_);
  or (_26044_, _26043_, _26040_);
  and (_26045_, _26044_, _02857_);
  and (_26046_, _26045_, _26017_);
  not (_26047_, _14063_);
  nor (_26048_, _13756_, _07684_);
  and (_26049_, _13756_, _07684_);
  or (_26050_, _26049_, _26048_);
  and (_26051_, _26050_, _26047_);
  nor (_26052_, _26050_, _26047_);
  nor (_26054_, _26052_, _26051_);
  and (_26055_, _26054_, _14367_);
  nor (_26056_, _26054_, _14367_);
  nor (_26057_, _26056_, _26055_);
  nor (_26058_, _26057_, _14664_);
  and (_26059_, _26057_, _14664_);
  or (_26060_, _26059_, _26058_);
  nor (_26061_, _26060_, _14960_);
  and (_26062_, _26060_, _14960_);
  or (_26063_, _26062_, _26061_);
  nor (_26065_, _26063_, _15005_);
  and (_26066_, _26063_, _15005_);
  or (_26067_, _26066_, _26065_);
  and (_26068_, _26067_, _08099_);
  nor (_26069_, _26067_, _08099_);
  or (_26070_, _26069_, _26068_);
  and (_26071_, _26070_, _02856_);
  or (_26072_, _26071_, _26046_);
  and (_26073_, _26072_, _08074_);
  not (_26074_, _08829_);
  and (_26076_, _26074_, _07762_);
  nor (_26077_, _26074_, _07762_);
  nor (_26078_, _26077_, _26076_);
  and (_26079_, _26078_, _14068_);
  nor (_26080_, _26078_, _14068_);
  nor (_26081_, _26080_, _26079_);
  and (_26082_, _26081_, _14373_);
  nor (_26083_, _26081_, _14373_);
  nor (_26084_, _26083_, _26082_);
  nor (_26085_, _26084_, _14669_);
  and (_26087_, _26084_, _14669_);
  or (_26088_, _26087_, _26085_);
  and (_26089_, _26088_, _14967_);
  nor (_26090_, _26088_, _14967_);
  nor (_26091_, _26090_, _26089_);
  nor (_26092_, _26091_, _15275_);
  and (_26093_, _26091_, _15275_);
  nor (_26094_, _26093_, _26092_);
  nand (_26095_, _26094_, _08132_);
  or (_26096_, _26094_, _08132_);
  and (_26098_, _26096_, _08073_);
  nand (_26099_, _26098_, _26095_);
  nand (_26100_, _26099_, _24747_);
  or (_26101_, _26100_, _26073_);
  nand (_26102_, _26101_, _24748_);
  nand (_26103_, _26102_, _05747_);
  or (_26104_, _24742_, _05747_);
  and (_26105_, _26104_, _03138_);
  and (_26106_, _26105_, _26103_);
  and (_26107_, _24944_, _03133_);
  or (_26109_, _26107_, _08138_);
  or (_26110_, _26109_, _26106_);
  not (_26111_, _08144_);
  and (_26112_, _13838_, _26111_);
  and (_26113_, _26112_, \oc8051_golden_model_1.ACC [3]);
  nor (_26114_, _26112_, \oc8051_golden_model_1.ACC [3]);
  nor (_26115_, _26114_, _26113_);
  and (_26116_, _26115_, _14682_);
  nor (_26117_, _26115_, _14682_);
  nor (_26118_, _26117_, _26116_);
  and (_26120_, _14977_, _06762_);
  nor (_26121_, _14977_, _06762_);
  nor (_26122_, _26121_, _26120_);
  nor (_26123_, _26122_, _26118_);
  and (_26124_, _26122_, _26118_);
  or (_26125_, _26124_, _26123_);
  nor (_26126_, _26125_, _08150_);
  and (_26127_, _26125_, _08150_);
  nor (_26128_, _26127_, _26126_);
  nand (_26129_, _26128_, _08138_);
  and (_26131_, _26129_, _09716_);
  and (_26132_, _26131_, _26110_);
  and (_26133_, \oc8051_golden_model_1.PSW [7], \oc8051_golden_model_1.ACC [7]);
  nor (_26134_, _26133_, _07455_);
  nand (_26135_, _26134_, _25979_);
  or (_26136_, _26134_, _25979_);
  and (_26137_, _26136_, _26135_);
  nand (_26138_, _26137_, _08143_);
  nand (_26139_, _26138_, _03907_);
  or (_26140_, _26139_, _26132_);
  or (_26142_, _24742_, _03907_);
  and (_26143_, _26142_, _03142_);
  and (_26144_, _26143_, _26140_);
  and (_26145_, _25081_, _02778_);
  or (_26146_, _26145_, _03698_);
  or (_26147_, _26146_, _26144_);
  or (_26148_, _24742_, _05214_);
  nand (_26149_, _26148_, _26147_);
  nor (_26150_, _04125_, _03912_);
  and (_26151_, _26150_, _04113_);
  nand (_26153_, _26151_, _26149_);
  or (_26154_, _26151_, _24742_);
  and (_26155_, _26154_, _02853_);
  and (_26156_, _26155_, _26153_);
  not (_26157_, _14395_);
  nor (_26158_, _14693_, _26157_);
  and (_26159_, _14693_, _26157_);
  nor (_26160_, _26159_, _26158_);
  nor (_26161_, _26160_, _15298_);
  and (_26162_, _26160_, _15298_);
  nor (_26164_, _26162_, _26161_);
  nor (_26165_, _13781_, _13330_);
  and (_26166_, _13781_, _13330_);
  nor (_26167_, _26166_, _26165_);
  and (_26168_, _26167_, _14090_);
  nor (_26169_, _26167_, _14090_);
  nor (_26170_, _26169_, _26168_);
  and (_26171_, _26170_, _14989_);
  nor (_26172_, _26170_, _14989_);
  or (_26173_, _26172_, _26171_);
  and (_26175_, _26173_, _08163_);
  nor (_26176_, _26173_, _08163_);
  or (_26177_, _26176_, _26175_);
  not (_26178_, _26177_);
  nand (_26179_, _26178_, _26164_);
  or (_26180_, _26178_, _26164_);
  and (_26181_, _26180_, _02852_);
  and (_26182_, _26181_, _26179_);
  or (_26183_, _26182_, _26156_);
  and (_26184_, _26183_, _08161_);
  not (_26186_, _08168_);
  and (_26187_, _13838_, _26186_);
  and (_26188_, _26187_, _02605_);
  nor (_26189_, _26187_, _02605_);
  nor (_26190_, _26189_, _26188_);
  nor (_26191_, _26190_, _14698_);
  and (_26192_, _26190_, _14698_);
  or (_26193_, _26192_, _26191_);
  or (_26194_, _26193_, _14994_);
  nand (_26195_, _26193_, _14994_);
  and (_26197_, _26195_, _26194_);
  or (_26198_, _26197_, _15304_);
  nand (_26199_, _26197_, _15304_);
  and (_26200_, _26199_, _26198_);
  nor (_26201_, _26200_, _08175_);
  and (_26202_, _26200_, _08175_);
  or (_26203_, _26202_, _26201_);
  nand (_26204_, _26203_, _08160_);
  nor (_26205_, _08167_, _02982_);
  and (_26206_, _26205_, _22822_);
  nand (_26208_, _26206_, _26204_);
  or (_26209_, _26208_, _26184_);
  or (_26210_, _26206_, _24742_);
  and (_26211_, _26210_, _34446_);
  and (_26212_, _26211_, _26209_);
  or (_26213_, _26212_, _24727_);
  and (_35630_[0], _26213_, _35583_);
  nand (_26214_, _04658_, _03660_);
  nor (_26215_, _04658_, \oc8051_golden_model_1.PSW [1]);
  nor (_26216_, _26215_, _05261_);
  and (_26218_, _26216_, _26214_);
  not (_26219_, _05289_);
  nor (_26220_, _10662_, _26219_);
  not (_26221_, \oc8051_golden_model_1.PSW [1]);
  nor (_26222_, _05289_, _26221_);
  or (_26223_, _26222_, _02966_);
  or (_26224_, _26223_, _26220_);
  and (_26225_, _10622_, _04658_);
  nor (_26226_, _26225_, _26215_);
  or (_26227_, _26226_, _06162_);
  not (_26229_, _02939_);
  and (_26230_, _04658_, _02477_);
  nor (_26231_, _26230_, _26215_);
  nand (_26232_, _26231_, _02837_);
  nor (_26233_, _02837_, _26221_);
  nor (_26234_, _26233_, _02932_);
  and (_26235_, _26234_, _26232_);
  nor (_26236_, _26235_, _26229_);
  and (_26237_, _26236_, _26227_);
  nor (_26238_, _04658_, _26221_);
  nor (_26240_, _09746_, _03989_);
  or (_26241_, _26240_, _26238_);
  and (_26242_, _26241_, _02930_);
  and (_26243_, _10617_, _05289_);
  or (_26244_, _26243_, _26222_);
  and (_26245_, _26244_, _02799_);
  or (_26246_, _26245_, _26242_);
  or (_26247_, _26246_, _02928_);
  or (_26248_, _26247_, _26237_);
  or (_26249_, _26231_, _02943_);
  and (_26251_, _26249_, _26248_);
  or (_26252_, _26251_, _02796_);
  and (_26253_, _10620_, _05289_);
  or (_26254_, _26253_, _26222_);
  or (_26255_, _26254_, _02927_);
  and (_26256_, _26255_, _06189_);
  and (_26257_, _26256_, _26252_);
  and (_26258_, _26243_, _10616_);
  or (_26259_, _26258_, _26222_);
  and (_26260_, _26259_, _02790_);
  or (_26262_, _26260_, _02785_);
  or (_26263_, _26262_, _26257_);
  and (_26264_, _26263_, _26224_);
  or (_26265_, _26264_, _03861_);
  or (_26266_, _26241_, _03860_);
  and (_26267_, _26266_, _26265_);
  or (_26268_, _26267_, _03850_);
  and (_26269_, _06113_, _04658_);
  or (_26270_, _26238_, _06726_);
  or (_26271_, _26270_, _26269_);
  and (_26273_, _26271_, _02970_);
  and (_26274_, _26273_, _26268_);
  nor (_26275_, _10719_, _09746_);
  or (_26276_, _26275_, _26238_);
  and (_26277_, _26276_, _02524_);
  or (_26278_, _26277_, _26274_);
  and (_26279_, _26278_, _05261_);
  or (_26280_, _26279_, _26218_);
  and (_26281_, _26280_, _03882_);
  or (_26282_, _10613_, _09746_);
  nor (_26284_, _26215_, _03881_);
  and (_26285_, _26284_, _26282_);
  or (_26286_, _10610_, _09746_);
  nor (_26287_, _26215_, _07104_);
  and (_26288_, _26287_, _26286_);
  or (_26289_, _10614_, _09746_);
  nor (_26290_, _26215_, _07092_);
  and (_26291_, _26290_, _26289_);
  or (_26292_, _26291_, _26288_);
  or (_26293_, _26292_, _26285_);
  or (_26295_, _26293_, _26281_);
  and (_26296_, _26295_, _06161_);
  or (_26297_, _26238_, _04988_);
  and (_26298_, _26231_, _03094_);
  and (_26299_, _26298_, _26297_);
  or (_26300_, _26299_, _26296_);
  and (_26301_, _26300_, _03100_);
  nand (_26302_, _26230_, _04987_);
  nor (_26303_, _26215_, _07118_);
  and (_26304_, _26303_, _26302_);
  or (_26306_, _26304_, _03133_);
  or (_26307_, _26214_, _04988_);
  nor (_26308_, _26215_, _07120_);
  and (_26309_, _26308_, _26307_);
  or (_26310_, _26309_, _26306_);
  or (_26311_, _26310_, _26301_);
  or (_26312_, _26226_, _03138_);
  and (_26313_, _26312_, _03142_);
  and (_26314_, _26313_, _26311_);
  and (_26315_, _26254_, _02778_);
  or (_26317_, _26315_, _02852_);
  or (_26318_, _26317_, _26314_);
  or (_26319_, _26238_, _02853_);
  or (_26320_, _26319_, _26225_);
  and (_26321_, _26320_, _26318_);
  or (_26322_, _26321_, _34450_);
  or (_26323_, _34446_, \oc8051_golden_model_1.PSW [1]);
  and (_26324_, _26323_, _35583_);
  and (_35630_[1], _26324_, _26322_);
  not (_26325_, \oc8051_golden_model_1.PSW [2]);
  nor (_26327_, _05289_, _26325_);
  and (_26328_, _10818_, _05289_);
  nor (_26329_, _26328_, _26327_);
  and (_26330_, _26329_, _02778_);
  nor (_26331_, _04658_, _26325_);
  not (_26332_, _26331_);
  or (_26333_, _09746_, _04413_);
  and (_26334_, _26333_, _26332_);
  and (_26335_, _26334_, _03861_);
  nor (_26336_, _10824_, _09746_);
  nor (_26338_, _26336_, _26331_);
  and (_26339_, _26338_, _02932_);
  and (_26340_, _04658_, \oc8051_golden_model_1.ACC [2]);
  nor (_26341_, _26340_, _26331_);
  or (_26342_, _26341_, _09167_);
  nor (_26343_, _02837_, _26325_);
  nor (_26344_, _26343_, _02932_);
  and (_26345_, _26344_, _26342_);
  or (_26346_, _26345_, _26229_);
  or (_26347_, _26346_, _26339_);
  or (_26349_, _26334_, _03693_);
  not (_26350_, _26327_);
  nand (_26351_, _10815_, _05289_);
  and (_26352_, _26351_, _26350_);
  or (_26353_, _26352_, _03186_);
  and (_26354_, _26353_, _26349_);
  and (_26355_, _26354_, _02943_);
  and (_26356_, _26355_, _26347_);
  and (_26357_, _26341_, _02928_);
  or (_26358_, _26357_, _26356_);
  and (_26360_, _26358_, _02927_);
  and (_26361_, _26329_, _02796_);
  or (_26362_, _26361_, _02790_);
  or (_26363_, _26362_, _26360_);
  and (_26364_, _26350_, _09771_);
  or (_26365_, _26364_, _06189_);
  or (_26366_, _26365_, _26352_);
  and (_26367_, _26366_, _26363_);
  and (_26368_, _26367_, _06201_);
  or (_26369_, _12638_, _12531_);
  or (_26371_, _26369_, _12752_);
  or (_26372_, _26371_, _12866_);
  or (_26373_, _26372_, _12982_);
  or (_26374_, _26373_, _13096_);
  or (_26375_, _26374_, _06712_);
  or (_26376_, _26375_, _13209_);
  nand (_26377_, _26376_, _07400_);
  or (_26378_, _26377_, _26368_);
  and (_26379_, _09999_, _07246_);
  nor (_26380_, _09999_, _07246_);
  or (_26382_, _26380_, _26379_);
  nor (_26383_, _26382_, _07531_);
  and (_26384_, _26382_, _07531_);
  or (_26385_, _26384_, _26383_);
  or (_26386_, _26385_, _07400_);
  and (_26387_, _26386_, _26378_);
  or (_26388_, _26387_, _07329_);
  nor (_26389_, _07334_, \oc8051_golden_model_1.ACC [7]);
  nor (_26390_, _07332_, _25590_);
  nor (_26391_, _26390_, _26389_);
  nor (_26393_, _26391_, _07338_);
  nor (_26394_, _09756_, _07333_);
  or (_26395_, _26394_, _26393_);
  nor (_26396_, _26395_, _07393_);
  and (_26397_, _26395_, _07393_);
  or (_26398_, _26397_, _26396_);
  or (_26399_, _26398_, _07330_);
  and (_26400_, _26399_, _26388_);
  or (_26401_, _26400_, _02898_);
  nor (_26402_, _10026_, _07969_);
  or (_26404_, _26402_, _07970_);
  nor (_26405_, _07960_, \oc8051_golden_model_1.ACC [7]);
  nor (_26406_, _07959_, _10130_);
  nor (_26407_, _26406_, _26405_);
  nor (_26408_, _26407_, _07965_);
  nor (_26409_, _10030_, _07961_);
  or (_26410_, _26409_, _26408_);
  nor (_26411_, _26410_, _26404_);
  and (_26412_, _26410_, _26404_);
  or (_26413_, _26412_, _02899_);
  or (_26415_, _26413_, _26411_);
  and (_26416_, _26415_, _07541_);
  and (_26417_, _26416_, _26401_);
  nor (_26418_, _07705_, _09717_);
  nor (_26419_, _07706_, \oc8051_golden_model_1.ACC [7]);
  nor (_26420_, _26419_, _26418_);
  not (_26421_, _26420_);
  or (_26422_, _26421_, _10043_);
  nand (_26423_, _26421_, _10043_);
  and (_26424_, _26423_, _26422_);
  nand (_26426_, _26424_, _07779_);
  or (_26427_, _26424_, _07779_);
  and (_26428_, _26427_, _26426_);
  and (_26429_, _26428_, _07540_);
  or (_26430_, _26429_, _02785_);
  or (_26431_, _26430_, _26417_);
  or (_26432_, _10866_, _26219_);
  and (_26433_, _26432_, _26350_);
  or (_26434_, _26433_, _02966_);
  and (_26435_, _26434_, _03860_);
  and (_26437_, _26435_, _26431_);
  or (_26438_, _26437_, _26335_);
  and (_26439_, _26438_, _06726_);
  or (_26440_, _05980_, _09746_);
  nor (_26441_, _26331_, _06726_);
  and (_26442_, _26441_, _26440_);
  or (_26443_, _26442_, _02524_);
  or (_26444_, _26443_, _26439_);
  or (_26445_, _10922_, _09746_);
  and (_26446_, _26445_, _26332_);
  or (_26448_, _26446_, _02970_);
  and (_26449_, _26448_, _06737_);
  and (_26450_, _26449_, _26444_);
  nor (_26451_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  nand (_26452_, _26451_, _06761_);
  and (_26453_, _26452_, _06731_);
  or (_26454_, _26453_, _26450_);
  and (_26455_, _26454_, _05261_);
  and (_26456_, _04658_, _05690_);
  nor (_26457_, _26456_, _26331_);
  and (_26459_, _26457_, _02974_);
  or (_26460_, _26459_, _02977_);
  or (_26461_, _26460_, _26455_);
  nand (_26462_, _10936_, _04658_);
  nor (_26463_, _26331_, _03107_);
  and (_26464_, _26463_, _26462_);
  or (_26465_, _26464_, _03108_);
  and (_26466_, _26465_, _26461_);
  nand (_26467_, _10942_, _04658_);
  nor (_26468_, _26331_, _07104_);
  and (_26469_, _26468_, _26467_);
  or (_26470_, _26469_, _02991_);
  or (_26471_, _26470_, _26466_);
  and (_26472_, _26332_, _05085_);
  or (_26473_, _26457_, _03881_);
  or (_26474_, _26473_, _26472_);
  and (_26475_, _26474_, _26471_);
  or (_26476_, _26475_, _03094_);
  or (_26477_, _26341_, _06161_);
  or (_26478_, _26477_, _26472_);
  and (_26481_, _26478_, _07120_);
  and (_26482_, _26481_, _26476_);
  or (_26483_, _10935_, _09746_);
  nor (_26484_, _26331_, _07120_);
  and (_26485_, _26484_, _26483_);
  or (_26486_, _26485_, _03099_);
  or (_26487_, _26486_, _26482_);
  or (_26488_, _10941_, _09746_);
  and (_26489_, _26488_, _26332_);
  nor (_26490_, _26489_, _07118_);
  nor (_26492_, _26490_, _10095_);
  and (_26493_, _26492_, _26487_);
  not (_26494_, _07195_);
  nor (_26495_, _07244_, _26494_);
  nor (_26496_, _07245_, \oc8051_golden_model_1.ACC [7]);
  nor (_26497_, _26496_, _09735_);
  nor (_26498_, _26497_, _26495_);
  nand (_26499_, _26498_, _07313_);
  nand (_26500_, _26495_, _07310_);
  and (_26501_, _26500_, _26499_);
  and (_26503_, _26501_, _10095_);
  or (_26504_, _26503_, _03513_);
  or (_26505_, _26504_, _26493_);
  or (_26506_, _26501_, _09732_);
  and (_26507_, _26506_, _07917_);
  and (_26508_, _26507_, _26505_);
  nor (_26509_, _26389_, _09728_);
  nor (_26510_, _26509_, _26390_);
  nand (_26511_, _26510_, _07942_);
  nand (_26512_, _26390_, _07939_);
  and (_26514_, _26512_, _07236_);
  and (_26515_, _26514_, _26511_);
  or (_26516_, _26515_, _03103_);
  or (_26517_, _26516_, _26508_);
  nand (_26518_, _26406_, _08020_);
  not (_26519_, _26407_);
  nor (_26520_, _26519_, _10105_);
  nor (_26521_, _26520_, _26406_);
  nand (_26522_, _26521_, _08023_);
  and (_26523_, _26522_, _26518_);
  or (_26525_, _26523_, _03104_);
  and (_26526_, _26525_, _08029_);
  and (_26527_, _26526_, _26517_);
  and (_26528_, _26420_, _09723_);
  or (_26529_, _26528_, _26418_);
  and (_26530_, _26529_, _08054_);
  nor (_26531_, _26529_, _08054_);
  or (_26532_, _26531_, _26530_);
  and (_26533_, _26532_, _07946_);
  or (_26534_, _26533_, _13285_);
  or (_26536_, _26534_, _26527_);
  nor (_26537_, _07230_, _07194_);
  and (_26538_, _07230_, _26494_);
  or (_26539_, _26538_, _26537_);
  or (_26540_, _26539_, _07193_);
  and (_26541_, _26540_, _08792_);
  nand (_26542_, _26541_, _26536_);
  not (_26543_, _07145_);
  nor (_26544_, _07179_, _26543_);
  and (_26545_, _07179_, _07146_);
  or (_26547_, _26545_, _08792_);
  or (_26548_, _26547_, _26544_);
  and (_26549_, _26548_, _20297_);
  and (_26550_, _26549_, _26542_);
  and (_26551_, _08129_, _09717_);
  not (_26552_, _26551_);
  and (_26553_, _26552_, _09719_);
  nor (_26554_, _08096_, _07542_);
  not (_26555_, _26554_);
  and (_26556_, _26555_, _10132_);
  nor (_26558_, _26556_, _26553_);
  not (_26559_, _26558_);
  nor (_26560_, _26559_, _26550_);
  nor (_26561_, _26560_, _03133_);
  nor (_26562_, _26338_, _03138_);
  or (_26563_, _26562_, _02778_);
  nor (_26564_, _26563_, _26561_);
  nor (_26565_, _26564_, _26330_);
  and (_26566_, _26565_, _02853_);
  and (_26567_, _10988_, _04658_);
  nor (_26569_, _26567_, _26331_);
  nor (_26570_, _26569_, _02853_);
  or (_26571_, _26570_, _26566_);
  or (_26572_, _26571_, _34450_);
  or (_26573_, _34446_, \oc8051_golden_model_1.PSW [2]);
  and (_26574_, _26573_, _35583_);
  and (_35630_[2], _26574_, _26572_);
  not (_26575_, _03095_);
  nor (_26576_, _04658_, _02937_);
  and (_26577_, _11134_, _04658_);
  nor (_26579_, _26577_, _26576_);
  nor (_26580_, _26579_, _07104_);
  nor (_26581_, _09746_, _04226_);
  nor (_26582_, _26581_, _26576_);
  and (_26583_, _26582_, _03861_);
  nor (_26584_, _11058_, _26219_);
  nor (_26585_, _05289_, _02937_);
  or (_26586_, _26585_, _02966_);
  or (_26587_, _26586_, _26584_);
  nor (_26588_, _11014_, _09746_);
  nor (_26590_, _26588_, _26576_);
  and (_26591_, _26590_, _02932_);
  and (_26592_, _04658_, \oc8051_golden_model_1.ACC [3]);
  nor (_26593_, _26592_, _26576_);
  or (_26594_, _26593_, _09167_);
  nor (_26595_, _02837_, _02937_);
  nor (_26596_, _26595_, _02932_);
  and (_26597_, _26596_, _26594_);
  or (_26598_, _26597_, _26229_);
  nor (_26599_, _26598_, _26591_);
  nor (_26601_, _26582_, _03693_);
  and (_26602_, _11011_, _05289_);
  nor (_26603_, _26602_, _26585_);
  nor (_26604_, _26603_, _03186_);
  nor (_26605_, _26604_, _26601_);
  nand (_26606_, _26605_, _02943_);
  or (_26607_, _26606_, _26599_);
  nand (_26608_, _26593_, _02928_);
  and (_26609_, _26608_, _26607_);
  and (_26610_, _26609_, _02927_);
  and (_26612_, _11009_, _05289_);
  nor (_26613_, _26612_, _26585_);
  nor (_26614_, _26613_, _02927_);
  or (_26615_, _26614_, _26610_);
  and (_26616_, _26615_, _06189_);
  or (_26617_, _26585_, _11040_);
  nor (_26618_, _26603_, _06189_);
  and (_26619_, _26618_, _26617_);
  or (_26620_, _26619_, _02785_);
  or (_26621_, _26620_, _26616_);
  and (_26623_, _26621_, _26587_);
  nor (_26624_, _26623_, _03861_);
  nor (_26625_, _26624_, _26583_);
  nor (_26626_, _26625_, _03850_);
  and (_26627_, _06116_, _04658_);
  nor (_26628_, _26576_, _06726_);
  not (_26629_, _26628_);
  nor (_26630_, _26629_, _26627_);
  or (_26631_, _26630_, _02524_);
  nor (_26632_, _26631_, _26626_);
  nor (_26634_, _11114_, _09746_);
  nor (_26635_, _26634_, _26576_);
  nor (_26636_, _26635_, _02970_);
  or (_26637_, _26636_, _02974_);
  or (_26638_, _26637_, _26632_);
  and (_26639_, _04658_, _05616_);
  nor (_26640_, _26639_, _26576_);
  nand (_26641_, _26640_, _02974_);
  and (_26642_, _26641_, _26638_);
  and (_26643_, _26642_, _07092_);
  and (_26645_, _11128_, _04658_);
  nor (_26646_, _26645_, _26576_);
  nor (_26647_, _26646_, _07092_);
  or (_26648_, _26647_, _26643_);
  and (_26649_, _26648_, _07104_);
  nor (_26650_, _26649_, _26580_);
  or (_26651_, _26650_, _26575_);
  nor (_26652_, _26576_, _04939_);
  or (_26653_, _26593_, _06161_);
  or (_26654_, _26640_, _03881_);
  and (_26656_, _26654_, _26653_);
  or (_26657_, _26656_, _26652_);
  and (_26658_, _26657_, _07120_);
  and (_26659_, _26658_, _26651_);
  nor (_26660_, _11127_, _09746_);
  or (_26661_, _26576_, _07120_);
  nor (_26662_, _26661_, _26660_);
  or (_26663_, _26662_, _03099_);
  nor (_26664_, _26663_, _26659_);
  nor (_26665_, _11133_, _09746_);
  nor (_26667_, _26665_, _26576_);
  nor (_26668_, _26667_, _07118_);
  or (_26669_, _26668_, _26664_);
  and (_26670_, _26669_, _03138_);
  nor (_26671_, _26590_, _03138_);
  or (_26672_, _26671_, _26670_);
  and (_26673_, _26672_, _03142_);
  nor (_26674_, _26613_, _03142_);
  or (_26675_, _26674_, _26673_);
  and (_26676_, _26675_, _02853_);
  and (_26678_, _11185_, _04658_);
  nor (_26679_, _26678_, _26576_);
  nor (_26680_, _26679_, _02853_);
  or (_26681_, _26680_, _26676_);
  or (_26682_, _26681_, _34450_);
  or (_26683_, _34446_, \oc8051_golden_model_1.PSW [3]);
  and (_26684_, _26683_, _35583_);
  and (_35630_[3], _26684_, _26682_);
  not (_26685_, \oc8051_golden_model_1.PSW [4]);
  nor (_26686_, _04658_, _26685_);
  and (_26688_, _11333_, _04658_);
  nor (_26689_, _26688_, _26686_);
  nor (_26690_, _26689_, _07104_);
  nor (_26691_, _05143_, _09746_);
  nor (_26692_, _26691_, _26686_);
  and (_26693_, _26692_, _03861_);
  nor (_26694_, _05289_, _26685_);
  nor (_26695_, _26694_, _11239_);
  and (_26696_, _11224_, _05289_);
  nor (_26697_, _26696_, _26694_);
  or (_26699_, _26697_, _06189_);
  nor (_26700_, _26699_, _26695_);
  nor (_26701_, _11207_, _09746_);
  nor (_26702_, _26701_, _26686_);
  and (_26703_, _26702_, _02932_);
  and (_26704_, _04658_, \oc8051_golden_model_1.ACC [4]);
  nor (_26705_, _26704_, _26686_);
  or (_26706_, _26705_, _09167_);
  nor (_26707_, _02837_, _26685_);
  nor (_26708_, _26707_, _02932_);
  and (_26710_, _26708_, _26706_);
  or (_26711_, _26710_, _26229_);
  nor (_26712_, _26711_, _26703_);
  nor (_26713_, _26692_, _03693_);
  nor (_26714_, _26697_, _03186_);
  nor (_26715_, _26714_, _26713_);
  nand (_26716_, _26715_, _02943_);
  or (_26717_, _26716_, _26712_);
  nand (_26718_, _26705_, _02928_);
  and (_26719_, _26718_, _26717_);
  and (_26721_, _26719_, _02927_);
  and (_26722_, _11203_, _05289_);
  nor (_26723_, _26722_, _26694_);
  nor (_26724_, _26723_, _02927_);
  or (_26725_, _26724_, _26721_);
  and (_26726_, _26725_, _06189_);
  nor (_26727_, _26726_, _26700_);
  nor (_26728_, _26727_, _02785_);
  nor (_26729_, _11257_, _26219_);
  nor (_26730_, _26729_, _26694_);
  nor (_26732_, _26730_, _02966_);
  nor (_26733_, _26732_, _03861_);
  not (_26734_, _26733_);
  nor (_26735_, _26734_, _26728_);
  nor (_26736_, _26735_, _26693_);
  nor (_26737_, _26736_, _03850_);
  and (_26738_, _06121_, _04658_);
  nor (_26739_, _26686_, _06726_);
  not (_26740_, _26739_);
  nor (_26741_, _26740_, _26738_);
  or (_26743_, _26741_, _02524_);
  nor (_26744_, _26743_, _26737_);
  nor (_26745_, _11313_, _09746_);
  nor (_26746_, _26745_, _26686_);
  nor (_26747_, _26746_, _02970_);
  or (_26748_, _26747_, _02974_);
  or (_26749_, _26748_, _26744_);
  and (_26750_, _05629_, _04658_);
  nor (_26751_, _26750_, _26686_);
  nand (_26752_, _26751_, _02974_);
  and (_26754_, _26752_, _26749_);
  and (_26755_, _26754_, _07092_);
  and (_26756_, _11327_, _04658_);
  nor (_26757_, _26756_, _26686_);
  nor (_26758_, _26757_, _07092_);
  or (_26759_, _26758_, _26755_);
  and (_26760_, _26759_, _07104_);
  nor (_26761_, _26760_, _26690_);
  or (_26762_, _26761_, _26575_);
  nor (_26763_, _26686_, _05190_);
  or (_26764_, _26705_, _06161_);
  or (_26765_, _26751_, _03881_);
  and (_26766_, _26765_, _26764_);
  or (_26767_, _26766_, _26763_);
  and (_26768_, _26767_, _07120_);
  and (_26769_, _26768_, _26762_);
  nor (_26770_, _11326_, _09746_);
  or (_26771_, _26686_, _07120_);
  nor (_26772_, _26771_, _26770_);
  or (_26773_, _26772_, _03099_);
  nor (_26776_, _26773_, _26769_);
  nor (_26777_, _11332_, _09746_);
  nor (_26778_, _26777_, _26686_);
  nor (_26779_, _26778_, _07118_);
  or (_26780_, _26779_, _26776_);
  and (_26781_, _26780_, _03138_);
  nor (_26782_, _26702_, _03138_);
  or (_26783_, _26782_, _26781_);
  and (_26784_, _26783_, _03142_);
  nor (_26785_, _26723_, _03142_);
  or (_26787_, _26785_, _26784_);
  and (_26788_, _26787_, _02853_);
  and (_26789_, _11383_, _04658_);
  nor (_26790_, _26789_, _26686_);
  nor (_26791_, _26790_, _02853_);
  or (_26792_, _26791_, _26788_);
  or (_26793_, _26792_, _34450_);
  or (_26794_, _34446_, \oc8051_golden_model_1.PSW [4]);
  and (_26795_, _26794_, _35583_);
  and (_35630_[4], _26795_, _26793_);
  not (_26797_, \oc8051_golden_model_1.PSW [5]);
  nor (_26798_, _04658_, _26797_);
  and (_26799_, _11531_, _04658_);
  nor (_26800_, _26799_, _26798_);
  nor (_26801_, _26800_, _07104_);
  and (_26802_, _06120_, _04658_);
  or (_26803_, _26802_, _26798_);
  and (_26804_, _26803_, _03850_);
  nor (_26805_, _11408_, _09746_);
  nor (_26806_, _26805_, _26798_);
  and (_26808_, _26806_, _02932_);
  and (_26809_, _04658_, \oc8051_golden_model_1.ACC [5]);
  nor (_26810_, _26809_, _26798_);
  or (_26811_, _26810_, _09167_);
  nor (_26812_, _02837_, _26797_);
  nor (_26813_, _26812_, _02932_);
  and (_26814_, _26813_, _26811_);
  or (_26815_, _26814_, _26229_);
  nor (_26816_, _26815_, _26808_);
  nor (_26817_, _04839_, _09746_);
  nor (_26819_, _26817_, _26798_);
  nor (_26820_, _26819_, _03693_);
  nor (_26821_, _05289_, _26797_);
  and (_26822_, _11422_, _05289_);
  nor (_26823_, _26822_, _26821_);
  nor (_26824_, _26823_, _03186_);
  nor (_26825_, _26824_, _26820_);
  nand (_26826_, _26825_, _02943_);
  or (_26827_, _26826_, _26816_);
  nand (_26828_, _26810_, _02928_);
  and (_26830_, _26828_, _26827_);
  and (_26831_, _26830_, _02927_);
  and (_26832_, _11405_, _05289_);
  nor (_26833_, _26832_, _26821_);
  nor (_26834_, _26833_, _02927_);
  or (_26835_, _26834_, _26831_);
  and (_26836_, _26835_, _06189_);
  and (_26837_, _11438_, _05289_);
  nor (_26838_, _26837_, _26821_);
  nor (_26839_, _26838_, _06189_);
  nor (_26841_, _26839_, _26836_);
  nor (_26842_, _26841_, _02785_);
  nor (_26843_, _11455_, _26219_);
  nor (_26844_, _26843_, _26821_);
  nor (_26845_, _26844_, _02966_);
  nor (_26846_, _26845_, _03861_);
  not (_26847_, _26846_);
  nor (_26848_, _26847_, _26842_);
  and (_26849_, _26819_, _03861_);
  or (_26850_, _26849_, _03850_);
  nor (_26852_, _26850_, _26848_);
  or (_26853_, _26852_, _26804_);
  and (_26854_, _26853_, _02970_);
  nor (_26855_, _11511_, _09746_);
  nor (_26856_, _26855_, _26798_);
  nor (_26857_, _26856_, _02970_);
  or (_26858_, _26857_, _02974_);
  or (_26859_, _26858_, _26854_);
  and (_26860_, _05633_, _04658_);
  nor (_26861_, _26860_, _26798_);
  nand (_26863_, _26861_, _02974_);
  and (_26864_, _26863_, _26859_);
  and (_26865_, _26864_, _07092_);
  and (_26866_, _11525_, _04658_);
  nor (_26867_, _26866_, _26798_);
  nor (_26868_, _26867_, _07092_);
  or (_26869_, _26868_, _26865_);
  and (_26870_, _26869_, _07104_);
  nor (_26871_, _26870_, _26801_);
  or (_26872_, _26871_, _26575_);
  nor (_26873_, _26798_, _04890_);
  or (_26874_, _26810_, _06161_);
  or (_26875_, _26861_, _03881_);
  and (_26876_, _26875_, _26874_);
  or (_26877_, _26876_, _26873_);
  and (_26878_, _26877_, _07120_);
  and (_26879_, _26878_, _26872_);
  nor (_26880_, _11524_, _09746_);
  or (_26881_, _26798_, _07120_);
  nor (_26882_, _26881_, _26880_);
  or (_26885_, _26882_, _03099_);
  nor (_26886_, _26885_, _26879_);
  nor (_26887_, _11530_, _09746_);
  nor (_26888_, _26887_, _26798_);
  nor (_26889_, _26888_, _07118_);
  or (_26890_, _26889_, _26886_);
  and (_26891_, _26890_, _03138_);
  nor (_26892_, _26806_, _03138_);
  or (_26893_, _26892_, _26891_);
  and (_26894_, _26893_, _03142_);
  nor (_26896_, _26833_, _03142_);
  or (_26897_, _26896_, _26894_);
  and (_26898_, _26897_, _02853_);
  and (_26899_, _11580_, _04658_);
  nor (_26900_, _26899_, _26798_);
  nor (_26901_, _26900_, _02853_);
  or (_26902_, _26901_, _26898_);
  or (_26903_, _26902_, _34450_);
  or (_26904_, _34446_, \oc8051_golden_model_1.PSW [5]);
  and (_26905_, _26904_, _35583_);
  and (_35630_[5], _26905_, _26903_);
  not (_26907_, _07702_);
  and (_26908_, _08045_, _26907_);
  nor (_26909_, _26908_, _08029_);
  not (_26910_, _07190_);
  and (_26911_, _03004_, _02591_);
  not (_26912_, _07265_);
  and (_26913_, _07304_, _26912_);
  not (_26914_, _26913_);
  and (_26915_, _26914_, _26911_);
  nor (_26917_, _04658_, _14153_);
  and (_26918_, _11601_, _04658_);
  nor (_26919_, _26918_, _26917_);
  nor (_26920_, _26919_, _07104_);
  nor (_26921_, _04735_, _09746_);
  nor (_26922_, _26921_, _26917_);
  and (_26923_, _26922_, _03861_);
  nor (_26924_, _07772_, _07702_);
  nor (_26925_, _26924_, _07541_);
  nor (_26926_, _07388_, _07352_);
  or (_26928_, _26926_, _07330_);
  or (_26929_, _07265_, _07400_);
  nor (_26930_, _26929_, _07527_);
  nor (_26931_, _11610_, _09746_);
  nor (_26932_, _26931_, _26917_);
  and (_26933_, _26932_, _02932_);
  and (_26934_, _04658_, \oc8051_golden_model_1.ACC [6]);
  nor (_26935_, _26934_, _26917_);
  or (_26936_, _26935_, _09167_);
  nor (_26937_, _02837_, _14153_);
  nor (_26939_, _26937_, _02932_);
  and (_26940_, _26939_, _26936_);
  or (_26941_, _26940_, _26229_);
  nor (_26942_, _26941_, _26933_);
  nor (_26943_, _26922_, _03693_);
  nor (_26944_, _05289_, _14153_);
  and (_26945_, _11604_, _05289_);
  nor (_26946_, _26945_, _26944_);
  nor (_26947_, _26946_, _03186_);
  nor (_26948_, _26947_, _26943_);
  nand (_26950_, _26948_, _02943_);
  or (_26951_, _26950_, _26942_);
  nand (_26952_, _26935_, _02928_);
  and (_26953_, _26952_, _26951_);
  and (_26954_, _26953_, _02927_);
  and (_26955_, _11633_, _05289_);
  nor (_26956_, _26955_, _26944_);
  nor (_26957_, _26956_, _02927_);
  or (_26958_, _26957_, _26954_);
  and (_26959_, _26958_, _06189_);
  nor (_26961_, _26944_, _11603_);
  or (_26962_, _26946_, _06189_);
  or (_26963_, _26962_, _26961_);
  and (_26964_, _26963_, _07400_);
  not (_26965_, _26964_);
  nor (_26966_, _26965_, _26959_);
  or (_26967_, _26966_, _07329_);
  or (_26968_, _26967_, _26930_);
  and (_26969_, _26968_, _02899_);
  and (_26970_, _26969_, _26928_);
  nor (_26972_, _10023_, _07956_);
  and (_26973_, _26972_, _02898_);
  nor (_26974_, _26973_, _26970_);
  and (_26975_, _26974_, _07541_);
  nor (_26976_, _26975_, _26925_);
  nor (_26977_, _26976_, _02785_);
  nor (_26978_, _11655_, _26219_);
  nor (_26979_, _26978_, _26944_);
  nor (_26980_, _26979_, _02966_);
  nor (_26981_, _26980_, _03861_);
  not (_26983_, _26981_);
  nor (_26984_, _26983_, _26977_);
  nor (_26985_, _26984_, _26923_);
  nor (_26986_, _26985_, _03850_);
  and (_26987_, _05798_, _04658_);
  nor (_26988_, _26917_, _06726_);
  not (_26989_, _26988_);
  nor (_26990_, _26989_, _26987_);
  nor (_26991_, _26990_, _02524_);
  not (_26992_, _26991_);
  nor (_26994_, _26992_, _26986_);
  nor (_26995_, _11711_, _09746_);
  nor (_26996_, _26995_, _26917_);
  nor (_26997_, _26996_, _02970_);
  or (_26998_, _26997_, _02974_);
  or (_26999_, _26998_, _26994_);
  and (_27000_, _11718_, _04658_);
  nor (_27001_, _27000_, _26917_);
  nand (_27002_, _27001_, _02974_);
  and (_27003_, _27002_, _26999_);
  and (_27005_, _27003_, _07092_);
  and (_27006_, _11728_, _04658_);
  nor (_27007_, _27006_, _26917_);
  nor (_27008_, _27007_, _07092_);
  or (_27009_, _27008_, _27005_);
  and (_27010_, _27009_, _07104_);
  nor (_27011_, _27010_, _26920_);
  or (_27012_, _27011_, _26575_);
  nor (_27013_, _26917_, _04784_);
  or (_27014_, _26935_, _06161_);
  or (_27016_, _27001_, _03881_);
  and (_27017_, _27016_, _27014_);
  or (_27018_, _27017_, _27013_);
  and (_27019_, _27018_, _07120_);
  and (_27020_, _27019_, _27012_);
  nor (_27021_, _11726_, _09746_);
  or (_27022_, _26917_, _07120_);
  nor (_27023_, _27022_, _27021_);
  nor (_27024_, _27023_, _27020_);
  nor (_27025_, _27024_, _03099_);
  nor (_27027_, _11600_, _09746_);
  nor (_27028_, _27027_, _26917_);
  and (_27029_, _27028_, _03099_);
  nor (_27030_, _27029_, _26911_);
  not (_27031_, _27030_);
  nor (_27032_, _27031_, _27025_);
  nor (_27033_, _03517_, _03251_);
  not (_27034_, _27033_);
  or (_27035_, _27034_, _27032_);
  nor (_27036_, _27035_, _26915_);
  and (_27038_, _27034_, _26913_);
  and (_27039_, _03681_, _02519_);
  nor (_27040_, _27039_, _27038_);
  not (_27041_, _27040_);
  nor (_27042_, _27041_, _27036_);
  and (_27043_, _27039_, _26914_);
  nor (_27044_, _27043_, _07240_);
  not (_27045_, _27044_);
  nor (_27046_, _27045_, _27042_);
  and (_27047_, _26913_, _07240_);
  or (_27049_, _27047_, _07236_);
  or (_27050_, _27049_, _27046_);
  not (_27051_, _07352_);
  and (_27052_, _07933_, _27051_);
  or (_27053_, _27052_, _07917_);
  and (_27054_, _27053_, _03104_);
  and (_27055_, _27054_, _27050_);
  nor (_27056_, _07956_, _03104_);
  and (_27057_, _27056_, _08014_);
  nor (_27058_, _27057_, _07946_);
  not (_27060_, _27058_);
  nor (_27061_, _27060_, _27055_);
  or (_27062_, _27061_, _26910_);
  nor (_27063_, _27062_, _26909_);
  and (_27064_, _07224_, _26910_);
  or (_27065_, _27064_, _27063_);
  and (_27066_, _27065_, _07192_);
  and (_27067_, _07224_, _07191_);
  or (_27068_, _27067_, _07183_);
  nor (_27069_, _27068_, _27066_);
  and (_27071_, _07183_, _07173_);
  nor (_27072_, _27071_, _03124_);
  not (_27073_, _27072_);
  nor (_27074_, _27073_, _27069_);
  nor (_27075_, _08090_, _03125_);
  or (_27076_, _27075_, _08073_);
  nor (_27077_, _27076_, _27074_);
  and (_27078_, _08123_, _08073_);
  or (_27079_, _27078_, _27077_);
  and (_27080_, _27079_, _03138_);
  nor (_27082_, _26932_, _03138_);
  or (_27083_, _27082_, _27080_);
  and (_27084_, _27083_, _03142_);
  nor (_27085_, _26956_, _03142_);
  or (_27086_, _27085_, _27084_);
  and (_27087_, _27086_, _02853_);
  and (_27088_, _11778_, _04658_);
  nor (_27089_, _27088_, _26917_);
  nor (_27090_, _27089_, _02853_);
  or (_27091_, _27090_, _27087_);
  or (_27092_, _27091_, _34450_);
  or (_27093_, _34446_, \oc8051_golden_model_1.PSW [6]);
  and (_27094_, _27093_, _35583_);
  and (_35630_[6], _27094_, _27092_);
  and (_35628_[0], \oc8051_golden_model_1.PCON [0], _35583_);
  and (_35628_[1], \oc8051_golden_model_1.PCON [1], _35583_);
  and (_35628_[2], \oc8051_golden_model_1.PCON [2], _35583_);
  and (_35628_[3], \oc8051_golden_model_1.PCON [3], _35583_);
  and (_35628_[4], \oc8051_golden_model_1.PCON [4], _35583_);
  and (_35628_[5], \oc8051_golden_model_1.PCON [5], _35583_);
  and (_35628_[6], \oc8051_golden_model_1.PCON [6], _35583_);
  and (_35631_[0], \oc8051_golden_model_1.SBUF [0], _35583_);
  and (_35631_[1], \oc8051_golden_model_1.SBUF [1], _35583_);
  and (_35631_[2], \oc8051_golden_model_1.SBUF [2], _35583_);
  and (_35631_[3], \oc8051_golden_model_1.SBUF [3], _35583_);
  and (_35631_[4], \oc8051_golden_model_1.SBUF [4], _35583_);
  and (_35631_[5], \oc8051_golden_model_1.SBUF [5], _35583_);
  and (_35631_[6], \oc8051_golden_model_1.SBUF [6], _35583_);
  and (_35632_[0], \oc8051_golden_model_1.SCON [0], _35583_);
  and (_35632_[1], \oc8051_golden_model_1.SCON [1], _35583_);
  and (_35632_[2], \oc8051_golden_model_1.SCON [2], _35583_);
  and (_35632_[3], \oc8051_golden_model_1.SCON [3], _35583_);
  and (_35632_[4], \oc8051_golden_model_1.SCON [4], _35583_);
  and (_35632_[5], \oc8051_golden_model_1.SCON [5], _35583_);
  and (_35632_[6], \oc8051_golden_model_1.SCON [6], _35583_);
  nor (_27098_, _04667_, _02787_);
  nor (_27099_, _05036_, _10164_);
  or (_27100_, _27099_, _27098_);
  or (_27101_, _27100_, _03330_);
  or (_27102_, _10546_, _10164_);
  nor (_27104_, _04667_, \oc8051_golden_model_1.SP [0]);
  nor (_27105_, _27104_, _07104_);
  and (_27106_, _27105_, _27102_);
  and (_27107_, _27100_, _02932_);
  not (_27108_, _27104_);
  nand (_27109_, _04667_, _02658_);
  and (_27110_, _27109_, _27108_);
  and (_27111_, _27110_, _02837_);
  nor (_27112_, _02837_, _02787_);
  or (_27113_, _27112_, _27111_);
  and (_27115_, _27113_, _06162_);
  or (_27116_, _27115_, _02930_);
  or (_27117_, _27116_, _27107_);
  and (_27118_, _04667_, _03805_);
  or (_27119_, _27118_, _27104_);
  or (_27120_, _27119_, _03693_);
  and (_27121_, _27120_, _27117_);
  or (_27122_, _27121_, _02928_);
  or (_27123_, _27110_, _02943_);
  and (_27124_, _27123_, _03932_);
  and (_27126_, _27124_, _27122_);
  nand (_27127_, _03860_, _03834_);
  or (_27128_, _27127_, _27126_);
  or (_27129_, _27098_, _03860_);
  or (_27130_, _27129_, _27118_);
  and (_27131_, _27130_, _27128_);
  or (_27132_, _27131_, _03850_);
  and (_27133_, _27132_, _02970_);
  and (_27134_, _06114_, _04667_);
  or (_27135_, _27098_, _06726_);
  or (_27137_, _27135_, _27134_);
  and (_27138_, _27137_, _27133_);
  nand (_27139_, _10530_, _04667_);
  nor (_27140_, _27104_, _02970_);
  and (_27141_, _27140_, _27139_);
  or (_27142_, _27141_, _02974_);
  or (_27143_, _27142_, _27138_);
  nand (_27144_, _04667_, _03471_);
  and (_27145_, _27144_, _27108_);
  or (_27146_, _27145_, _05261_);
  and (_27148_, _27146_, _07092_);
  and (_27149_, _27148_, _27143_);
  or (_27150_, _10427_, _10164_);
  nor (_27151_, _27104_, _07092_);
  and (_27152_, _27151_, _27150_);
  or (_27153_, _27152_, _27149_);
  and (_27154_, _27153_, _07104_);
  or (_27155_, _27154_, _27106_);
  and (_27156_, _27155_, _03095_);
  nand (_27157_, _27110_, _03094_);
  nor (_27159_, _27157_, _27099_);
  nand (_27160_, _27145_, _02991_);
  nor (_27161_, _27160_, _27099_);
  or (_27162_, _27161_, _27159_);
  or (_27163_, _27162_, _27156_);
  and (_27164_, _27163_, _03100_);
  or (_27165_, _27109_, _05036_);
  nor (_27166_, _27104_, _07118_);
  and (_27167_, _27166_, _27165_);
  or (_27168_, _27144_, _05036_);
  nor (_27170_, _27104_, _07120_);
  and (_27171_, _27170_, _27168_);
  or (_27172_, _27171_, _15390_);
  or (_27173_, _27172_, _27167_);
  or (_27174_, _27173_, _27164_);
  and (_27175_, _27174_, _27101_);
  and (_27176_, _27175_, _34446_);
  nor (_27177_, \oc8051_golden_model_1.SP [0], rst);
  nor (_27178_, _27177_, _00000_);
  or (_35633_[0], _27178_, _27176_);
  nor (_27180_, _04667_, _03692_);
  and (_27181_, _10622_, _04667_);
  nor (_27182_, _27181_, _27180_);
  nor (_27183_, _27182_, _02853_);
  or (_27184_, _10610_, _10164_);
  nor (_27185_, _04667_, \oc8051_golden_model_1.SP [1]);
  nor (_27186_, _27185_, _07104_);
  and (_27187_, _27186_, _27184_);
  nor (_27188_, _10164_, _03989_);
  or (_27189_, _27180_, _03850_);
  nor (_27191_, _27189_, _27188_);
  nor (_27192_, _27191_, _09305_);
  nor (_27193_, _27185_, _27181_);
  or (_27194_, _27193_, _06162_);
  or (_27195_, _02546_, _03692_);
  and (_27196_, _04667_, _02477_);
  nor (_27197_, _27196_, _27185_);
  and (_27198_, _27197_, _02837_);
  nor (_27199_, _02837_, _03692_);
  or (_27200_, _27199_, _02804_);
  or (_27202_, _27200_, _27198_);
  and (_27203_, _27202_, _27195_);
  or (_27204_, _27203_, _02932_);
  and (_27205_, _27204_, _02540_);
  and (_27206_, _27205_, _27194_);
  nor (_27207_, _02540_, \oc8051_golden_model_1.SP [1]);
  or (_27208_, _27207_, _02930_);
  or (_27209_, _27208_, _27206_);
  nor (_27210_, _04667_, _03927_);
  or (_27211_, _27210_, _27188_);
  or (_27213_, _27211_, _03693_);
  and (_27214_, _27213_, _27209_);
  or (_27215_, _27214_, _02928_);
  or (_27216_, _27197_, _02943_);
  and (_27217_, _27216_, _03932_);
  and (_27218_, _27217_, _27215_);
  or (_27219_, _10211_, _03931_);
  or (_27220_, _27219_, _27218_);
  or (_27221_, _04133_, _03692_);
  and (_27222_, _27221_, _03860_);
  and (_27224_, _27222_, _27220_);
  or (_27225_, _27224_, _27192_);
  and (_27226_, _06113_, _04667_);
  or (_27227_, _27180_, _06726_);
  or (_27228_, _27227_, _27226_);
  and (_27229_, _27228_, _02970_);
  and (_27230_, _27229_, _27225_);
  nor (_27231_, _10719_, _10164_);
  or (_27232_, _27231_, _27180_);
  and (_27233_, _27232_, _02524_);
  or (_27235_, _27233_, _27230_);
  and (_27236_, _27235_, _05261_);
  nand (_27237_, _04667_, _03660_);
  nor (_27238_, _27185_, _05261_);
  and (_27239_, _27238_, _27237_);
  or (_27240_, _27239_, _02585_);
  or (_27241_, _27240_, _27236_);
  and (_27242_, _02585_, \oc8051_golden_model_1.SP [1]);
  nor (_27243_, _27242_, _02977_);
  and (_27244_, _27243_, _27241_);
  or (_27246_, _10614_, _10164_);
  nor (_27247_, _27185_, _07092_);
  and (_27248_, _27247_, _27246_);
  or (_27249_, _27248_, _27244_);
  and (_27250_, _27249_, _07104_);
  or (_27251_, _27250_, _27187_);
  and (_27252_, _27251_, _03881_);
  or (_27253_, _10613_, _10164_);
  nor (_27254_, _27185_, _03881_);
  and (_27255_, _27254_, _27253_);
  or (_27257_, _27255_, _27252_);
  and (_27258_, _27257_, _08809_);
  and (_27259_, _02594_, _03692_);
  or (_27260_, _27180_, _04988_);
  and (_27261_, _27197_, _03094_);
  and (_27262_, _27261_, _27260_);
  or (_27263_, _27262_, _27259_);
  or (_27264_, _27263_, _27258_);
  and (_27265_, _27264_, _03100_);
  or (_27266_, _27237_, _04988_);
  nor (_27268_, _27185_, _07120_);
  and (_27269_, _27268_, _27266_);
  nand (_27270_, _27196_, _04987_);
  nor (_27271_, _27185_, _07118_);
  and (_27272_, _27271_, _27270_);
  or (_27273_, _27272_, _27269_);
  or (_27274_, _27273_, _27265_);
  and (_27275_, _27274_, _10309_);
  nor (_27276_, _10309_, \oc8051_golden_model_1.SP [1]);
  nor (_27277_, _27276_, _02854_);
  not (_27279_, _27277_);
  nor (_27280_, _27279_, _27275_);
  and (_27281_, _02854_, \oc8051_golden_model_1.SP [1]);
  nor (_27282_, _27281_, _03133_);
  not (_27283_, _27282_);
  nor (_27284_, _27283_, _27280_);
  nor (_27285_, _27193_, _04331_);
  nor (_27286_, _27285_, _10372_);
  nor (_27287_, _27286_, _27284_);
  nor (_27288_, _03907_, _03692_);
  nor (_27290_, _27288_, _02852_);
  not (_27291_, _27290_);
  nor (_27292_, _27291_, _27287_);
  nor (_27293_, _27292_, _27183_);
  nor (_27294_, _27293_, _34450_);
  nor (_27295_, \oc8051_golden_model_1.SP [1], rst);
  nor (_27296_, _27295_, _00000_);
  or (_35633_[1], _27296_, _27294_);
  and (_27297_, _10988_, _04667_);
  nor (_27298_, _04667_, _03256_);
  or (_27300_, _27298_, _02853_);
  or (_27301_, _27300_, _27297_);
  and (_27302_, _10942_, _04667_);
  or (_27303_, _27302_, _27298_);
  and (_27304_, _27303_, _03107_);
  nand (_27305_, _12141_, _02585_);
  nor (_27306_, _10164_, _04413_);
  or (_27307_, _27298_, _03860_);
  or (_27308_, _27307_, _27306_);
  nor (_27309_, _10824_, _10164_);
  or (_27311_, _27309_, _27298_);
  or (_27312_, _27311_, _06162_);
  and (_27313_, _04667_, \oc8051_golden_model_1.ACC [2]);
  or (_27314_, _27313_, _27298_);
  or (_27315_, _27314_, _09167_);
  or (_27316_, _02837_, \oc8051_golden_model_1.SP [2]);
  and (_27317_, _27316_, _02546_);
  and (_27318_, _27317_, _27315_);
  and (_27319_, _04505_, _02804_);
  or (_27320_, _27319_, _02932_);
  or (_27322_, _27320_, _27318_);
  and (_27323_, _27322_, _02540_);
  and (_27324_, _27323_, _27312_);
  nor (_27325_, _12141_, _02540_);
  or (_27326_, _27325_, _02930_);
  or (_27327_, _27326_, _27324_);
  nor (_27328_, _05358_, _04667_);
  or (_27329_, _27328_, _27306_);
  or (_27330_, _27329_, _03693_);
  and (_27331_, _27330_, _27327_);
  or (_27332_, _27331_, _02928_);
  or (_27333_, _27314_, _02943_);
  and (_27334_, _27333_, _03932_);
  and (_27335_, _27334_, _27332_);
  or (_27336_, _27335_, _04357_);
  and (_27337_, _27336_, _04133_);
  or (_27338_, _12141_, _04133_);
  nand (_27339_, _27338_, _03860_);
  or (_27340_, _27339_, _27337_);
  and (_27341_, _27340_, _27308_);
  or (_27344_, _27341_, _03850_);
  and (_27345_, _06117_, _04667_);
  or (_27346_, _27298_, _06726_);
  or (_27347_, _27346_, _27345_);
  and (_27348_, _27347_, _02970_);
  and (_27349_, _27348_, _27344_);
  nor (_27350_, _10922_, _10164_);
  or (_27351_, _27350_, _27298_);
  and (_27352_, _27351_, _02524_);
  or (_27353_, _27352_, _02974_);
  or (_27355_, _27353_, _27349_);
  and (_27356_, _04667_, _05690_);
  or (_27357_, _27356_, _27298_);
  or (_27358_, _27357_, _05261_);
  and (_27359_, _27358_, _27355_);
  or (_27360_, _27359_, _02585_);
  and (_27361_, _27360_, _27305_);
  or (_27362_, _27361_, _02977_);
  and (_27363_, _10936_, _04667_);
  or (_27364_, _27298_, _07092_);
  or (_27366_, _27364_, _27363_);
  and (_27367_, _27366_, _07104_);
  and (_27368_, _27367_, _27362_);
  or (_27369_, _27368_, _27304_);
  and (_27370_, _27369_, _03881_);
  or (_27371_, _27298_, _05086_);
  and (_27372_, _27357_, _02991_);
  and (_27373_, _27372_, _27371_);
  or (_27374_, _27373_, _27370_);
  and (_27375_, _27374_, _08809_);
  and (_27377_, _04505_, _02594_);
  or (_27378_, _27377_, _02994_);
  and (_27379_, _27314_, _03094_);
  and (_27380_, _27379_, _27371_);
  or (_27381_, _27380_, _27378_);
  or (_27382_, _27381_, _27375_);
  nor (_27383_, _10935_, _10164_);
  or (_27384_, _27383_, _27298_);
  or (_27385_, _27384_, _07120_);
  and (_27386_, _27385_, _27382_);
  or (_27388_, _27386_, _03099_);
  nor (_27389_, _10941_, _10164_);
  or (_27390_, _27298_, _07118_);
  or (_27391_, _27390_, _27389_);
  and (_27392_, _27391_, _10159_);
  and (_27393_, _27392_, _27388_);
  and (_27394_, _12141_, _03113_);
  or (_27395_, _27394_, _02592_);
  or (_27396_, _27395_, _27393_);
  nand (_27397_, _12141_, _02592_);
  and (_27399_, _27397_, _02855_);
  and (_27400_, _27399_, _27396_);
  and (_27401_, _12141_, _02854_);
  or (_27402_, _27401_, _03133_);
  or (_27403_, _27402_, _27400_);
  or (_27404_, _27311_, _03138_);
  and (_27405_, _27404_, _03907_);
  and (_27406_, _27405_, _27403_);
  nor (_27407_, _12141_, _03907_);
  or (_27408_, _27407_, _02852_);
  or (_27410_, _27408_, _27406_);
  and (_27411_, _27410_, _27301_);
  and (_27412_, _27411_, _34446_);
  nor (_27413_, \oc8051_golden_model_1.SP [2], rst);
  nor (_27414_, _27413_, _00000_);
  or (_35633_[2], _27414_, _27412_);
  nor (_27415_, _04667_, _03129_);
  and (_27416_, _11185_, _04667_);
  nor (_27417_, _27416_, _27415_);
  nor (_27418_, _27417_, _02853_);
  and (_27420_, _11134_, _04667_);
  nor (_27421_, _27420_, _27415_);
  nor (_27422_, _27421_, _07104_);
  and (_27423_, _11954_, _02585_);
  nor (_27424_, _10164_, _04226_);
  or (_27425_, _27415_, _03850_);
  nor (_27426_, _27425_, _27424_);
  nor (_27427_, _27426_, _09305_);
  nor (_27428_, _02837_, _03129_);
  and (_27429_, _04667_, \oc8051_golden_model_1.ACC [3]);
  nor (_27431_, _27429_, _27415_);
  nor (_27432_, _27431_, _09167_);
  or (_27433_, _27432_, _27428_);
  and (_27434_, _27433_, _02546_);
  and (_27435_, _04508_, _02804_);
  nor (_27436_, _27435_, _27434_);
  nor (_27437_, _27436_, _02932_);
  nor (_27438_, _11014_, _10164_);
  nor (_27439_, _27438_, _27415_);
  nor (_27440_, _27439_, _06162_);
  or (_27442_, _27440_, _27437_);
  and (_27443_, _27442_, _02540_);
  nor (_27444_, _11954_, _02540_);
  or (_27445_, _27444_, _27443_);
  and (_27446_, _27445_, _03693_);
  nor (_27447_, _05346_, _04667_);
  nor (_27448_, _27447_, _27424_);
  nor (_27449_, _27448_, _03693_);
  or (_27450_, _27449_, _27446_);
  and (_27451_, _27450_, _02943_);
  nor (_27453_, _27431_, _02943_);
  or (_27454_, _27453_, _27451_);
  and (_27455_, _27454_, _03932_);
  or (_27456_, _27455_, _10211_);
  nor (_27457_, _27456_, _04277_);
  nor (_27458_, _04508_, _04133_);
  or (_27459_, _27458_, _03861_);
  nor (_27460_, _27459_, _27457_);
  nor (_27461_, _27460_, _27427_);
  and (_27462_, _06116_, _04667_);
  nor (_27464_, _27415_, _06726_);
  not (_27465_, _27464_);
  nor (_27466_, _27465_, _27462_);
  or (_27467_, _27466_, _02524_);
  nor (_27468_, _27467_, _27461_);
  nor (_27469_, _11114_, _10164_);
  nor (_27470_, _27469_, _27415_);
  nor (_27471_, _27470_, _02970_);
  or (_27472_, _27471_, _02974_);
  or (_27473_, _27472_, _27468_);
  and (_27475_, _04667_, _05616_);
  nor (_27476_, _27475_, _27415_);
  nand (_27477_, _27476_, _02974_);
  and (_27478_, _27477_, _27473_);
  nor (_27479_, _27478_, _02585_);
  nor (_27480_, _27479_, _27423_);
  and (_27481_, _27480_, _07092_);
  and (_27482_, _11128_, _04667_);
  nor (_27483_, _27482_, _27415_);
  nor (_27484_, _27483_, _07092_);
  or (_27486_, _27484_, _27481_);
  and (_27487_, _27486_, _07104_);
  nor (_27488_, _27487_, _27422_);
  nor (_27489_, _27488_, _02991_);
  nor (_27490_, _27415_, _04939_);
  not (_27491_, _27490_);
  nor (_27492_, _27476_, _03881_);
  and (_27493_, _27492_, _27491_);
  nor (_27494_, _27493_, _27489_);
  nor (_27495_, _27494_, _10160_);
  and (_27497_, _04508_, _02594_);
  or (_27498_, _27490_, _06161_);
  nor (_27499_, _27498_, _27431_);
  nor (_27500_, _27499_, _27497_);
  and (_27501_, _27500_, _07120_);
  not (_27502_, _27501_);
  nor (_27503_, _27502_, _27495_);
  nor (_27504_, _11127_, _10164_);
  nor (_27505_, _27504_, _27415_);
  and (_27506_, _27505_, _02994_);
  nor (_27508_, _27506_, _27503_);
  and (_27509_, _27508_, _07118_);
  nor (_27510_, _11133_, _10164_);
  nor (_27511_, _27510_, _27415_);
  nor (_27512_, _27511_, _07118_);
  or (_27513_, _27512_, _27509_);
  and (_27514_, _27513_, _10159_);
  nor (_27515_, _05343_, _03129_);
  nor (_27516_, _27515_, _05344_);
  nor (_27517_, _27516_, _10159_);
  or (_27519_, _27517_, _02592_);
  nor (_27520_, _27519_, _27514_);
  and (_27521_, _11954_, _02592_);
  nor (_27522_, _27521_, _27520_);
  and (_27523_, _27522_, _02855_);
  nor (_27524_, _27516_, _02855_);
  or (_27525_, _27524_, _27523_);
  and (_27526_, _27525_, _03138_);
  nor (_27527_, _27439_, _03138_);
  or (_27528_, _27527_, _04331_);
  nor (_27530_, _27528_, _27526_);
  nor (_27531_, _04508_, _03907_);
  nor (_27532_, _27531_, _02852_);
  not (_27533_, _27532_);
  nor (_27534_, _27533_, _27530_);
  nor (_27535_, _27534_, _27418_);
  nand (_27536_, _27535_, _34446_);
  or (_27537_, _34446_, \oc8051_golden_model_1.SP [3]);
  and (_27538_, _27537_, _35583_);
  and (_35633_[3], _27538_, _27536_);
  nor (_27540_, _04667_, _10195_);
  and (_27541_, _11383_, _04667_);
  nor (_27542_, _27541_, _27540_);
  nor (_27543_, _27542_, _02853_);
  nor (_27544_, _04235_, \oc8051_golden_model_1.SP [4]);
  nor (_27545_, _27544_, _10175_);
  and (_27546_, _27545_, _02594_);
  nor (_27547_, _27546_, _02994_);
  and (_27548_, _11333_, _04667_);
  nor (_27549_, _27548_, _27540_);
  nor (_27551_, _27549_, _07104_);
  nor (_27552_, _05143_, _10164_);
  or (_27553_, _27540_, _03850_);
  nor (_27554_, _27553_, _27552_);
  nor (_27555_, _27554_, _09305_);
  nor (_27556_, _04236_, _10195_);
  and (_27557_, _04236_, _10195_);
  nor (_27558_, _27557_, _27556_);
  and (_27559_, _27558_, _02795_);
  nor (_27560_, _02837_, _10195_);
  and (_27562_, _04667_, \oc8051_golden_model_1.ACC [4]);
  nor (_27563_, _27562_, _27540_);
  nor (_27564_, _27563_, _09167_);
  or (_27565_, _27564_, _27560_);
  and (_27566_, _27565_, _02546_);
  and (_27567_, _27545_, _02804_);
  nor (_27568_, _27567_, _27566_);
  nor (_27569_, _27568_, _02932_);
  nor (_27570_, _11207_, _10164_);
  nor (_27571_, _27570_, _27540_);
  nor (_27573_, _27571_, _06162_);
  or (_27574_, _27573_, _27569_);
  and (_27575_, _27574_, _02540_);
  not (_27576_, _27545_);
  nor (_27577_, _27576_, _02540_);
  or (_27578_, _27577_, _27575_);
  and (_27579_, _27578_, _03693_);
  and (_27580_, _10196_, _02787_);
  nor (_27581_, _05345_, _10195_);
  nor (_27582_, _27581_, _27580_);
  nor (_27584_, _27582_, _04667_);
  nor (_27585_, _27584_, _27552_);
  nor (_27586_, _27585_, _03693_);
  or (_27587_, _27586_, _27579_);
  and (_27588_, _27587_, _02943_);
  nor (_27589_, _27563_, _02943_);
  or (_27590_, _27589_, _27588_);
  and (_27591_, _27590_, _03932_);
  or (_27592_, _27591_, _10211_);
  nor (_27593_, _27592_, _27559_);
  nor (_27595_, _27545_, _04133_);
  or (_27596_, _27595_, _03861_);
  nor (_27597_, _27596_, _27593_);
  nor (_27598_, _27597_, _27555_);
  and (_27599_, _06121_, _04667_);
  nor (_27600_, _27540_, _06726_);
  not (_27601_, _27600_);
  nor (_27602_, _27601_, _27599_);
  or (_27603_, _27602_, _02524_);
  nor (_27604_, _27603_, _27598_);
  nor (_27606_, _11313_, _10164_);
  nor (_27607_, _27606_, _27540_);
  nor (_27608_, _27607_, _02970_);
  or (_27609_, _27608_, _02974_);
  or (_27610_, _27609_, _27604_);
  and (_27611_, _05629_, _04667_);
  nor (_27612_, _27611_, _27540_);
  nand (_27613_, _27612_, _02974_);
  and (_27614_, _27613_, _27610_);
  nor (_27615_, _27614_, _02585_);
  and (_27616_, _27576_, _02585_);
  nor (_27617_, _27616_, _27615_);
  and (_27618_, _27617_, _07092_);
  and (_27619_, _11327_, _04667_);
  nor (_27620_, _27619_, _27540_);
  nor (_27621_, _27620_, _07092_);
  or (_27622_, _27621_, _27618_);
  and (_27623_, _27622_, _07104_);
  nor (_27624_, _27623_, _27551_);
  nor (_27625_, _27624_, _02991_);
  nor (_27628_, _27540_, _05190_);
  not (_27629_, _27628_);
  nor (_27630_, _27612_, _03881_);
  and (_27631_, _27630_, _27629_);
  nor (_27632_, _27631_, _27625_);
  nor (_27633_, _27632_, _10160_);
  nor (_27634_, _27563_, _06161_);
  and (_27635_, _27634_, _27629_);
  nor (_27636_, _27635_, _27633_);
  and (_27637_, _27636_, _27547_);
  nor (_27639_, _11326_, _10164_);
  nor (_27640_, _27639_, _27540_);
  and (_27641_, _27640_, _02994_);
  nor (_27642_, _27641_, _27637_);
  and (_27643_, _27642_, _07118_);
  nor (_27644_, _11332_, _10164_);
  nor (_27645_, _27644_, _27540_);
  nor (_27646_, _27645_, _07118_);
  or (_27647_, _27646_, _27643_);
  and (_27648_, _27647_, _10159_);
  nor (_27650_, _05344_, _10195_);
  nor (_27651_, _27650_, _10196_);
  nor (_27652_, _27651_, _10159_);
  or (_27653_, _27652_, _02592_);
  nor (_27654_, _27653_, _27648_);
  and (_27655_, _27576_, _02592_);
  nor (_27656_, _27655_, _27654_);
  and (_27657_, _27656_, _02855_);
  nor (_27658_, _27651_, _02855_);
  or (_27659_, _27658_, _27657_);
  and (_27661_, _27659_, _03138_);
  nor (_27662_, _27571_, _03138_);
  or (_27663_, _27662_, _04331_);
  nor (_27664_, _27663_, _27661_);
  nor (_27665_, _27545_, _03907_);
  nor (_27666_, _27665_, _02852_);
  not (_27667_, _27666_);
  nor (_27668_, _27667_, _27664_);
  nor (_27669_, _27668_, _27543_);
  nand (_27670_, _27669_, _34446_);
  or (_27672_, _34446_, \oc8051_golden_model_1.SP [4]);
  and (_27673_, _27672_, _35583_);
  and (_35633_[4], _27673_, _27670_);
  nor (_27674_, _04667_, _10194_);
  and (_27675_, _11580_, _04667_);
  nor (_27676_, _27675_, _27674_);
  nor (_27677_, _27676_, _02853_);
  nor (_27678_, _27674_, _04890_);
  not (_27679_, _27678_);
  and (_27680_, _05633_, _04667_);
  nor (_27682_, _27680_, _27674_);
  nor (_27683_, _27682_, _03881_);
  and (_27684_, _27683_, _27679_);
  and (_27685_, _10176_, \oc8051_golden_model_1.SP [0]);
  nor (_27686_, _27556_, \oc8051_golden_model_1.SP [5]);
  nor (_27687_, _27686_, _27685_);
  and (_27688_, _27687_, _02795_);
  nor (_27689_, _02837_, _10194_);
  and (_27690_, _04667_, \oc8051_golden_model_1.ACC [5]);
  nor (_27691_, _27690_, _27674_);
  nor (_27693_, _27691_, _09167_);
  or (_27694_, _27693_, _27689_);
  and (_27695_, _27694_, _02546_);
  nor (_27696_, _10175_, \oc8051_golden_model_1.SP [5]);
  nor (_27697_, _27696_, _10176_);
  and (_27698_, _27697_, _02804_);
  nor (_27699_, _27698_, _27695_);
  nor (_27700_, _27699_, _02932_);
  nor (_27701_, _11408_, _10164_);
  nor (_27702_, _27701_, _27674_);
  nor (_27704_, _27702_, _06162_);
  or (_27705_, _27704_, _27700_);
  and (_27706_, _27705_, _02540_);
  not (_27707_, _27697_);
  nor (_27708_, _27707_, _02540_);
  or (_27709_, _27708_, _27706_);
  and (_27710_, _27709_, _03693_);
  nor (_27711_, _04839_, _10164_);
  and (_27712_, _10197_, _02787_);
  nor (_27713_, _27580_, _10194_);
  nor (_27715_, _27713_, _27712_);
  nor (_27716_, _27715_, _04667_);
  nor (_27717_, _27716_, _27711_);
  nor (_27718_, _27717_, _03693_);
  or (_27719_, _27718_, _27710_);
  and (_27720_, _27719_, _02943_);
  nor (_27721_, _27691_, _02943_);
  or (_27722_, _27721_, _27720_);
  and (_27723_, _27722_, _03932_);
  or (_27724_, _27723_, _10211_);
  nor (_27726_, _27724_, _27688_);
  nor (_27727_, _27697_, _04133_);
  or (_27728_, _27727_, _27726_);
  and (_27729_, _27728_, _03860_);
  nor (_27730_, _27674_, _03860_);
  not (_27731_, _27730_);
  nor (_27732_, _27731_, _27711_);
  nor (_27733_, _27732_, _27729_);
  nor (_27734_, _27733_, _03850_);
  and (_27735_, _06120_, _04667_);
  nor (_27737_, _27674_, _06726_);
  not (_27738_, _27737_);
  nor (_27739_, _27738_, _27735_);
  nor (_27740_, _27739_, _27734_);
  nor (_27741_, _27740_, _02524_);
  nor (_27742_, _11511_, _10164_);
  nor (_27743_, _27742_, _27674_);
  and (_27744_, _27743_, _02524_);
  nor (_27745_, _27744_, _27741_);
  and (_27746_, _27745_, _05261_);
  nor (_27748_, _27682_, _05261_);
  or (_27749_, _27748_, _27746_);
  and (_27750_, _27749_, _04131_);
  and (_27751_, _27697_, _02585_);
  or (_27752_, _27751_, _27750_);
  and (_27753_, _27752_, _07092_);
  and (_27754_, _11525_, _04667_);
  nor (_27755_, _27754_, _27674_);
  nor (_27756_, _27755_, _07092_);
  or (_27757_, _27756_, _27753_);
  and (_27759_, _27757_, _07104_);
  and (_27760_, _11531_, _04667_);
  nor (_27761_, _27760_, _27674_);
  nor (_27762_, _27761_, _07104_);
  or (_27763_, _27762_, _27759_);
  and (_27764_, _27763_, _03881_);
  nor (_27765_, _27764_, _27684_);
  nor (_27766_, _27765_, _10160_);
  nor (_27767_, _27691_, _06161_);
  and (_27768_, _27767_, _27679_);
  and (_27770_, _27697_, _02594_);
  nor (_27771_, _27770_, _27768_);
  and (_27772_, _27771_, _07120_);
  not (_27773_, _27772_);
  nor (_27774_, _27773_, _27766_);
  nor (_27775_, _11524_, _10164_);
  or (_27776_, _27674_, _07120_);
  nor (_27777_, _27776_, _27775_);
  nor (_27778_, _27777_, _27774_);
  and (_27779_, _27778_, _07118_);
  nor (_27781_, _11530_, _10164_);
  nor (_27782_, _27781_, _27674_);
  nor (_27783_, _27782_, _07118_);
  or (_27784_, _27783_, _27779_);
  and (_27785_, _27784_, _10159_);
  nor (_27786_, _10196_, _10194_);
  nor (_27787_, _27786_, _10197_);
  nor (_27788_, _27787_, _10159_);
  or (_27789_, _27788_, _02592_);
  nor (_27790_, _27789_, _27785_);
  and (_27792_, _27707_, _02592_);
  nor (_27793_, _27792_, _27790_);
  and (_27794_, _27793_, _02855_);
  nor (_27795_, _27787_, _02855_);
  or (_27796_, _27795_, _27794_);
  and (_27797_, _27796_, _03138_);
  nor (_27798_, _27702_, _03138_);
  or (_27799_, _27798_, _04331_);
  nor (_27800_, _27799_, _27797_);
  nor (_27801_, _27697_, _03907_);
  nor (_27803_, _27801_, _02852_);
  not (_27804_, _27803_);
  nor (_27805_, _27804_, _27800_);
  nor (_27806_, _27805_, _27677_);
  nand (_27807_, _27806_, _34446_);
  or (_27808_, _34446_, \oc8051_golden_model_1.SP [5]);
  and (_27809_, _27808_, _35583_);
  and (_35633_[5], _27809_, _27807_);
  and (_27810_, _11778_, _04667_);
  nor (_27811_, _04667_, _10193_);
  or (_27813_, _27811_, _02853_);
  or (_27814_, _27813_, _27810_);
  and (_27815_, _11601_, _04667_);
  or (_27816_, _27815_, _27811_);
  and (_27817_, _27816_, _03107_);
  nor (_27818_, _04735_, _10164_);
  or (_27819_, _27811_, _03860_);
  or (_27820_, _27819_, _27818_);
  nor (_27821_, _11610_, _10164_);
  or (_27822_, _27821_, _27811_);
  or (_27824_, _27822_, _06162_);
  and (_27825_, _04667_, \oc8051_golden_model_1.ACC [6]);
  or (_27826_, _27825_, _27811_);
  or (_27827_, _27826_, _09167_);
  or (_27828_, _02837_, \oc8051_golden_model_1.SP [6]);
  and (_27829_, _27828_, _02546_);
  and (_27830_, _27829_, _27827_);
  nor (_27831_, _10176_, \oc8051_golden_model_1.SP [6]);
  nor (_27832_, _27831_, _10177_);
  and (_27833_, _27832_, _02804_);
  or (_27835_, _27833_, _02932_);
  or (_27836_, _27835_, _27830_);
  and (_27837_, _27836_, _02540_);
  and (_27838_, _27837_, _27824_);
  and (_27839_, _27832_, _04239_);
  or (_27840_, _27839_, _02930_);
  or (_27841_, _27840_, _27838_);
  nor (_27842_, _27712_, _10193_);
  nor (_27843_, _27842_, _10199_);
  nor (_27844_, _27843_, _04667_);
  or (_27846_, _27844_, _27818_);
  or (_27847_, _27846_, _03693_);
  and (_27848_, _27847_, _27841_);
  or (_27849_, _27848_, _02928_);
  or (_27850_, _27826_, _02943_);
  and (_27851_, _27850_, _03932_);
  and (_27852_, _27851_, _27849_);
  nor (_27853_, _27685_, \oc8051_golden_model_1.SP [6]);
  nor (_27854_, _27853_, _10212_);
  and (_27855_, _27854_, _02795_);
  or (_27857_, _27855_, _27852_);
  and (_27858_, _27857_, _04133_);
  nand (_27859_, _27832_, _10211_);
  nand (_27860_, _27859_, _03860_);
  or (_27861_, _27860_, _27858_);
  and (_27862_, _27861_, _27820_);
  or (_27863_, _27862_, _03850_);
  and (_27864_, _05798_, _04667_);
  or (_27865_, _27864_, _06726_);
  or (_27866_, _27865_, _27811_);
  and (_27868_, _27866_, _02970_);
  and (_27869_, _27868_, _27863_);
  nor (_27870_, _11711_, _10164_);
  or (_27871_, _27870_, _27811_);
  and (_27872_, _27871_, _02524_);
  or (_27873_, _27872_, _02974_);
  or (_27874_, _27873_, _27869_);
  and (_27875_, _11718_, _04667_);
  or (_27876_, _27875_, _27811_);
  or (_27877_, _27876_, _05261_);
  and (_27879_, _27877_, _27874_);
  or (_27880_, _27879_, _02585_);
  or (_27881_, _27832_, _04131_);
  and (_27882_, _27881_, _27880_);
  or (_27883_, _27882_, _02977_);
  and (_27884_, _11728_, _04667_);
  or (_27885_, _27811_, _07092_);
  or (_27886_, _27885_, _27884_);
  and (_27887_, _27886_, _07104_);
  and (_27888_, _27887_, _27883_);
  or (_27890_, _27888_, _27817_);
  and (_27891_, _27890_, _03881_);
  or (_27892_, _27811_, _04784_);
  and (_27893_, _27876_, _02991_);
  and (_27894_, _27893_, _27892_);
  or (_27895_, _27894_, _27891_);
  and (_27896_, _27895_, _08809_);
  and (_27897_, _27826_, _03094_);
  and (_27898_, _27897_, _27892_);
  and (_27899_, _27832_, _02594_);
  or (_27901_, _27899_, _02994_);
  or (_27902_, _27901_, _27898_);
  or (_27903_, _27902_, _27896_);
  nor (_27904_, _11726_, _10164_);
  or (_27905_, _27904_, _27811_);
  or (_27906_, _27905_, _07120_);
  and (_27907_, _27906_, _27903_);
  or (_27908_, _27907_, _03099_);
  nor (_27909_, _11600_, _10164_);
  or (_27910_, _27811_, _07118_);
  or (_27912_, _27910_, _27909_);
  and (_27913_, _27912_, _10159_);
  and (_27914_, _27913_, _27908_);
  nor (_27915_, _10197_, _10193_);
  or (_27916_, _27915_, _10198_);
  and (_27917_, _27916_, _03113_);
  or (_27918_, _27917_, _02592_);
  or (_27919_, _27918_, _27914_);
  or (_27920_, _27832_, _05741_);
  and (_27921_, _27920_, _02855_);
  and (_27923_, _27921_, _27919_);
  and (_27924_, _27916_, _02854_);
  or (_27925_, _27924_, _03133_);
  or (_27926_, _27925_, _27923_);
  or (_27927_, _27822_, _03138_);
  and (_27928_, _27927_, _03907_);
  and (_27929_, _27928_, _27926_);
  and (_27930_, _27832_, _04331_);
  or (_27931_, _27930_, _02852_);
  or (_27932_, _27931_, _27929_);
  and (_27934_, _27932_, _27814_);
  or (_27935_, _27934_, _34450_);
  or (_27936_, _34446_, \oc8051_golden_model_1.SP [6]);
  and (_27937_, _27936_, _35583_);
  and (_35633_[6], _27937_, _27935_);
  and (_35634_[0], \oc8051_golden_model_1.TCON [0], _35583_);
  and (_35634_[1], \oc8051_golden_model_1.TCON [1], _35583_);
  and (_35634_[2], \oc8051_golden_model_1.TCON [2], _35583_);
  and (_35634_[3], \oc8051_golden_model_1.TCON [3], _35583_);
  and (_35634_[4], \oc8051_golden_model_1.TCON [4], _35583_);
  and (_35634_[5], \oc8051_golden_model_1.TCON [5], _35583_);
  and (_35634_[6], \oc8051_golden_model_1.TCON [6], _35583_);
  and (_35635_[0], \oc8051_golden_model_1.TH0 [0], _35583_);
  and (_35635_[1], \oc8051_golden_model_1.TH0 [1], _35583_);
  and (_35635_[2], \oc8051_golden_model_1.TH0 [2], _35583_);
  and (_35635_[3], \oc8051_golden_model_1.TH0 [3], _35583_);
  and (_35635_[4], \oc8051_golden_model_1.TH0 [4], _35583_);
  and (_35635_[5], \oc8051_golden_model_1.TH0 [5], _35583_);
  and (_35635_[6], \oc8051_golden_model_1.TH0 [6], _35583_);
  and (_35636_[0], \oc8051_golden_model_1.TH1 [0], _35583_);
  and (_35636_[1], \oc8051_golden_model_1.TH1 [1], _35583_);
  and (_35636_[2], \oc8051_golden_model_1.TH1 [2], _35583_);
  and (_35636_[3], \oc8051_golden_model_1.TH1 [3], _35583_);
  and (_35636_[4], \oc8051_golden_model_1.TH1 [4], _35583_);
  and (_35636_[5], \oc8051_golden_model_1.TH1 [5], _35583_);
  and (_35636_[6], \oc8051_golden_model_1.TH1 [6], _35583_);
  and (_35637_[0], \oc8051_golden_model_1.TL0 [0], _35583_);
  and (_35637_[1], \oc8051_golden_model_1.TL0 [1], _35583_);
  and (_35637_[2], \oc8051_golden_model_1.TL0 [2], _35583_);
  and (_35637_[3], \oc8051_golden_model_1.TL0 [3], _35583_);
  and (_35637_[4], \oc8051_golden_model_1.TL0 [4], _35583_);
  and (_35637_[5], \oc8051_golden_model_1.TL0 [5], _35583_);
  and (_35637_[6], \oc8051_golden_model_1.TL0 [6], _35583_);
  and (_35638_[0], \oc8051_golden_model_1.TL1 [0], _35583_);
  and (_35638_[1], \oc8051_golden_model_1.TL1 [1], _35583_);
  and (_35638_[2], \oc8051_golden_model_1.TL1 [2], _35583_);
  and (_35638_[3], \oc8051_golden_model_1.TL1 [3], _35583_);
  and (_35638_[4], \oc8051_golden_model_1.TL1 [4], _35583_);
  and (_35638_[5], \oc8051_golden_model_1.TL1 [5], _35583_);
  and (_35638_[6], \oc8051_golden_model_1.TL1 [6], _35583_);
  and (_35639_[0], \oc8051_golden_model_1.TMOD [0], _35583_);
  and (_35639_[1], \oc8051_golden_model_1.TMOD [1], _35583_);
  and (_35639_[2], \oc8051_golden_model_1.TMOD [2], _35583_);
  and (_35639_[3], \oc8051_golden_model_1.TMOD [3], _35583_);
  and (_35639_[4], \oc8051_golden_model_1.TMOD [4], _35583_);
  and (_35639_[5], \oc8051_golden_model_1.TMOD [5], _35583_);
  and (_35639_[6], \oc8051_golden_model_1.TMOD [6], _35583_);
  and (_27942_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [0]);
  and (_27943_, _07425_, \oc8051_golden_model_1.DPL [0]);
  nor (_27944_, _07425_, _09178_);
  or (_27946_, _09162_, _07432_);
  and (_27947_, _27946_, _03805_);
  and (_27948_, _20718_, _09158_);
  and (_27949_, _09156_, \oc8051_golden_model_1.DPL [0]);
  and (_27950_, _09168_, _09163_);
  and (_27951_, _10364_, \oc8051_golden_model_1.XRAM_ADDR [0]);
  and (_27952_, _27951_, _27950_);
  or (_27953_, _27952_, _27949_);
  and (_27954_, _27953_, _27948_);
  or (_27955_, _27954_, _27947_);
  and (_27957_, _27955_, _27944_);
  or (_27958_, _27957_, _27943_);
  and (_27959_, _10312_, _05324_);
  and (_27960_, _27959_, _10324_);
  and (_27961_, _10304_, _09927_);
  and (_27962_, _27961_, _27960_);
  and (_27963_, _09319_, _05268_);
  and (_27964_, _27963_, _10326_);
  and (_27965_, _10332_, _07808_);
  and (_27966_, _27965_, _10351_);
  and (_27968_, _27966_, _27964_);
  and (_27969_, _27968_, _27962_);
  and (_27970_, _09289_, _07330_);
  and (_27971_, _27970_, _10331_);
  and (_27972_, _27971_, _09759_);
  and (_27973_, _27972_, _07400_);
  and (_27974_, _27973_, _10308_);
  and (_27975_, _27974_, _10344_);
  and (_27976_, _27975_, _27969_);
  and (_27977_, _10382_, _10370_);
  and (_27979_, _10358_, _10328_);
  nor (_27980_, _03236_, _02990_);
  and (_27981_, _10316_, _10296_);
  nor (_27982_, _07191_, _07185_);
  and (_27983_, _27982_, _07189_);
  and (_27984_, _27983_, _27981_);
  and (_27985_, _27984_, _19640_);
  and (_27986_, _27985_, _27980_);
  and (_27987_, _10346_, _02571_);
  nor (_27988_, _27987_, _03557_);
  not (_27990_, _06081_);
  and (_27991_, _10753_, _27990_);
  and (_27992_, _27991_, _27988_);
  and (_27993_, _27992_, _27986_);
  and (_27994_, _10310_, _10371_);
  not (_27995_, _03260_);
  and (_27996_, _25985_, _08028_);
  and (_27997_, _27996_, _27995_);
  and (_27998_, _10373_, _03560_);
  and (_27999_, _27998_, _27997_);
  and (_28001_, _27999_, _27994_);
  and (_28002_, _28001_, _27993_);
  and (_28003_, _28002_, _27979_);
  and (_28004_, _28003_, _27977_);
  and (_28005_, _28004_, _27976_);
  and (_28006_, _28005_, _27958_);
  or (_28007_, _28006_, _27942_);
  and (_35640_[0], _28007_, _35583_);
  and (_28008_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [1]);
  and (_28009_, _07425_, \oc8051_golden_model_1.DPL [1]);
  and (_28010_, _27946_, _03990_);
  and (_28011_, _09156_, \oc8051_golden_model_1.DPL [1]);
  and (_28012_, _10364_, \oc8051_golden_model_1.XRAM_ADDR [1]);
  and (_28013_, _28012_, _27950_);
  or (_28014_, _28013_, _28011_);
  and (_28015_, _28014_, _27948_);
  or (_28016_, _28015_, _28010_);
  and (_28017_, _28016_, _27944_);
  or (_28018_, _28017_, _28009_);
  and (_28019_, _28018_, _28005_);
  or (_28022_, _28019_, _28008_);
  and (_35640_[1], _28022_, _35583_);
  and (_28023_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [2]);
  and (_28024_, _07425_, \oc8051_golden_model_1.DPL [2]);
  and (_28025_, _27946_, _04414_);
  and (_28026_, _09156_, \oc8051_golden_model_1.DPL [2]);
  and (_28027_, _10364_, \oc8051_golden_model_1.XRAM_ADDR [2]);
  and (_28028_, _28027_, _27950_);
  or (_28029_, _28028_, _28026_);
  and (_28030_, _28029_, _27948_);
  or (_28032_, _28030_, _28025_);
  and (_28033_, _28032_, _27944_);
  or (_28034_, _28033_, _28024_);
  and (_28035_, _28034_, _28005_);
  or (_28036_, _28035_, _28023_);
  and (_35640_[2], _28036_, _35583_);
  and (_28037_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [3]);
  and (_28038_, _07425_, \oc8051_golden_model_1.DPL [3]);
  and (_28039_, _27946_, _07272_);
  and (_28040_, _09156_, \oc8051_golden_model_1.DPL [3]);
  and (_28042_, _10364_, \oc8051_golden_model_1.XRAM_ADDR [3]);
  and (_28043_, _28042_, _27950_);
  or (_28044_, _28043_, _28040_);
  and (_28045_, _28044_, _27948_);
  or (_28046_, _28045_, _28039_);
  and (_28047_, _28046_, _27944_);
  or (_28048_, _28047_, _28038_);
  and (_28049_, _28048_, _28005_);
  or (_28050_, _28049_, _28037_);
  and (_35640_[3], _28050_, _35583_);
  and (_28052_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [4]);
  and (_28053_, _07425_, \oc8051_golden_model_1.DPL [4]);
  and (_28054_, _27946_, _05200_);
  and (_28055_, _09156_, \oc8051_golden_model_1.DPL [4]);
  and (_28056_, _10364_, \oc8051_golden_model_1.XRAM_ADDR [4]);
  and (_28057_, _28056_, _27950_);
  or (_28058_, _28057_, _28055_);
  and (_28059_, _28058_, _27948_);
  or (_28060_, _28059_, _28054_);
  and (_28061_, _28060_, _27944_);
  or (_28063_, _28061_, _28053_);
  and (_28064_, _28063_, _28005_);
  or (_28065_, _28064_, _28052_);
  and (_35640_[4], _28065_, _35583_);
  and (_28066_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [5]);
  and (_28067_, _07425_, \oc8051_golden_model_1.DPL [5]);
  and (_28068_, _27946_, _05199_);
  and (_28069_, _09156_, \oc8051_golden_model_1.DPL [5]);
  and (_28070_, _10364_, \oc8051_golden_model_1.XRAM_ADDR [5]);
  and (_28071_, _28070_, _27950_);
  or (_28073_, _28071_, _28069_);
  and (_28074_, _28073_, _27948_);
  or (_28075_, _28074_, _28068_);
  and (_28076_, _28075_, _27944_);
  or (_28077_, _28076_, _28067_);
  and (_28078_, _28077_, _28005_);
  or (_28079_, _28078_, _28066_);
  and (_35640_[5], _28079_, _35583_);
  and (_28080_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [6]);
  and (_28081_, _07425_, \oc8051_golden_model_1.DPL [6]);
  and (_28083_, _27946_, _07242_);
  and (_28084_, _09156_, \oc8051_golden_model_1.DPL [6]);
  and (_28085_, _10364_, \oc8051_golden_model_1.XRAM_ADDR [6]);
  and (_28086_, _28085_, _27950_);
  or (_28087_, _28086_, _28084_);
  and (_28088_, _28087_, _27948_);
  or (_28089_, _28088_, _28083_);
  and (_28090_, _28089_, _27944_);
  or (_28091_, _28090_, _28081_);
  and (_28092_, _28091_, _28005_);
  or (_28094_, _28092_, _28080_);
  and (_35640_[6], _28094_, _35583_);
  and (_28095_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [7]);
  and (_28096_, _07425_, \oc8051_golden_model_1.DPL [7]);
  and (_28097_, _27946_, _05198_);
  and (_28098_, _09156_, \oc8051_golden_model_1.DPL [7]);
  and (_28099_, _10364_, \oc8051_golden_model_1.XRAM_ADDR [7]);
  and (_28100_, _28099_, _27950_);
  or (_28101_, _28100_, _28098_);
  and (_28102_, _28101_, _27948_);
  or (_28104_, _28102_, _28097_);
  and (_28105_, _28104_, _27944_);
  or (_28106_, _28105_, _28096_);
  and (_28107_, _28106_, _28005_);
  or (_28108_, _28107_, _28095_);
  and (_35640_[7], _28108_, _35583_);
  and (_28109_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [8]);
  and (_28110_, _10362_, \oc8051_golden_model_1.DPH [0]);
  and (_28111_, _02545_, \oc8051_golden_model_1.XRAM_ADDR [8]);
  and (_28112_, _28111_, _02543_);
  or (_28114_, _28112_, _28110_);
  and (_28115_, _28114_, _28004_);
  and (_28116_, _28115_, _27976_);
  or (_28117_, _28116_, _28109_);
  and (_35640_[8], _28117_, _35583_);
  and (_28118_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [9]);
  and (_28119_, _10377_, _10378_);
  and (_28120_, _27962_, _28119_);
  and (_28121_, _10308_, _10331_);
  and (_28122_, _27966_, _28121_);
  and (_28124_, _27963_, _10380_);
  and (_28125_, _27970_, _10753_);
  and (_28126_, _28125_, _27980_);
  and (_28127_, _28126_, _27999_);
  not (_28128_, _27987_);
  and (_28129_, _10756_, _28128_);
  and (_28130_, _28129_, _10328_);
  and (_28131_, _28130_, _28127_);
  and (_28132_, _28131_, _28124_);
  and (_28133_, _28132_, _28122_);
  and (_28135_, _10362_, \oc8051_golden_model_1.DPH [1]);
  and (_28136_, _02545_, \oc8051_golden_model_1.XRAM_ADDR [9]);
  and (_28137_, _28136_, _02543_);
  or (_28138_, _28137_, _28135_);
  and (_28139_, _10345_, _07400_);
  and (_28140_, _10370_, _10358_);
  and (_28141_, _27994_, _10326_);
  and (_28142_, _27985_, _28141_);
  and (_28143_, _28142_, _28140_);
  and (_28144_, _28143_, _28139_);
  and (_28146_, _28144_, _28138_);
  and (_28147_, _28146_, _28133_);
  and (_28148_, _28147_, _28120_);
  or (_28149_, _28148_, _28118_);
  and (_35640_[9], _28149_, _35583_);
  and (_28150_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [10]);
  and (_28151_, _27974_, _27998_);
  and (_28152_, _28151_, _27993_);
  and (_28153_, _28152_, _27977_);
  and (_28154_, _10362_, \oc8051_golden_model_1.DPH [2]);
  and (_28156_, _02545_, \oc8051_golden_model_1.XRAM_ADDR [10]);
  and (_28157_, _28156_, _02543_);
  or (_28158_, _28157_, _28154_);
  and (_28159_, _27994_, _10352_);
  and (_28160_, _27997_, _10328_);
  and (_28161_, _28160_, _28159_);
  and (_28162_, _28161_, _10357_);
  and (_28163_, _28162_, _10344_);
  and (_28164_, _28163_, _27969_);
  and (_28165_, _28164_, _28158_);
  and (_28167_, _28165_, _28153_);
  or (_28168_, _28167_, _28150_);
  and (_35640_[10], _28168_, _35583_);
  and (_28169_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [11]);
  and (_28170_, _10362_, \oc8051_golden_model_1.DPH [3]);
  and (_28171_, _02545_, \oc8051_golden_model_1.XRAM_ADDR [11]);
  and (_28172_, _28171_, _02543_);
  or (_28173_, _28172_, _28170_);
  and (_28174_, _28173_, _28004_);
  and (_28175_, _28174_, _27976_);
  or (_28177_, _28175_, _28169_);
  and (_35640_[11], _28177_, _35583_);
  and (_28178_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [12]);
  and (_28179_, _10362_, \oc8051_golden_model_1.DPH [4]);
  and (_28180_, _02545_, \oc8051_golden_model_1.XRAM_ADDR [12]);
  and (_28181_, _28180_, _02543_);
  or (_28182_, _28181_, _28179_);
  and (_28183_, _28182_, _28005_);
  or (_28184_, _28183_, _28178_);
  and (_35640_[12], _28184_, _35583_);
  and (_28185_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [13]);
  and (_28186_, _10362_, \oc8051_golden_model_1.DPH [5]);
  and (_28187_, _02545_, \oc8051_golden_model_1.XRAM_ADDR [13]);
  and (_28188_, _28187_, _02543_);
  or (_28189_, _28188_, _28186_);
  and (_28190_, _28189_, _28005_);
  or (_28191_, _28190_, _28185_);
  and (_35640_[13], _28191_, _35583_);
  and (_28192_, _34450_, \oc8051_golden_model_1.XRAM_ADDR [14]);
  and (_28193_, _10362_, \oc8051_golden_model_1.DPH [6]);
  and (_28196_, _02545_, \oc8051_golden_model_1.XRAM_ADDR [14]);
  and (_28197_, _28196_, _02543_);
  or (_28198_, _28197_, _28193_);
  and (_28199_, _28198_, _28164_);
  and (_28200_, _28199_, _28153_);
  or (_28201_, _28200_, _28192_);
  and (_35640_[14], _28201_, _35583_);
  and (_28202_, _34450_, \oc8051_golden_model_1.XRAM_DATA_OUT [0]);
  and (_28203_, _09162_, \oc8051_golden_model_1.ACC [0]);
  and (_28204_, _27950_, \oc8051_golden_model_1.XRAM_DATA_OUT [0]);
  or (_28206_, _28204_, _28203_);
  and (_28207_, _28206_, _10364_);
  and (_28208_, _09156_, \oc8051_golden_model_1.ACC [0]);
  or (_28209_, _28208_, _28207_);
  and (_28210_, _27986_, _10304_);
  and (_28211_, _28210_, _28209_);
  and (_28212_, _27991_, _27994_);
  and (_28213_, _10328_, _09927_);
  and (_28214_, _28213_, _27988_);
  and (_28215_, _28214_, _10326_);
  and (_28217_, _28215_, _09158_);
  and (_28218_, _28217_, _27999_);
  and (_28219_, _28218_, _28212_);
  and (_28220_, _27944_, _20718_);
  and (_28221_, _28220_, _27960_);
  and (_28222_, _28221_, _27963_);
  and (_28223_, _28222_, _28219_);
  and (_28224_, _28223_, _10358_);
  and (_28225_, _28224_, _28211_);
  and (_28226_, _28225_, _28122_);
  and (_28227_, _28139_, _27970_);
  and (_28228_, _27977_, _28227_);
  and (_28229_, _28228_, _28226_);
  or (_28230_, _28229_, _28202_);
  and (_35642_[0], _28230_, _35583_);
  and (_28231_, _34450_, \oc8051_golden_model_1.XRAM_DATA_OUT [1]);
  and (_28232_, _10382_, _10358_);
  and (_28233_, _27968_, _10344_);
  and (_28234_, _28233_, _28232_);
  and (_28235_, _27960_, _02543_);
  and (_28237_, _28235_, _27961_);
  and (_28238_, _24746_, _20297_);
  and (_28239_, _28238_, _08794_);
  and (_28240_, _28239_, _05748_);
  and (_28241_, _27994_, _10373_);
  and (_28242_, _28241_, _10328_);
  and (_28243_, _27996_, _03544_);
  and (_28244_, _28243_, _28242_);
  and (_28245_, _28244_, _28240_);
  and (_28246_, _28245_, _10370_);
  and (_28248_, _09162_, \oc8051_golden_model_1.ACC [1]);
  and (_28249_, _27950_, \oc8051_golden_model_1.XRAM_DATA_OUT [1]);
  or (_28250_, _28249_, _28248_);
  and (_28251_, _28250_, _10364_);
  and (_28252_, _09156_, \oc8051_golden_model_1.ACC [1]);
  or (_28253_, _28252_, _28251_);
  and (_28254_, _28253_, _27974_);
  and (_28255_, _28254_, _28246_);
  and (_28256_, _28255_, _28237_);
  and (_28257_, _28256_, _28234_);
  or (_28259_, _28257_, _28231_);
  and (_35642_[1], _28259_, _35583_);
  and (_28260_, _34450_, \oc8051_golden_model_1.XRAM_DATA_OUT [2]);
  and (_28261_, _28245_, _10344_);
  and (_28262_, _09162_, \oc8051_golden_model_1.ACC [2]);
  and (_28263_, _27950_, \oc8051_golden_model_1.XRAM_DATA_OUT [2]);
  or (_28264_, _28263_, _28262_);
  and (_28265_, _28264_, _10364_);
  and (_28266_, _09156_, \oc8051_golden_model_1.ACC [2]);
  or (_28267_, _28266_, _28265_);
  and (_28269_, _28267_, _27974_);
  and (_28270_, _28269_, _28261_);
  and (_28271_, _28270_, _10382_);
  and (_28272_, _28140_, _27968_);
  and (_28273_, _28272_, _28237_);
  and (_28274_, _28273_, _28271_);
  or (_28275_, _28274_, _28260_);
  and (_35642_[2], _28275_, _35583_);
  and (_28276_, _34450_, \oc8051_golden_model_1.XRAM_DATA_OUT [3]);
  and (_28277_, _10319_, _05261_);
  and (_28279_, _28277_, _09158_);
  and (_28280_, _10328_, _10354_);
  and (_28281_, _28280_, _09927_);
  and (_28282_, _28281_, _28243_);
  and (_28283_, _28282_, _28279_);
  and (_28284_, _28241_, _10326_);
  and (_28285_, _28240_, _28284_);
  and (_28286_, _28285_, _28283_);
  and (_28287_, _28286_, _28221_);
  and (_28288_, _10356_, _10352_);
  and (_28290_, _09162_, \oc8051_golden_model_1.ACC [3]);
  and (_28291_, _27950_, \oc8051_golden_model_1.XRAM_DATA_OUT [3]);
  or (_28292_, _28291_, _28290_);
  and (_28293_, _28292_, _10364_);
  and (_28294_, _09156_, \oc8051_golden_model_1.ACC [3]);
  or (_28295_, _28294_, _28293_);
  and (_28296_, _28295_, _28288_);
  and (_28297_, _28296_, _28287_);
  and (_28298_, _10381_, _10306_);
  and (_28299_, _28298_, _28297_);
  and (_28301_, _10377_, _10370_);
  and (_28302_, _28122_, _10349_);
  and (_28303_, _28302_, _28301_);
  and (_28304_, _28303_, _28299_);
  or (_28305_, _28304_, _28276_);
  and (_35642_[3], _28305_, _35583_);
  and (_28306_, _34450_, \oc8051_golden_model_1.XRAM_DATA_OUT [4]);
  and (_28307_, _27964_, _10351_);
  and (_28308_, _28307_, _28288_);
  and (_28309_, _28308_, _10381_);
  and (_28311_, _28241_, _27965_);
  and (_28312_, _28243_, _28311_);
  and (_28313_, _28281_, _27944_);
  and (_28314_, _28313_, _27948_);
  and (_28315_, _28240_, _27960_);
  and (_28316_, _28315_, _28314_);
  and (_28317_, _28316_, _28312_);
  and (_28318_, _10344_, _10304_);
  and (_28319_, _09162_, \oc8051_golden_model_1.ACC [4]);
  and (_28320_, _27950_, \oc8051_golden_model_1.XRAM_DATA_OUT [4]);
  or (_28322_, _28320_, _28319_);
  and (_28323_, _28322_, _10364_);
  and (_28324_, _09156_, \oc8051_golden_model_1.ACC [4]);
  or (_28325_, _28324_, _28323_);
  and (_28326_, _28325_, _27974_);
  and (_28327_, _28326_, _28318_);
  and (_28328_, _28327_, _28317_);
  and (_28329_, _28328_, _28301_);
  and (_28330_, _28329_, _28309_);
  or (_28331_, _28330_, _28306_);
  and (_35642_[4], _28331_, _35583_);
  and (_28333_, _34450_, \oc8051_golden_model_1.XRAM_DATA_OUT [5]);
  and (_28334_, _09162_, \oc8051_golden_model_1.ACC [5]);
  and (_28335_, _27950_, \oc8051_golden_model_1.XRAM_DATA_OUT [5]);
  or (_28336_, _28335_, _28334_);
  and (_28337_, _28336_, _10364_);
  and (_28338_, _09156_, \oc8051_golden_model_1.ACC [5]);
  or (_28339_, _28338_, _28337_);
  and (_28340_, _27974_, _28245_);
  and (_28341_, _28340_, _28339_);
  and (_28343_, _28341_, _10370_);
  and (_28344_, _28343_, _28237_);
  and (_28345_, _28344_, _28234_);
  or (_28346_, _28345_, _28333_);
  and (_35642_[5], _28346_, _35583_);
  and (_28347_, _34450_, \oc8051_golden_model_1.XRAM_DATA_OUT [6]);
  and (_28348_, _09162_, \oc8051_golden_model_1.ACC [6]);
  and (_28349_, _27950_, \oc8051_golden_model_1.XRAM_DATA_OUT [6]);
  or (_28350_, _28349_, _28348_);
  and (_28351_, _28350_, _10364_);
  and (_28353_, _09156_, \oc8051_golden_model_1.ACC [6]);
  or (_28354_, _28353_, _28351_);
  and (_28355_, _28235_, _25083_);
  and (_28356_, _28355_, _28354_);
  and (_28357_, _28280_, _27971_);
  and (_28358_, _28357_, _07400_);
  and (_28359_, _28358_, _28240_);
  and (_28360_, _28359_, _10303_);
  and (_28361_, _28312_, _10308_);
  and (_28362_, _28361_, _28360_);
  and (_28364_, _28362_, _10345_);
  and (_28365_, _28364_, _28356_);
  and (_28366_, _28365_, _28301_);
  and (_28367_, _28366_, _28309_);
  or (_28368_, _28367_, _28347_);
  and (_35642_[6], _28368_, _35583_);
  and (_28369_, _34450_, \oc8051_golden_model_1.P0INREG [0]);
  or (_28370_, _28369_, _00536_);
  and (_35620_[0], _28370_, _35583_);
  and (_28371_, _34450_, \oc8051_golden_model_1.P0INREG [1]);
  or (_28373_, _28371_, _00569_);
  and (_35620_[1], _28373_, _35583_);
  and (_28374_, _34450_, \oc8051_golden_model_1.P0INREG [2]);
  or (_28375_, _28374_, _00552_);
  and (_35620_[2], _28375_, _35583_);
  and (_28376_, _34450_, \oc8051_golden_model_1.P0INREG [3]);
  or (_28377_, _28376_, _00521_);
  and (_35620_[3], _28377_, _35583_);
  and (_28378_, _34450_, \oc8051_golden_model_1.P0INREG [4]);
  or (_28379_, _28378_, _00529_);
  and (_35620_[4], _28379_, _35583_);
  and (_28381_, _34450_, \oc8051_golden_model_1.P0INREG [5]);
  or (_28382_, _28381_, _00562_);
  and (_35620_[5], _28382_, _35583_);
  and (_28383_, _34450_, \oc8051_golden_model_1.P0INREG [6]);
  or (_28384_, _28383_, _00545_);
  and (_35620_[6], _28384_, _35583_);
  and (_28385_, _34450_, \oc8051_golden_model_1.P1INREG [0]);
  or (_28386_, _28385_, _00452_);
  and (_35622_[0], _28386_, _35583_);
  and (_28388_, _34450_, \oc8051_golden_model_1.P1INREG [1]);
  or (_28389_, _28388_, _00476_);
  and (_35622_[1], _28389_, _35583_);
  and (_28390_, _34450_, \oc8051_golden_model_1.P1INREG [2]);
  or (_28391_, _28390_, _00492_);
  and (_35622_[2], _28391_, _35583_);
  and (_28392_, _34450_, \oc8051_golden_model_1.P1INREG [3]);
  or (_28393_, _28392_, _00461_);
  and (_35622_[3], _28393_, _35583_);
  and (_28394_, _34450_, \oc8051_golden_model_1.P1INREG [4]);
  or (_28396_, _28394_, _00445_);
  and (_35622_[4], _28396_, _35583_);
  and (_28397_, _34450_, \oc8051_golden_model_1.P1INREG [5]);
  or (_28398_, _28397_, _00469_);
  and (_35622_[5], _28398_, _35583_);
  and (_28399_, _34450_, \oc8051_golden_model_1.P1INREG [6]);
  or (_28400_, _28399_, _00485_);
  and (_35622_[6], _28400_, _35583_);
  and (_28401_, _34450_, \oc8051_golden_model_1.P2INREG [0]);
  or (_28402_, _28401_, _00618_);
  and (_35624_[0], _28402_, _35583_);
  and (_28404_, _34450_, \oc8051_golden_model_1.P2INREG [1]);
  or (_28405_, _28404_, _00659_);
  and (_35624_[1], _28405_, _35583_);
  and (_28406_, _34450_, \oc8051_golden_model_1.P2INREG [2]);
  or (_28407_, _28406_, _00643_);
  and (_35624_[2], _28407_, _35583_);
  and (_28408_, _34450_, \oc8051_golden_model_1.P2INREG [3]);
  or (_28409_, _28408_, _00627_);
  and (_35624_[3], _28409_, _35583_);
  and (_28411_, _34450_, \oc8051_golden_model_1.P2INREG [4]);
  or (_28412_, _28411_, _00611_);
  and (_35624_[4], _28412_, _35583_);
  and (_28413_, _34450_, \oc8051_golden_model_1.P2INREG [5]);
  or (_28414_, _28413_, _00652_);
  and (_35624_[5], _28414_, _35583_);
  and (_28415_, _34450_, \oc8051_golden_model_1.P2INREG [6]);
  or (_28416_, _28415_, _00636_);
  and (_35624_[6], _28416_, _35583_);
  and (_28417_, _34450_, \oc8051_golden_model_1.P3INREG [0]);
  or (_28419_, _28417_, _00710_);
  and (_35626_[0], _28419_, _35583_);
  and (_28420_, _34450_, \oc8051_golden_model_1.P3INREG [1]);
  or (_28421_, _28420_, _00751_);
  and (_35626_[1], _28421_, _35583_);
  and (_28422_, _34450_, \oc8051_golden_model_1.P3INREG [2]);
  or (_28423_, _28422_, _00735_);
  and (_35626_[2], _28423_, _35583_);
  and (_28424_, _34450_, \oc8051_golden_model_1.P3INREG [3]);
  or (_28425_, _28424_, _00719_);
  and (_35626_[3], _28425_, _35583_);
  and (_28427_, _34450_, \oc8051_golden_model_1.P3INREG [4]);
  or (_28428_, _28427_, _00703_);
  and (_35626_[4], _28428_, _35583_);
  and (_28429_, _34450_, \oc8051_golden_model_1.P3INREG [5]);
  or (_28430_, _28429_, _00744_);
  and (_35626_[5], _28430_, _35583_);
  and (_28431_, _34450_, \oc8051_golden_model_1.P3INREG [6]);
  or (_28432_, _28431_, _00728_);
  and (_35626_[6], _28432_, _35583_);
  and (_35641_[0], \oc8051_golden_model_1.XRAM_DATA_IN [0], _35583_);
  and (_35641_[1], \oc8051_golden_model_1.XRAM_DATA_IN [1], _35583_);
  and (_35641_[2], \oc8051_golden_model_1.XRAM_DATA_IN [2], _35583_);
  and (_35641_[3], \oc8051_golden_model_1.XRAM_DATA_IN [3], _35583_);
  and (_35641_[4], \oc8051_golden_model_1.XRAM_DATA_IN [4], _35583_);
  and (_35641_[5], \oc8051_golden_model_1.XRAM_DATA_IN [5], _35583_);
  and (_35641_[6], \oc8051_golden_model_1.XRAM_DATA_IN [6], _35583_);
  and (_00005_[6], _00729_, _35583_);
  and (_00005_[5], _00745_, _35583_);
  and (_00005_[4], _00704_, _35583_);
  and (_00005_[3], _00720_, _35583_);
  and (_00005_[2], _00736_, _35583_);
  and (_00005_[1], _00752_, _35583_);
  and (_00005_[0], _00711_, _35583_);
  and (_00004_[6], _00637_, _35583_);
  and (_00004_[5], _00653_, _35583_);
  and (_00004_[4], _00612_, _35583_);
  and (_00004_[3], _00628_, _35583_);
  and (_00004_[2], _00644_, _35583_);
  and (_00004_[1], _00660_, _35583_);
  and (_00004_[0], _00619_, _35583_);
  and (_00003_[6], _00486_, _35583_);
  and (_00003_[5], _00470_, _35583_);
  and (_00003_[4], _00446_, _35583_);
  and (_00003_[3], _00462_, _35583_);
  and (_00003_[2], _00493_, _35583_);
  and (_00003_[1], _00477_, _35583_);
  and (_00003_[0], _00453_, _35583_);
  and (_00002_[6], _00546_, _35583_);
  and (_00002_[5], _00563_, _35583_);
  and (_00002_[4], _00530_, _35583_);
  and (_00002_[3], _00522_, _35583_);
  and (_00002_[2], _00553_, _35583_);
  and (_00002_[1], _00570_, _35583_);
  and (_00002_[0], _00537_, _35583_);
  and (_28437_, _07433_, _03183_);
  and (_28438_, _28437_, _09018_);
  and (_28439_, _03142_, op0_cnst);
  nor (_28440_, _08827_, _02785_);
  and (_28441_, _28440_, _28439_);
  and (_28443_, _02939_, _02895_);
  and (_28444_, _28443_, _28441_);
  and (_28445_, _10388_, _09903_);
  and (_28446_, _28445_, _03188_);
  and (_28447_, _28446_, _28444_);
  and (_28448_, _28447_, _28438_);
  and (_28449_, _28448_, _34446_);
  and (_28450_, _28449_, _35583_);
  nor (_28451_, _27934_, _30854_);
  and (_28452_, _27934_, _30854_);
  or (_28454_, _28452_, _28451_);
  and (_28455_, _10291_, _30810_);
  nor (_28456_, _10291_, _30810_);
  or (_28457_, _28456_, _28455_);
  or (_28458_, _28457_, _28454_);
  and (_28459_, _27806_, _32171_);
  nor (_28460_, _27806_, _32171_);
  and (_28461_, _27535_, _32063_);
  and (_28462_, _27411_, _30830_);
  nor (_28463_, _27535_, _32063_);
  or (_28465_, _28463_, _28462_);
  or (_28466_, _28465_, _28461_);
  and (_28467_, _27669_, _32274_);
  nor (_28468_, _27669_, _32274_);
  or (_28469_, _27293_, _30824_);
  nand (_28470_, _27293_, _30824_);
  and (_28471_, _28470_, _28469_);
  nor (_28472_, _27175_, _30818_);
  and (_28473_, _27175_, _30818_);
  or (_28474_, _28473_, _28472_);
  or (_28476_, _28474_, _28471_);
  nor (_28477_, _27411_, _30830_);
  or (_28478_, _28477_, _28476_);
  or (_28479_, _28478_, _28468_);
  or (_28480_, _28479_, _28467_);
  or (_28481_, _28480_, _28466_);
  or (_28482_, _28481_, _28460_);
  or (_28483_, _28482_, _28459_);
  or (_28484_, _28483_, _28458_);
  and (_00007_, _28484_, _28450_);
  or (_28486_, _10150_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand (_28487_, _10150_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_28488_, _28487_, _28486_);
  nor (_28489_, _26571_, _31231_);
  and (_28490_, _26571_, _31231_);
  or (_28491_, _28490_, _28489_);
  nor (_28492_, _27091_, _30054_);
  and (_28493_, _27091_, _30054_);
  or (_28494_, _28493_, _28492_);
  not (_28495_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_28497_, _26902_, _28495_);
  nor (_28498_, _26902_, _28495_);
  or (_28499_, _28498_, _28497_);
  or (_28500_, _26792_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nand (_28501_, _26792_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_28502_, _28501_, _28500_);
  or (_28503_, _26321_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand (_28504_, _26321_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_28505_, _28504_, _28503_);
  and (_28506_, _26681_, _31267_);
  nor (_28508_, _26681_, _31267_);
  or (_28509_, _28508_, _28506_);
  or (_28510_, _28509_, _28505_);
  or (_28511_, _28510_, _28502_);
  or (_28512_, _28511_, _28499_);
  or (_28513_, _28512_, _28494_);
  or (_28514_, _28513_, _28491_);
  or (_28515_, _28514_, _28488_);
  and (_00006_, _28515_, _28450_);
  or (_00001_, _28448_, rst);
  and (_00005_[7], _00697_, _35583_);
  and (_00004_[7], _00605_, _35583_);
  and (_00003_[7], _00502_, _35583_);
  and (_00002_[7], _00515_, _35583_);
  and (_28517_, _02836_, _31959_);
  nor (_28518_, _02836_, _31959_);
  or (_28519_, _28518_, _28517_);
  not (_28520_, _32239_);
  nor (_28521_, _03742_, _28520_);
  and (_28522_, _03742_, _28520_);
  or (_28524_, _28522_, _28521_);
  or (_28525_, _28524_, _28519_);
  not (_28526_, _32184_);
  nor (_28527_, _03179_, _28526_);
  and (_28528_, _03179_, _28526_);
  or (_28529_, _28528_, _28527_);
  nor (_28530_, _04597_, _32288_);
  and (_28531_, _04597_, _32288_);
  or (_28532_, _28531_, _28530_);
  or (_28533_, _28532_, _28529_);
  or (_28535_, _28533_, _28525_);
  and (_28536_, _02774_, _32079_);
  nor (_28537_, _02774_, _32079_);
  or (_28538_, _28537_, _28536_);
  nand (_28539_, _03320_, _32132_);
  or (_28540_, _03320_, _32132_);
  and (_28541_, _28540_, _28539_);
  or (_28542_, _28541_, _28538_);
  nand (_28543_, _02889_, _32350_);
  or (_28544_, _02889_, _32350_);
  and (_28546_, _28544_, _28543_);
  and (_28547_, _02858_, _32028_);
  nor (_28548_, _02858_, _32028_);
  or (_28549_, _28548_, _28547_);
  or (_28550_, _28549_, _28546_);
  or (_28551_, _28550_, _28542_);
  or (_28552_, _28551_, _28535_);
  nor (_28553_, _09044_, _02598_);
  or (_28554_, _23948_, _02499_);
  and (_28555_, _23793_, _02556_);
  and (_28557_, _09043_, _02548_);
  nor (_28558_, _28557_, _28555_);
  nand (_28559_, _28558_, _02499_);
  and (_28560_, _28559_, _02525_);
  and (_28561_, _28560_, _28554_);
  nor (_28562_, _09044_, _02525_);
  or (_28563_, _28562_, _02476_);
  nor (_28564_, _28563_, _28561_);
  not (_28565_, _28564_);
  and (_28566_, _22129_, \oc8051_golden_model_1.ACC [7]);
  nor (_28568_, _22129_, \oc8051_golden_model_1.ACC [7]);
  nor (_28569_, _28568_, _28566_);
  not (_28570_, _28569_);
  and (_28571_, _21774_, \oc8051_golden_model_1.ACC [6]);
  nor (_28572_, _21774_, \oc8051_golden_model_1.ACC [6]);
  nor (_28573_, _28572_, _28571_);
  and (_28574_, _21401_, \oc8051_golden_model_1.ACC [5]);
  nor (_28575_, _21401_, \oc8051_golden_model_1.ACC [5]);
  and (_28576_, _21041_, \oc8051_golden_model_1.ACC [4]);
  nor (_28577_, _02610_, _02604_);
  nor (_28579_, _28577_, _02609_);
  nor (_28580_, _21041_, \oc8051_golden_model_1.ACC [4]);
  nor (_28581_, _28580_, _28576_);
  not (_28582_, _28581_);
  nor (_28583_, _28582_, _28579_);
  nor (_28584_, _28583_, _28576_);
  nor (_28585_, _28584_, _28575_);
  or (_28586_, _28585_, _28574_);
  and (_28587_, _28586_, _28573_);
  nor (_28588_, _28587_, _28571_);
  nor (_28590_, _28588_, _28570_);
  nor (_28591_, _28590_, _28566_);
  nor (_28592_, _28591_, _22542_);
  and (_28593_, _28592_, \oc8051_golden_model_1.PC [9]);
  and (_28594_, _28593_, _23160_);
  and (_28595_, _28594_, \oc8051_golden_model_1.PC [11]);
  and (_28596_, _28595_, _23793_);
  nor (_28597_, _28595_, _23793_);
  nor (_28598_, _28597_, _28596_);
  nor (_28599_, _28598_, _02552_);
  nor (_28601_, _28599_, _02657_);
  and (_28602_, _28601_, _28565_);
  nor (_28603_, _28602_, _28553_);
  and (_28604_, _34688_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_28605_, _28604_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_28606_, _28605_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_28607_, _28606_, _34683_);
  and (_28608_, _28607_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_28609_, _28608_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_28610_, _28608_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_28612_, _28610_, _28609_);
  nand (_28613_, _28612_, _28603_);
  or (_28614_, _28612_, _28603_);
  nor (_28615_, _09055_, _02598_);
  nor (_28616_, _23329_, _02499_);
  not (_28617_, _02525_);
  and (_28618_, _23161_, _02556_);
  and (_28619_, _09055_, _02548_);
  nor (_28620_, _28619_, _28618_);
  nor (_28621_, _28620_, _07700_);
  nor (_28623_, _28621_, _28617_);
  not (_28624_, _28623_);
  nor (_28625_, _28624_, _28616_);
  nor (_28626_, _09055_, _02525_);
  or (_28627_, _28626_, _02476_);
  nor (_28628_, _28627_, _28625_);
  not (_28629_, _28628_);
  nor (_28630_, _28593_, _23160_);
  nor (_28631_, _28630_, _28594_);
  nor (_28632_, _28631_, _02552_);
  nor (_28634_, _28632_, _02657_);
  and (_28635_, _28634_, _28629_);
  nor (_28636_, _28635_, _28615_);
  and (_28637_, _28606_, _34622_);
  nor (_28638_, _28637_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_28639_, _28638_, _28607_);
  nand (_28640_, _28639_, _28636_);
  or (_28641_, _28639_, _28636_);
  or (_28642_, _28606_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_28643_, _28606_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not (_28644_, _28643_);
  and (_28645_, _28644_, _28642_);
  not (_28646_, _28645_);
  and (_28647_, _22679_, _07700_);
  and (_28648_, _09067_, _02548_);
  and (_28649_, _22495_, _02556_);
  nor (_28650_, _28649_, _28648_);
  nor (_28651_, _28650_, _07700_);
  nor (_28652_, _28651_, _28617_);
  not (_28653_, _28652_);
  nor (_28656_, _28653_, _28647_);
  nor (_28657_, _09067_, _02525_);
  nor (_28658_, _28657_, _02476_);
  not (_28659_, _28658_);
  nor (_28660_, _28659_, _28656_);
  and (_28661_, _28591_, _22542_);
  nor (_28662_, _28661_, _28592_);
  and (_28663_, _28662_, _02476_);
  nor (_28664_, _28663_, _28660_);
  nor (_28665_, _28664_, _02657_);
  nor (_28667_, _09068_, _02598_);
  or (_28668_, _28667_, _28665_);
  nand (_28669_, _28668_, _28646_);
  or (_28670_, _28668_, _28646_);
  nor (_28671_, _28605_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_28672_, _28671_, _28606_);
  and (_28673_, _02598_, _02557_);
  or (_28674_, _05318_, _28673_);
  and (_28675_, _28588_, _28570_);
  nor (_28676_, _28675_, _28590_);
  or (_28678_, _28676_, _02552_);
  and (_28679_, _02525_, _02552_);
  nor (_28680_, _22328_, _02499_);
  and (_28681_, _22138_, _02499_);
  and (_28682_, _28681_, _02556_);
  or (_28683_, _28682_, _28680_);
  nand (_28684_, _28683_, _28679_);
  and (_28685_, _28684_, _28678_);
  or (_28686_, _28685_, _02657_);
  and (_28687_, _28686_, _28674_);
  not (_28689_, _28687_);
  nand (_28690_, _28689_, _28672_);
  or (_28691_, _28689_, _28672_);
  nand (_28692_, _34686_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_28693_, _28692_, _35051_);
  and (_28694_, _28693_, _35055_);
  nor (_28695_, _28693_, _35055_);
  nor (_28696_, _28695_, _28694_);
  nor (_28697_, _28574_, _28575_);
  nor (_28698_, _28697_, _28584_);
  and (_28700_, _28697_, _28584_);
  or (_28701_, _28700_, _28698_);
  or (_28702_, _28701_, _02552_);
  nor (_28703_, _21610_, _02499_);
  and (_28704_, _21415_, _02499_);
  and (_28705_, _28704_, _02556_);
  or (_28706_, _28705_, _28703_);
  nand (_28707_, _28706_, _28679_);
  and (_28708_, _28707_, _28702_);
  or (_28709_, _28708_, _02657_);
  or (_28710_, _09083_, _28673_);
  and (_28711_, _28710_, _28709_);
  or (_28712_, _28711_, _28696_);
  nand (_28713_, _28711_, _28696_);
  and (_28714_, _28713_, _28712_);
  and (_28715_, _34687_, _35055_);
  nor (_28716_, _34687_, _35055_);
  or (_28717_, _28716_, _28715_);
  or (_28718_, _09084_, _03018_);
  nand (_28719_, _21401_, _03018_);
  and (_28721_, _28719_, _28718_);
  or (_28722_, _28721_, _28717_);
  and (_28723_, _08791_, _03018_);
  nor (_28724_, _09138_, _03018_);
  nor (_28725_, _28724_, _28723_);
  or (_28726_, _28725_, _34697_);
  and (_28727_, _23794_, _03018_);
  nor (_28728_, _09043_, _03018_);
  or (_28729_, _28728_, _28727_);
  or (_28730_, _28729_, _35509_);
  and (_28732_, _28730_, _28726_);
  and (_28733_, _28732_, _28722_);
  nor (_28734_, _34686_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  or (_28735_, _28734_, _34687_);
  nor (_28736_, _09089_, _03018_);
  and (_28737_, _21041_, _03018_);
  or (_28738_, _28737_, _28736_);
  or (_28739_, _28738_, _28735_);
  and (_28740_, _24424_, _03018_);
  nor (_28741_, _09030_, _03018_);
  or (_28743_, _28741_, _28740_);
  or (_28744_, _28743_, _35557_);
  and (_28745_, _28744_, _28739_);
  nand (_28746_, _28725_, _34697_);
  or (_28747_, _03021_, _35035_);
  and (_28748_, _28747_, _28746_);
  and (_28749_, _28748_, _28745_);
  and (_28750_, _28749_, _28733_);
  and (_28751_, _28750_, _28714_);
  and (_28752_, _28751_, _28691_);
  and (_28754_, _28752_, _28690_);
  and (_28755_, _28754_, _28670_);
  and (_28756_, _28755_, _28669_);
  and (_28757_, _28756_, _28641_);
  and (_28758_, _28757_, _28640_);
  and (_28759_, _28758_, _28614_);
  and (_28760_, _28759_, _28613_);
  not (_28761_, _34338_);
  nor (_28762_, _03471_, _28761_);
  and (_28763_, _03471_, _28761_);
  or (_28765_, _28763_, _28762_);
  not (_28766_, _34355_);
  nor (_28767_, _03660_, _28766_);
  and (_28768_, _03660_, _28766_);
  or (_28769_, _28768_, _28767_);
  or (_28770_, _28769_, _28765_);
  not (_28771_, _34423_);
  nor (_28772_, _05612_, _28771_);
  and (_28773_, _05612_, _28771_);
  or (_28774_, _28773_, _28772_);
  not (_28776_, _34406_);
  nor (_28777_, _05581_, _28776_);
  and (_28778_, _05581_, _28776_);
  or (_28779_, _28778_, _28777_);
  or (_28780_, _28779_, _28774_);
  or (_28781_, _28780_, _28770_);
  nand (_28782_, _03223_, _34372_);
  or (_28783_, _03223_, _34372_);
  and (_28784_, _28783_, _28782_);
  not (_28785_, _34389_);
  nor (_28787_, _03087_, _28785_);
  and (_28788_, _03087_, _28785_);
  or (_28789_, _28788_, _28787_);
  or (_28790_, _28789_, _28784_);
  nand (_28791_, _05549_, _34440_);
  or (_28792_, _05549_, _34440_);
  and (_28793_, _28792_, _28791_);
  not (_28794_, _34321_);
  nor (_28795_, _05256_, _28794_);
  and (_28796_, _05256_, _28794_);
  or (_28798_, _28796_, _28795_);
  or (_28799_, _28798_, _28793_);
  or (_28800_, _28799_, _28790_);
  or (_28801_, _28800_, _28781_);
  nor (_28802_, _28607_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_28803_, _28802_, _28608_);
  and (_28804_, _23522_, _02556_);
  and (_28805_, _09049_, _02548_);
  nor (_28806_, _28805_, _28804_);
  and (_28807_, _28806_, _02499_);
  and (_28809_, _23639_, _07700_);
  or (_28810_, _28809_, _28807_);
  nor (_28811_, _28810_, _28617_);
  nor (_28812_, _09048_, _02525_);
  nor (_28813_, _28812_, _02476_);
  not (_28814_, _28813_);
  nor (_28815_, _28814_, _28811_);
  nor (_28816_, _28594_, _23478_);
  not (_28817_, _28816_);
  nor (_28818_, _28595_, _02552_);
  and (_28820_, _28818_, _28817_);
  nor (_28821_, _28820_, _28815_);
  nor (_28822_, _28821_, _02657_);
  nor (_28823_, _09049_, _02598_);
  or (_28824_, _28823_, _28822_);
  not (_28825_, _28824_);
  nand (_28826_, _28825_, _28803_);
  or (_28827_, _28825_, _28803_);
  and (_28828_, _22841_, _02556_);
  and (_28829_, _09062_, _02548_);
  nor (_28831_, _28829_, _28828_);
  and (_28832_, _28831_, _02499_);
  and (_28833_, _23010_, _07700_);
  or (_28834_, _28833_, _28832_);
  nor (_28835_, _28834_, _28617_);
  nor (_28836_, _09061_, _02525_);
  nor (_28837_, _28836_, _02476_);
  not (_28838_, _28837_);
  nor (_28839_, _28838_, _28835_);
  nor (_28840_, _28592_, _22831_);
  not (_28842_, _28840_);
  nor (_28843_, _28593_, _02552_);
  and (_28844_, _28843_, _28842_);
  nor (_28845_, _28844_, _28839_);
  nor (_28846_, _28845_, _02657_);
  nor (_28847_, _09062_, _02598_);
  or (_28848_, _28847_, _28846_);
  not (_28849_, _28848_);
  and (_28850_, _28643_, _30879_);
  nor (_28851_, _28643_, _30879_);
  or (_28853_, _28851_, _28850_);
  nand (_28854_, _28853_, _28849_);
  or (_28855_, _28853_, _28849_);
  and (_28856_, _34685_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_28857_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_28858_, _28857_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_28859_, _28858_, _28856_);
  or (_28860_, _28859_, _02603_);
  nor (_28861_, _28604_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_28862_, _28861_, _28605_);
  nor (_28864_, _28586_, _28573_);
  nor (_28865_, _28864_, _28587_);
  and (_28866_, _28865_, _02476_);
  not (_28867_, _28679_);
  and (_28868_, _21969_, _07700_);
  and (_28869_, _21774_, _02499_);
  and (_28870_, _28869_, _02556_);
  nor (_28871_, _28870_, _28868_);
  nor (_28872_, _28871_, _28867_);
  nor (_28873_, _28872_, _28866_);
  nor (_28875_, _28873_, _02657_);
  nor (_28876_, _09077_, _28673_);
  nor (_28877_, _28876_, _28875_);
  nand (_28878_, _28877_, _28862_);
  or (_28879_, _28877_, _28862_);
  and (_28880_, _28879_, _28878_);
  and (_28881_, _28880_, _28860_);
  nand (_28882_, _28859_, _02603_);
  or (_28883_, _02689_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_28884_, _28883_, _28882_);
  and (_28886_, _28884_, _28881_);
  nor (_28887_, \oc8051_golden_model_1.PC [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_28888_, \oc8051_golden_model_1.PC [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_28889_, _28888_, _28887_);
  or (_28890_, _28889_, _03020_);
  or (_28891_, _02441_, _30535_);
  nand (_28892_, _02441_, _30535_);
  and (_28893_, _28892_, _28891_);
  or (_28894_, _02472_, _30437_);
  nand (_28895_, _02472_, _30437_);
  and (_28897_, _28895_, _28894_);
  or (_28898_, _28897_, _28893_);
  or (_28899_, _02496_, _30502_);
  or (_28900_, _02314_, _30503_);
  and (_28901_, _28900_, _28899_);
  or (_28902_, _02527_, _30365_);
  nand (_28903_, _02527_, _30365_);
  and (_28904_, _28903_, _28902_);
  or (_28905_, _28904_, _28901_);
  or (_28906_, _28905_, _28898_);
  nor (_28908_, _02378_, _30459_);
  and (_28909_, _02378_, _30459_);
  or (_28910_, _28909_, _28908_);
  and (_28911_, _02409_, _30482_);
  nor (_28912_, _02409_, _30482_);
  or (_28913_, _28912_, _28911_);
  or (_28914_, _28913_, _28910_);
  and (_28915_, _02801_, _30411_);
  nor (_28916_, _02801_, _30411_);
  or (_28917_, _28916_, _28915_);
  and (_28919_, _02251_, _30389_);
  nor (_28920_, _02251_, _30389_);
  or (_28921_, _28920_, _28919_);
  or (_28922_, _28921_, _28917_);
  or (_28923_, _28922_, _28914_);
  or (_28924_, _28923_, _28906_);
  nor (_28925_, \oc8051_golden_model_1.PC [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_28926_, \oc8051_golden_model_1.PC [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_28927_, _28926_, _28925_);
  nor (_28928_, \oc8051_golden_model_1.PC [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_28930_, \oc8051_golden_model_1.PC [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_28931_, _28930_, _28928_);
  and (_28932_, _28931_, _28927_);
  or (_28933_, \oc8051_golden_model_1.PC [12], _30890_);
  nand (_28934_, \oc8051_golden_model_1.PC [12], _30890_);
  and (_28935_, _28934_, _28933_);
  or (_28936_, \oc8051_golden_model_1.PC [13], _30865_);
  or (_28937_, _24103_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_28938_, _28937_, _28936_);
  and (_28939_, _28938_, _28935_);
  and (_28941_, _28939_, _28932_);
  and (_28942_, \oc8051_golden_model_1.PC [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_28943_, \oc8051_golden_model_1.PC [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_28944_, _28943_, _28942_);
  nor (_28945_, \oc8051_golden_model_1.PC [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_28946_, \oc8051_golden_model_1.PC [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_28947_, _28946_, _28945_);
  and (_28948_, _28947_, _28944_);
  and (_28949_, \oc8051_golden_model_1.PC [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_28950_, \oc8051_golden_model_1.PC [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_28952_, _28950_, _28949_);
  nor (_28953_, \oc8051_golden_model_1.PC [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_28954_, \oc8051_golden_model_1.PC [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_28955_, _28954_, _28953_);
  and (_28956_, _28955_, _28952_);
  and (_28957_, _28956_, _28948_);
  and (_28958_, _28957_, _28941_);
  or (_28959_, \oc8051_golden_model_1.PC [0], _35035_);
  or (_28960_, _02225_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_28961_, _28960_, _28959_);
  nor (_28963_, _28961_, _28889_);
  or (_28964_, \oc8051_golden_model_1.PC [3], _35047_);
  or (_28965_, _02194_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_28966_, _28965_, _28964_);
  and (_28967_, \oc8051_golden_model_1.PC [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_28968_, \oc8051_golden_model_1.PC [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_28969_, _28968_, _28967_);
  and (_28970_, _28969_, _28966_);
  and (_28971_, _28970_, _28963_);
  or (_28972_, \oc8051_golden_model_1.PC [4], _35051_);
  or (_28974_, _21037_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_28975_, _28974_, _28972_);
  nand (_28976_, \oc8051_golden_model_1.PC [5], _35055_);
  or (_28977_, \oc8051_golden_model_1.PC [5], _35055_);
  and (_28978_, _28977_, _28976_);
  and (_28979_, _28978_, _28975_);
  or (_28980_, \oc8051_golden_model_1.PC [6], _35059_);
  nand (_28981_, \oc8051_golden_model_1.PC [6], _35059_);
  and (_28982_, _28981_, _28980_);
  and (_28983_, \oc8051_golden_model_1.PC [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_28985_, \oc8051_golden_model_1.PC [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  or (_28986_, _28985_, _28983_);
  and (_28987_, _28986_, _28982_);
  and (_28988_, _28987_, _28979_);
  and (_28989_, _28988_, _28971_);
  and (_28990_, _28989_, _28958_);
  and (_28991_, _28990_, _34446_);
  and (_28992_, _28991_, _28924_);
  and (_28993_, _28992_, _28890_);
  and (_28994_, _24109_, _03018_);
  nor (_28996_, _09038_, _03018_);
  nor (_28997_, _28996_, _28994_);
  nand (_28998_, _28997_, _35536_);
  or (_28999_, _28997_, _35536_);
  and (_29000_, _28999_, _28998_);
  nor (_29001_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_29002_, _29001_, _34685_);
  nand (_29003_, _29002_, _03029_);
  or (_29004_, _29002_, _03029_);
  and (_29005_, _29004_, _29003_);
  and (_29007_, _29005_, _29000_);
  and (_29008_, _28692_, _35051_);
  nor (_29009_, _29008_, _28693_);
  and (_29010_, _28582_, _28579_);
  nor (_29011_, _29010_, _28583_);
  or (_29012_, _29011_, _02552_);
  nor (_29013_, _21243_, _02499_);
  and (_29014_, _21042_, _02499_);
  and (_29015_, _29014_, _02556_);
  or (_29016_, _29015_, _29013_);
  nand (_29018_, _29016_, _28679_);
  and (_29019_, _29018_, _29012_);
  or (_29020_, _29019_, _02657_);
  or (_29021_, _09088_, _28673_);
  and (_29022_, _29021_, _29020_);
  not (_29023_, _29022_);
  nand (_29024_, _29023_, _29009_);
  nor (_29025_, _34685_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_29026_, _29025_, _34686_);
  or (_29027_, _29026_, _03032_);
  nand (_29029_, _29026_, _03032_);
  and (_29030_, _29029_, _29027_);
  and (_29031_, _29030_, _29024_);
  and (_29032_, _29031_, _29007_);
  and (_29033_, _23478_, _03018_);
  nor (_29034_, _09049_, _03018_);
  nor (_29035_, _29034_, _29033_);
  nand (_29036_, _29035_, _35477_);
  or (_29037_, _29035_, _35477_);
  and (_29038_, _29037_, _29036_);
  and (_29040_, _28856_, _35047_);
  nor (_29041_, _28856_, _35047_);
  nor (_29042_, _29041_, _29040_);
  or (_29043_, _29042_, _02696_);
  and (_29044_, _29043_, _29038_);
  or (_29045_, _29023_, _29009_);
  nand (_29046_, _29042_, _02696_);
  and (_29047_, _29046_, _29045_);
  and (_29048_, _29047_, _29044_);
  and (_29049_, _29048_, _29032_);
  and (_29051_, _29049_, _28993_);
  and (_29052_, _29051_, _28886_);
  and (_29053_, _02685_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_29054_, _02700_, _35039_);
  nor (_29055_, _29054_, _29053_);
  nand (_29056_, _29055_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_29057_, _29055_, _02666_);
  and (_29058_, _29057_, _29056_);
  and (_29059_, _29058_, _29052_);
  and (_29060_, _29059_, _28855_);
  and (_29062_, _29060_, _28854_);
  and (_29063_, _29062_, _28827_);
  and (_29064_, _29063_, _28826_);
  and (_29065_, _29064_, _28801_);
  and (_29066_, _29065_, _28760_);
  and (property_invalid_rom_pc, _29066_, _28552_);
  nor (_29067_, _30854_, \oc8051_golden_model_1.SP [6]);
  and (_29068_, _30854_, \oc8051_golden_model_1.SP [6]);
  or (_29069_, _29068_, _29067_);
  nor (_29070_, _30810_, _10154_);
  and (_29072_, _30810_, _10154_);
  or (_29073_, _29072_, _29070_);
  or (_29074_, _29073_, _29069_);
  nor (_29075_, _30848_, \oc8051_golden_model_1.SP [5]);
  and (_29076_, _30848_, \oc8051_golden_model_1.SP [5]);
  or (_29077_, _29076_, _29075_);
  and (_29078_, _30836_, \oc8051_golden_model_1.SP [3]);
  nor (_29079_, _30836_, \oc8051_golden_model_1.SP [3]);
  or (_29080_, _29079_, _29078_);
  and (_29081_, _30830_, \oc8051_golden_model_1.SP [2]);
  or (_29083_, _30818_, _02787_);
  nand (_29084_, _30818_, _02787_);
  and (_29085_, _29084_, _29083_);
  and (_29086_, _30824_, \oc8051_golden_model_1.SP [1]);
  nor (_29087_, _30824_, \oc8051_golden_model_1.SP [1]);
  or (_29088_, _29087_, _29086_);
  or (_29089_, _29088_, _29085_);
  nor (_29090_, _30830_, \oc8051_golden_model_1.SP [2]);
  or (_29091_, _29090_, _29089_);
  or (_29092_, _29091_, _29081_);
  or (_29094_, _29092_, _29080_);
  and (_29095_, _30842_, \oc8051_golden_model_1.SP [4]);
  nor (_29096_, _30842_, \oc8051_golden_model_1.SP [4]);
  or (_29097_, _29096_, _29095_);
  or (_29098_, _29097_, _29094_);
  or (_29099_, _29098_, _29077_);
  or (_29100_, _29099_, _29074_);
  and (_29101_, _28448_, inst_finished_r);
  and (_29102_, _29101_, property_invalid_sp_1_r);
  and (property_invalid_sp, _29102_, _29100_);
  and (_29104_, _26685_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_29105_, \oc8051_golden_model_1.PSW [4], _31281_);
  or (_29106_, _29105_, _29104_);
  and (_29107_, _02937_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_29108_, \oc8051_golden_model_1.PSW [3], _31267_);
  or (_29109_, _29108_, _29107_);
  or (_29110_, _29109_, _29106_);
  and (_29111_, _26221_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_29112_, \oc8051_golden_model_1.PSW [1], _31223_);
  or (_29113_, _29112_, _29111_);
  nand (_29115_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_29116_, \oc8051_golden_model_1.PSW [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_29117_, _29116_, _29115_);
  or (_29118_, _29117_, _29113_);
  or (_29119_, _29118_, _29110_);
  and (_29120_, _07294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_29121_, \oc8051_golden_model_1.PSW [7], _31206_);
  or (_29122_, _29121_, _29120_);
  and (_29123_, _26797_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_29124_, \oc8051_golden_model_1.PSW [5], _28495_);
  or (_29126_, _29124_, _29123_);
  nand (_29127_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_29128_, \oc8051_golden_model_1.PSW [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_29129_, _29128_, _29127_);
  or (_29130_, _29129_, _29126_);
  or (_29131_, _29130_, _29122_);
  or (_29132_, _29131_, _29119_);
  and (_29133_, _29132_, property_invalid_psw_1_r);
  and (property_invalid_psw, _29133_, _29101_);
  nand (_29134_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_29136_, \oc8051_golden_model_1.P3 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_29137_, _29136_, _29134_);
  and (_29138_, _19091_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_29139_, \oc8051_golden_model_1.P3 [2], _31790_);
  or (_29140_, _29139_, _29138_);
  or (_29141_, _29140_, _29137_);
  and (_29142_, \oc8051_golden_model_1.P3 [0], _31764_);
  and (_29143_, _18877_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_29144_, _29143_, _29142_);
  and (_29145_, _18981_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_29147_, \oc8051_golden_model_1.P3 [1], _31777_);
  or (_29148_, _29147_, _29145_);
  or (_29149_, _29148_, _29144_);
  or (_29150_, _29149_, _29141_);
  or (_29151_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand (_29152_, \oc8051_golden_model_1.P3 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_29153_, _29152_, _29151_);
  or (_29154_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand (_29155_, \oc8051_golden_model_1.P3 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_29156_, _29155_, _29154_);
  or (_29158_, _29156_, _29153_);
  and (_29159_, _08672_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_29160_, \oc8051_golden_model_1.P3 [7], _31482_);
  or (_29161_, _29160_, _29159_);
  nand (_29162_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_29163_, \oc8051_golden_model_1.P3 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_29164_, _29163_, _29162_);
  or (_29165_, _29164_, _29161_);
  or (_29166_, _29165_, _29158_);
  or (_29167_, _29166_, _29150_);
  and (property_invalid_p3, _29167_, _29101_);
  nand (_29169_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_29170_, \oc8051_golden_model_1.P2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_29171_, _29170_, _29169_);
  and (_29172_, _18334_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_29173_, \oc8051_golden_model_1.P2 [2], _31702_);
  or (_29174_, _29173_, _29172_);
  or (_29175_, _29174_, _29171_);
  and (_29176_, \oc8051_golden_model_1.P2 [0], _31676_);
  and (_29177_, _18121_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_29179_, _29177_, _29176_);
  and (_29180_, _18224_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_29181_, \oc8051_golden_model_1.P2 [1], _31689_);
  or (_29182_, _29181_, _29180_);
  or (_29183_, _29182_, _29179_);
  or (_29184_, _29183_, _29175_);
  or (_29185_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nand (_29186_, \oc8051_golden_model_1.P2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_29187_, _29186_, _29185_);
  or (_29188_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nand (_29189_, \oc8051_golden_model_1.P2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_29190_, _29189_, _29188_);
  or (_29191_, _29190_, _29187_);
  and (_29192_, _08572_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_29193_, \oc8051_golden_model_1.P2 [7], _31466_);
  or (_29194_, _29193_, _29192_);
  nand (_29195_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_29196_, \oc8051_golden_model_1.P2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_29197_, _29196_, _29195_);
  or (_29198_, _29197_, _29194_);
  or (_29201_, _29198_, _29191_);
  or (_29202_, _29201_, _29184_);
  and (property_invalid_p2, _29202_, _29101_);
  nand (_29203_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_29204_, \oc8051_golden_model_1.P1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_29205_, _29204_, _29203_);
  and (_29206_, _17578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_29207_, \oc8051_golden_model_1.P1 [2], _31614_);
  or (_29208_, _29207_, _29206_);
  or (_29209_, _29208_, _29205_);
  and (_29211_, \oc8051_golden_model_1.P1 [0], _31588_);
  and (_29212_, _17364_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_29213_, _29212_, _29211_);
  and (_29214_, _17468_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_29215_, \oc8051_golden_model_1.P1 [1], _31601_);
  or (_29216_, _29215_, _29214_);
  or (_29217_, _29216_, _29213_);
  or (_29218_, _29217_, _29209_);
  or (_29219_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nand (_29220_, \oc8051_golden_model_1.P1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_29222_, _29220_, _29219_);
  or (_29223_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nand (_29224_, \oc8051_golden_model_1.P1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_29225_, _29224_, _29223_);
  or (_29226_, _29225_, _29222_);
  and (_29227_, _08472_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_29228_, \oc8051_golden_model_1.P1 [7], _31447_);
  or (_29229_, _29228_, _29227_);
  nand (_29230_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_29231_, \oc8051_golden_model_1.P1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_29233_, _29231_, _29230_);
  or (_29234_, _29233_, _29229_);
  or (_29235_, _29234_, _29226_);
  or (_29236_, _29235_, _29218_);
  and (property_invalid_p1, _29236_, _29101_);
  nand (_29237_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_29238_, \oc8051_golden_model_1.P0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_29239_, _29238_, _29237_);
  and (_29240_, _16814_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_29241_, \oc8051_golden_model_1.P0 [2], _31525_);
  or (_29243_, _29241_, _29240_);
  or (_29244_, _29243_, _29239_);
  and (_29245_, \oc8051_golden_model_1.P0 [0], _31489_);
  and (_29246_, _16598_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_29247_, _29246_, _29245_);
  and (_29248_, _16703_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_29249_, \oc8051_golden_model_1.P0 [1], _31509_);
  or (_29250_, _29249_, _29248_);
  or (_29251_, _29250_, _29247_);
  or (_29252_, _29251_, _29244_);
  or (_29254_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand (_29255_, \oc8051_golden_model_1.P0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_29256_, _29255_, _29254_);
  or (_29257_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nand (_29258_, \oc8051_golden_model_1.P0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_29259_, _29258_, _29257_);
  or (_29260_, _29259_, _29256_);
  and (_29261_, _08371_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_29262_, \oc8051_golden_model_1.P0 [7], _31434_);
  or (_29263_, _29262_, _29261_);
  nand (_29265_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_29266_, \oc8051_golden_model_1.P0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_29267_, _29266_, _29265_);
  or (_29268_, _29267_, _29263_);
  or (_29269_, _29268_, _29260_);
  or (_29270_, _29269_, _29252_);
  and (property_invalid_p0, _29270_, _29101_);
  or (_29271_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_29272_, \oc8051_golden_model_1.IRAM[0] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  and (_29273_, _29272_, _29271_);
  nand (_29275_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or (_29276_, \oc8051_golden_model_1.IRAM[0] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  and (_29277_, _29276_, _29275_);
  or (_29278_, _29277_, _29273_);
  and (_29279_, \oc8051_golden_model_1.IRAM[0] [0], _32442_);
  and (_29280_, _03338_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or (_29281_, _29280_, _29279_);
  and (_29282_, _03933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  and (_29283_, \oc8051_golden_model_1.IRAM[0] [1], _32446_);
  or (_29284_, _29283_, _29282_);
  or (_29286_, _29284_, _29281_);
  or (_29287_, _29286_, _29278_);
  or (_29288_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nand (_29289_, \oc8051_golden_model_1.IRAM[0] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  and (_29290_, _29289_, _29288_);
  nand (_29291_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or (_29292_, \oc8051_golden_model_1.IRAM[0] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  and (_29293_, _29292_, _29291_);
  or (_29294_, _29293_, _29290_);
  or (_29295_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand (_29297_, \oc8051_golden_model_1.IRAM[0] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  and (_29298_, _29297_, _29295_);
  or (_29299_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand (_29300_, \oc8051_golden_model_1.IRAM[0] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  and (_29301_, _29300_, _29299_);
  or (_29302_, _29301_, _29298_);
  or (_29303_, _29302_, _29294_);
  or (_29304_, _29303_, _29287_);
  or (_29305_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_29306_, \oc8051_golden_model_1.IRAM[1] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  and (_29308_, _29306_, _29305_);
  or (_29309_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_29310_, \oc8051_golden_model_1.IRAM[1] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  and (_29311_, _29310_, _29309_);
  or (_29312_, _29311_, _29308_);
  or (_29313_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nand (_29314_, \oc8051_golden_model_1.IRAM[1] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  and (_29315_, _29314_, _29313_);
  nand (_29316_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  or (_29317_, \oc8051_golden_model_1.IRAM[1] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  and (_29319_, _29317_, _29316_);
  or (_29320_, _29319_, _29315_);
  or (_29321_, _29320_, _29312_);
  and (_29322_, _04786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  and (_29323_, \oc8051_golden_model_1.IRAM[1] [5], _32482_);
  or (_29324_, _29323_, _29322_);
  and (_29325_, _05090_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  and (_29326_, \oc8051_golden_model_1.IRAM[1] [4], _32479_);
  or (_29327_, _29326_, _29325_);
  or (_29328_, _29327_, _29324_);
  or (_29330_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nand (_29331_, \oc8051_golden_model_1.IRAM[1] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  and (_29332_, _29331_, _29330_);
  nand (_29333_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  or (_29334_, \oc8051_golden_model_1.IRAM[1] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  and (_29335_, _29334_, _29333_);
  or (_29336_, _29335_, _29332_);
  or (_29337_, _29336_, _29328_);
  or (_29338_, _29337_, _29321_);
  or (_29339_, _29338_, _29304_);
  or (_29341_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nand (_29342_, \oc8051_golden_model_1.IRAM[2] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and (_29343_, _29342_, _29341_);
  or (_29344_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nand (_29345_, \oc8051_golden_model_1.IRAM[2] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  and (_29346_, _29345_, _29344_);
  or (_29347_, _29346_, _29343_);
  and (_29348_, _04365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  and (_29349_, \oc8051_golden_model_1.IRAM[2] [2], _32497_);
  or (_29350_, _29349_, _29348_);
  nand (_29352_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or (_29353_, \oc8051_golden_model_1.IRAM[2] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  and (_29354_, _29353_, _29352_);
  or (_29355_, _29354_, _29350_);
  or (_29356_, _29355_, _29347_);
  and (_29357_, _05095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and (_29358_, \oc8051_golden_model_1.IRAM[2] [4], _32502_);
  or (_29359_, _29358_, _29357_);
  and (_29360_, _04791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and (_29361_, \oc8051_golden_model_1.IRAM[2] [5], _32505_);
  or (_29363_, _29361_, _29360_);
  or (_29364_, _29363_, _29359_);
  and (_29365_, \oc8051_golden_model_1.IRAM[2] [7], _32510_);
  and (_29366_, _04537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or (_29367_, _29366_, _29365_);
  nand (_29368_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or (_29369_, \oc8051_golden_model_1.IRAM[2] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  and (_29370_, _29369_, _29368_);
  or (_29371_, _29370_, _29367_);
  or (_29372_, _29371_, _29364_);
  or (_29374_, _29372_, _29356_);
  and (_29375_, \oc8051_golden_model_1.IRAM[3] [2], _32520_);
  and (_29376_, _04363_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  or (_29377_, _29376_, _29375_);
  nand (_29378_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  or (_29379_, \oc8051_golden_model_1.IRAM[3] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  and (_29380_, _29379_, _29378_);
  or (_29381_, _29380_, _29377_);
  and (_29382_, _03752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  and (_29383_, \oc8051_golden_model_1.IRAM[3] [0], _32514_);
  or (_29385_, _29383_, _29382_);
  and (_29386_, \oc8051_golden_model_1.IRAM[3] [1], _32517_);
  and (_29387_, _03938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  or (_29388_, _29387_, _29386_);
  or (_29389_, _29388_, _29385_);
  or (_29390_, _29389_, _29381_);
  and (_29391_, _04535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  and (_29392_, \oc8051_golden_model_1.IRAM[3] [7], _32375_);
  or (_29393_, _29392_, _29391_);
  nand (_29394_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  or (_29396_, \oc8051_golden_model_1.IRAM[3] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and (_29397_, _29396_, _29394_);
  or (_29398_, _29397_, _29393_);
  or (_29399_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_29400_, \oc8051_golden_model_1.IRAM[3] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  and (_29401_, _29400_, _29399_);
  or (_29402_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_29403_, \oc8051_golden_model_1.IRAM[3] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  and (_29404_, _29403_, _29402_);
  or (_29405_, _29404_, _29401_);
  or (_29407_, _29405_, _29398_);
  or (_29408_, _29407_, _29390_);
  or (_29409_, _29408_, _29374_);
  or (_29410_, _29409_, _29339_);
  and (_29411_, _03768_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and (_29412_, \oc8051_golden_model_1.IRAM[4] [0], _32538_);
  or (_29413_, _29412_, _29411_);
  and (_29414_, \oc8051_golden_model_1.IRAM[4] [1], _32541_);
  and (_29415_, _03951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or (_29416_, _29415_, _29414_);
  or (_29417_, _29416_, _29413_);
  or (_29418_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nand (_29419_, \oc8051_golden_model_1.IRAM[4] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  and (_29420_, _29419_, _29418_);
  nand (_29421_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or (_29422_, \oc8051_golden_model_1.IRAM[4] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and (_29423_, _29422_, _29421_);
  or (_29424_, _29423_, _29420_);
  or (_29425_, _29424_, _29417_);
  or (_29426_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nand (_29428_, \oc8051_golden_model_1.IRAM[4] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  and (_29429_, _29428_, _29426_);
  or (_29430_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nand (_29431_, \oc8051_golden_model_1.IRAM[4] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  and (_29432_, _29431_, _29430_);
  or (_29433_, _29432_, _29429_);
  or (_29434_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nand (_29435_, \oc8051_golden_model_1.IRAM[4] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  and (_29436_, _29435_, _29434_);
  nand (_29437_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or (_29439_, \oc8051_golden_model_1.IRAM[4] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  and (_29440_, _29439_, _29437_);
  or (_29441_, _29440_, _29436_);
  or (_29442_, _29441_, _29433_);
  or (_29443_, _29442_, _29425_);
  or (_29444_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nand (_29445_, \oc8051_golden_model_1.IRAM[5] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  and (_29446_, _29445_, _29444_);
  nand (_29447_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  or (_29448_, \oc8051_golden_model_1.IRAM[5] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  and (_29449_, _29448_, _29447_);
  or (_29450_, _29449_, _29446_);
  or (_29451_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_29452_, \oc8051_golden_model_1.IRAM[5] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  and (_29453_, _29452_, _29451_);
  or (_29454_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_29455_, \oc8051_golden_model_1.IRAM[5] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  and (_29456_, _29455_, _29454_);
  or (_29457_, _29456_, _29453_);
  or (_29458_, _29457_, _29450_);
  or (_29461_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nand (_29462_, \oc8051_golden_model_1.IRAM[5] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and (_29463_, _29462_, _29461_);
  nand (_29464_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  or (_29465_, \oc8051_golden_model_1.IRAM[5] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and (_29466_, _29465_, _29464_);
  or (_29467_, _29466_, _29463_);
  and (_29468_, _05109_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and (_29469_, \oc8051_golden_model_1.IRAM[5] [4], _32568_);
  or (_29470_, _29469_, _29468_);
  and (_29472_, _04805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and (_29473_, \oc8051_golden_model_1.IRAM[5] [5], _32571_);
  or (_29474_, _29473_, _29472_);
  or (_29475_, _29474_, _29470_);
  or (_29476_, _29475_, _29467_);
  or (_29477_, _29476_, _29458_);
  or (_29478_, _29477_, _29443_);
  and (_29479_, \oc8051_golden_model_1.IRAM[6] [2], _32585_);
  and (_29480_, _04373_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or (_29481_, _29480_, _29479_);
  nand (_29483_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or (_29484_, \oc8051_golden_model_1.IRAM[6] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and (_29485_, _29484_, _29483_);
  or (_29486_, _29485_, _29481_);
  or (_29487_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nand (_29488_, \oc8051_golden_model_1.IRAM[6] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and (_29489_, _29488_, _29487_);
  or (_29490_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nand (_29491_, \oc8051_golden_model_1.IRAM[6] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  and (_29492_, _29491_, _29490_);
  or (_29494_, _29492_, _29489_);
  or (_29495_, _29494_, _29486_);
  and (_29496_, _04545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  and (_29497_, \oc8051_golden_model_1.IRAM[6] [7], _32598_);
  or (_29498_, _29497_, _29496_);
  nand (_29499_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or (_29500_, \oc8051_golden_model_1.IRAM[6] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and (_29501_, _29500_, _29499_);
  or (_29502_, _29501_, _29498_);
  and (_29503_, _05103_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and (_29505_, \oc8051_golden_model_1.IRAM[6] [4], _32590_);
  or (_29506_, _29505_, _29503_);
  and (_29507_, \oc8051_golden_model_1.IRAM[6] [5], _32593_);
  and (_29508_, _04799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or (_29509_, _29508_, _29507_);
  or (_29510_, _29509_, _29506_);
  or (_29511_, _29510_, _29502_);
  or (_29512_, _29511_, _29495_);
  and (_29513_, _03945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and (_29514_, \oc8051_golden_model_1.IRAM[7] [1], _32605_);
  or (_29516_, _29514_, _29513_);
  and (_29517_, _03762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and (_29518_, \oc8051_golden_model_1.IRAM[7] [0], _32602_);
  or (_29519_, _29518_, _29517_);
  or (_29520_, _29519_, _29516_);
  and (_29521_, _04371_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  and (_29522_, \oc8051_golden_model_1.IRAM[7] [2], _32608_);
  or (_29523_, _29522_, _29521_);
  nand (_29524_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  or (_29525_, \oc8051_golden_model_1.IRAM[7] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and (_29527_, _29525_, _29524_);
  or (_29528_, _29527_, _29523_);
  or (_29529_, _29528_, _29520_);
  or (_29530_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_29531_, \oc8051_golden_model_1.IRAM[7] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and (_29532_, _29531_, _29530_);
  or (_29533_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_29534_, \oc8051_golden_model_1.IRAM[7] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and (_29535_, _29534_, _29533_);
  or (_29536_, _29535_, _29532_);
  and (_29538_, _04543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and (_29539_, \oc8051_golden_model_1.IRAM[7] [7], _32387_);
  or (_29540_, _29539_, _29538_);
  nand (_29541_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  or (_29542_, \oc8051_golden_model_1.IRAM[7] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and (_29543_, _29542_, _29541_);
  or (_29544_, _29543_, _29540_);
  or (_29545_, _29544_, _29536_);
  or (_29546_, _29545_, _29529_);
  or (_29547_, _29546_, _29512_);
  or (_29549_, _29547_, _29478_);
  or (_29550_, _29549_, _29410_);
  and (_29551_, _03784_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  and (_29552_, \oc8051_golden_model_1.IRAM[8] [0], _32626_);
  or (_29553_, _29552_, _29551_);
  and (_29554_, \oc8051_golden_model_1.IRAM[8] [1], _32629_);
  and (_29555_, _03966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  or (_29556_, _29555_, _29554_);
  or (_29557_, _29556_, _29553_);
  or (_29558_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nand (_29560_, \oc8051_golden_model_1.IRAM[8] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  and (_29561_, _29560_, _29558_);
  or (_29562_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nand (_29563_, \oc8051_golden_model_1.IRAM[8] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  and (_29564_, _29563_, _29562_);
  or (_29565_, _29564_, _29561_);
  or (_29566_, _29565_, _29557_);
  or (_29567_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nand (_29568_, \oc8051_golden_model_1.IRAM[8] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  and (_29569_, _29568_, _29567_);
  or (_29571_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nand (_29572_, \oc8051_golden_model_1.IRAM[8] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  and (_29573_, _29572_, _29571_);
  or (_29574_, _29573_, _29569_);
  or (_29575_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nand (_29576_, \oc8051_golden_model_1.IRAM[8] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  and (_29577_, _29576_, _29575_);
  or (_29578_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_29579_, \oc8051_golden_model_1.IRAM[8] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and (_29580_, _29579_, _29578_);
  or (_29582_, _29580_, _29577_);
  or (_29583_, _29582_, _29574_);
  or (_29584_, _29583_, _29566_);
  or (_29585_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nand (_29586_, \oc8051_golden_model_1.IRAM[9] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and (_29587_, _29586_, _29585_);
  nand (_29588_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  or (_29589_, \oc8051_golden_model_1.IRAM[9] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and (_29590_, _29589_, _29588_);
  or (_29591_, _29590_, _29587_);
  or (_29593_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nand (_29594_, \oc8051_golden_model_1.IRAM[9] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and (_29595_, _29594_, _29593_);
  or (_29596_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nand (_29597_, \oc8051_golden_model_1.IRAM[9] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and (_29598_, _29597_, _29596_);
  or (_29599_, _29598_, _29595_);
  or (_29600_, _29599_, _29591_);
  and (_29601_, _04819_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and (_29602_, \oc8051_golden_model_1.IRAM[9] [5], _32658_);
  or (_29604_, _29602_, _29601_);
  and (_29605_, _05123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  and (_29606_, \oc8051_golden_model_1.IRAM[9] [4], _32655_);
  or (_29607_, _29606_, _29605_);
  or (_29608_, _29607_, _29604_);
  or (_29609_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nand (_29610_, \oc8051_golden_model_1.IRAM[9] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and (_29611_, _29610_, _29609_);
  nand (_29612_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  or (_29613_, \oc8051_golden_model_1.IRAM[9] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and (_29615_, _29613_, _29612_);
  or (_29616_, _29615_, _29611_);
  or (_29617_, _29616_, _29608_);
  or (_29618_, _29617_, _29600_);
  or (_29619_, _29618_, _29584_);
  nand (_29620_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  or (_29621_, \oc8051_golden_model_1.IRAM[10] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and (_29622_, _29621_, _29620_);
  and (_29623_, _04389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and (_29624_, \oc8051_golden_model_1.IRAM[10] [2], _32671_);
  or (_29626_, _29624_, _29623_);
  or (_29627_, _29626_, _29622_);
  or (_29628_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nand (_29629_, \oc8051_golden_model_1.IRAM[10] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and (_29630_, _29629_, _29628_);
  or (_29631_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nand (_29632_, \oc8051_golden_model_1.IRAM[10] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and (_29633_, _29632_, _29631_);
  or (_29634_, _29633_, _29630_);
  or (_29635_, _29634_, _29627_);
  and (_29637_, \oc8051_golden_model_1.IRAM[10] [7], _32401_);
  and (_29638_, _04561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  or (_29639_, _29638_, _29637_);
  nand (_29640_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  or (_29641_, \oc8051_golden_model_1.IRAM[10] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and (_29642_, _29641_, _29640_);
  or (_29643_, _29642_, _29639_);
  and (_29644_, _05118_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and (_29645_, \oc8051_golden_model_1.IRAM[10] [4], _32676_);
  or (_29646_, _29645_, _29644_);
  and (_29648_, \oc8051_golden_model_1.IRAM[10] [5], _32679_);
  and (_29649_, _04814_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  or (_29650_, _29649_, _29648_);
  or (_29651_, _29650_, _29646_);
  or (_29652_, _29651_, _29643_);
  or (_29653_, _29652_, _29635_);
  and (_29654_, _03779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and (_29655_, \oc8051_golden_model_1.IRAM[11] [0], _32688_);
  or (_29656_, _29655_, _29654_);
  and (_29657_, \oc8051_golden_model_1.IRAM[11] [1], _32691_);
  and (_29659_, _03961_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  or (_29660_, _29659_, _29657_);
  or (_29661_, _29660_, _29656_);
  and (_29662_, \oc8051_golden_model_1.IRAM[11] [2], _32694_);
  and (_29663_, _04387_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  or (_29664_, _29663_, _29662_);
  nand (_29665_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  or (_29666_, \oc8051_golden_model_1.IRAM[11] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and (_29667_, _29666_, _29665_);
  or (_29668_, _29667_, _29664_);
  or (_29670_, _29668_, _29661_);
  or (_29671_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nand (_29672_, \oc8051_golden_model_1.IRAM[11] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and (_29673_, _29672_, _29671_);
  or (_29674_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand (_29675_, \oc8051_golden_model_1.IRAM[11] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  and (_29676_, _29675_, _29674_);
  or (_29677_, _29676_, _29673_);
  and (_29678_, _04559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and (_29679_, \oc8051_golden_model_1.IRAM[11] [7], _32707_);
  or (_29681_, _29679_, _29678_);
  or (_29682_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand (_29683_, \oc8051_golden_model_1.IRAM[11] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  and (_29684_, _29683_, _29682_);
  or (_29685_, _29684_, _29681_);
  or (_29686_, _29685_, _29677_);
  or (_29687_, _29686_, _29670_);
  or (_29688_, _29687_, _29653_);
  or (_29689_, _29688_, _29619_);
  or (_29690_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nand (_29692_, \oc8051_golden_model_1.IRAM[12] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and (_29693_, _29692_, _29690_);
  or (_29694_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nand (_29695_, \oc8051_golden_model_1.IRAM[12] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and (_29696_, _29695_, _29694_);
  or (_29697_, _29696_, _29693_);
  and (_29698_, \oc8051_golden_model_1.IRAM[12] [1], _32714_);
  and (_29699_, _03979_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  or (_29700_, _29699_, _29698_);
  and (_29701_, _03796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  and (_29703_, \oc8051_golden_model_1.IRAM[12] [0], _32711_);
  or (_29704_, _29703_, _29701_);
  or (_29705_, _29704_, _29700_);
  or (_29706_, _29705_, _29697_);
  or (_29707_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_29708_, \oc8051_golden_model_1.IRAM[12] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and (_29709_, _29708_, _29707_);
  or (_29710_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nand (_29711_, \oc8051_golden_model_1.IRAM[12] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  and (_29712_, _29711_, _29710_);
  or (_29714_, _29712_, _29709_);
  or (_29715_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nand (_29716_, \oc8051_golden_model_1.IRAM[12] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  and (_29717_, _29716_, _29715_);
  or (_29718_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nand (_29719_, \oc8051_golden_model_1.IRAM[12] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  and (_29720_, _29719_, _29718_);
  or (_29721_, _29720_, _29717_);
  or (_29722_, _29721_, _29714_);
  or (_29723_, _29722_, _29706_);
  or (_29725_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nand (_29726_, \oc8051_golden_model_1.IRAM[13] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and (_29727_, _29726_, _29725_);
  or (_29728_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nand (_29729_, \oc8051_golden_model_1.IRAM[13] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and (_29730_, _29729_, _29728_);
  or (_29731_, _29730_, _29727_);
  or (_29732_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nand (_29733_, \oc8051_golden_model_1.IRAM[13] [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and (_29734_, _29733_, _29732_);
  nand (_29736_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  or (_29737_, \oc8051_golden_model_1.IRAM[13] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and (_29738_, _29737_, _29736_);
  or (_29739_, _29738_, _29734_);
  or (_29740_, _29739_, _29731_);
  and (_29741_, _05135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and (_29742_, \oc8051_golden_model_1.IRAM[13] [4], _32741_);
  or (_29743_, _29742_, _29741_);
  and (_29744_, \oc8051_golden_model_1.IRAM[13] [5], _32744_);
  and (_29745_, _04831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  or (_29747_, _29745_, _29744_);
  or (_29748_, _29747_, _29743_);
  or (_29749_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nand (_29750_, \oc8051_golden_model_1.IRAM[13] [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and (_29751_, _29750_, _29749_);
  nand (_29752_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  or (_29753_, \oc8051_golden_model_1.IRAM[13] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and (_29754_, _29753_, _29752_);
  or (_29755_, _29754_, _29751_);
  or (_29756_, _29755_, _29748_);
  or (_29757_, _29756_, _29740_);
  or (_29758_, _29757_, _29723_);
  or (_29759_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nand (_29760_, \oc8051_golden_model_1.IRAM[14] [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and (_29761_, _29760_, _29759_);
  or (_29762_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nand (_29763_, \oc8051_golden_model_1.IRAM[14] [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  and (_29764_, _29763_, _29762_);
  or (_29765_, _29764_, _29761_);
  and (_29766_, \oc8051_golden_model_1.IRAM[14] [2], _32758_);
  and (_29769_, _04401_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  or (_29770_, _29769_, _29766_);
  nand (_29771_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  or (_29772_, \oc8051_golden_model_1.IRAM[14] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and (_29773_, _29772_, _29771_);
  or (_29774_, _29773_, _29770_);
  or (_29775_, _29774_, _29765_);
  and (_29776_, \oc8051_golden_model_1.IRAM[14] [5], _32766_);
  and (_29777_, _04826_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  or (_29778_, _29777_, _29776_);
  and (_29780_, _05130_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  and (_29781_, \oc8051_golden_model_1.IRAM[14] [4], _32763_);
  or (_29782_, _29781_, _29780_);
  or (_29783_, _29782_, _29778_);
  and (_29784_, _04573_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and (_29785_, \oc8051_golden_model_1.IRAM[14] [7], _32412_);
  or (_29786_, _29785_, _29784_);
  nand (_29787_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  or (_29788_, \oc8051_golden_model_1.IRAM[14] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and (_29789_, _29788_, _29787_);
  or (_29791_, _29789_, _29786_);
  or (_29792_, _29791_, _29783_);
  or (_29793_, _29792_, _29775_);
  or (_29794_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand (_29795_, \oc8051_golden_model_1.IRAM[15] [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and (_29796_, _29795_, _29794_);
  and (_29797_, _04399_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and (_29798_, \oc8051_golden_model_1.IRAM[15] [2], _32780_);
  or (_29799_, _29798_, _29797_);
  or (_29800_, _29799_, _29796_);
  and (_29802_, _03791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and (_29803_, \oc8051_golden_model_1.IRAM[15] [0], _32774_);
  or (_29804_, _29803_, _29802_);
  and (_29805_, _03973_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and (_29806_, \oc8051_golden_model_1.IRAM[15] [1], _32777_);
  or (_29807_, _29806_, _29805_);
  or (_29808_, _29807_, _29804_);
  or (_29809_, _29808_, _29800_);
  or (_29810_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand (_29811_, \oc8051_golden_model_1.IRAM[15] [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and (_29813_, _29811_, _29810_);
  and (_29814_, \oc8051_golden_model_1.IRAM[15] [7], _32434_);
  and (_29815_, _04571_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  or (_29816_, _29815_, _29814_);
  or (_29817_, _29816_, _29813_);
  or (_29818_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nand (_29819_, \oc8051_golden_model_1.IRAM[15] [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and (_29820_, _29819_, _29818_);
  or (_29821_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand (_29822_, \oc8051_golden_model_1.IRAM[15] [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and (_29824_, _29822_, _29821_);
  or (_29825_, _29824_, _29820_);
  or (_29826_, _29825_, _29817_);
  or (_29827_, _29826_, _29809_);
  or (_29828_, _29827_, _29793_);
  or (_29829_, _29828_, _29758_);
  or (_29830_, _29829_, _29689_);
  or (_29831_, _29830_, _29550_);
  and (property_invalid_iram, _29831_, _29101_);
  nand (_29832_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_29834_, \oc8051_golden_model_1.DPH [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_29835_, _29834_, _29832_);
  and (_29836_, _16136_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  nor (_29837_, _16136_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_29838_, _29837_, _29836_);
  or (_29839_, _29838_, _29835_);
  nor (_29840_, _09337_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_29841_, _09337_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_29842_, _29841_, _29840_);
  and (_29843_, _16042_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_29845_, _16042_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_29846_, _29845_, _29843_);
  or (_29847_, _29846_, _29842_);
  or (_29848_, _29847_, _29839_);
  or (_29849_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  nand (_29850_, \oc8051_golden_model_1.DPH [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_29851_, _29850_, _29849_);
  or (_29852_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nand (_29853_, \oc8051_golden_model_1.DPH [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_29854_, _29853_, _29852_);
  or (_29856_, _29854_, _29851_);
  and (_29857_, _08280_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  nor (_29858_, _08280_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_29859_, _29858_, _29857_);
  nand (_29860_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_29861_, \oc8051_golden_model_1.DPH [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_29862_, _29861_, _29860_);
  or (_29863_, _29862_, _29859_);
  or (_29864_, _29863_, _29856_);
  or (_29865_, _29864_, _29848_);
  and (property_invalid_dph, _29865_, _29101_);
  nand (_29867_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  or (_29868_, \oc8051_golden_model_1.DPL [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_29869_, _29868_, _29867_);
  and (_29870_, _15497_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_29871_, \oc8051_golden_model_1.DPL [2], _31187_);
  or (_29872_, _29871_, _29870_);
  or (_29873_, _29872_, _29869_);
  and (_29874_, \oc8051_golden_model_1.DPL [0], _31179_);
  and (_29875_, _15313_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or (_29877_, _29875_, _29874_);
  and (_29878_, _15401_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_29879_, \oc8051_golden_model_1.DPL [1], _31183_);
  or (_29880_, _29879_, _29878_);
  or (_29881_, _29880_, _29877_);
  or (_29882_, _29881_, _29873_);
  or (_29883_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand (_29884_, \oc8051_golden_model_1.DPL [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_29885_, _29884_, _29883_);
  or (_29886_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand (_29888_, \oc8051_golden_model_1.DPL [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_29889_, _29888_, _29886_);
  or (_29890_, _29889_, _29885_);
  and (_29891_, _08185_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_29892_, \oc8051_golden_model_1.DPL [7], _30958_);
  or (_29893_, _29892_, _29891_);
  nand (_29894_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_29895_, \oc8051_golden_model_1.DPL [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_29896_, _29895_, _29894_);
  or (_29897_, _29896_, _29893_);
  or (_29899_, _29897_, _29890_);
  or (_29900_, _29899_, _29882_);
  and (property_invalid_dpl, _29900_, _29101_);
  nand (_29901_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_29902_, \oc8051_golden_model_1.B [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_29903_, _29902_, _29901_);
  and (_29904_, _06753_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_29905_, \oc8051_golden_model_1.B [2], _29919_);
  or (_29906_, _29905_, _29904_);
  or (_29907_, _29906_, _29903_);
  and (_29909_, \oc8051_golden_model_1.B [0], _28589_);
  and (_29910_, _06743_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_29911_, _29910_, _29909_);
  and (_29912_, _06738_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_29913_, \oc8051_golden_model_1.B [1], _29274_);
  or (_29914_, _29913_, _29912_);
  or (_29915_, _29914_, _29911_);
  or (_29916_, _29915_, _29907_);
  or (_29917_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_29918_, \oc8051_golden_model_1.B [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_29920_, _29918_, _29917_);
  or (_29921_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_29922_, \oc8051_golden_model_1.B [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_29923_, _29922_, _29921_);
  or (_29924_, _29923_, _29920_);
  and (_29925_, _06159_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_29926_, \oc8051_golden_model_1.B [7], _27529_);
  or (_29927_, _29926_, _29925_);
  nand (_29928_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_29929_, \oc8051_golden_model_1.B [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_29931_, _29929_, _29928_);
  or (_29932_, _29931_, _29927_);
  or (_29933_, _29932_, _29924_);
  or (_29934_, _29933_, _29916_);
  and (property_invalid_b_reg, _29934_, _29101_);
  nand (_29935_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_29936_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_29937_, _29936_, _29935_);
  and (_29938_, _06908_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_29939_, \oc8051_golden_model_1.ACC [2], _31365_);
  or (_29941_, _29939_, _29938_);
  or (_29942_, _29941_, _29937_);
  nor (_29943_, _02477_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_29944_, _02477_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_29945_, _29944_, _29943_);
  and (_29946_, _02658_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_29947_, _02658_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_29948_, _29947_, _29946_);
  or (_29949_, _29948_, _29945_);
  or (_29950_, _29949_, _29942_);
  or (_29952_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_29953_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_29954_, _29953_, _29952_);
  or (_29955_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_29956_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_29957_, _29956_, _29955_);
  or (_29958_, _29957_, _29954_);
  and (_29959_, _06762_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_29960_, _06762_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_29961_, _29960_, _29959_);
  nand (_29963_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_29964_, \oc8051_golden_model_1.ACC [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_29965_, _29964_, _29963_);
  or (_29966_, _29965_, _29961_);
  or (_29967_, _29966_, _29958_);
  or (_29968_, _29967_, _29950_);
  and (property_invalid_acc, _29968_, _29101_);
  nor (_29969_, _20292_, _35039_);
  and (_29970_, _20292_, _35039_);
  nor (_29971_, _20662_, _35043_);
  and (_29973_, _20662_, _35043_);
  and (_29974_, _22122_, _35059_);
  nor (_29975_, _22122_, _35059_);
  nor (_29976_, _23154_, _30879_);
  and (_29977_, _23154_, _30879_);
  nand (_29978_, _22825_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_29979_, _22825_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_29980_, _29979_, _29978_);
  and (_29981_, _24099_, _30890_);
  nor (_29982_, _24099_, _30890_);
  nor (_29984_, _19902_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_29985_, _19902_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_29986_, _29985_, _29984_);
  or (_29987_, _29986_, _29982_);
  or (_29988_, _29987_, _29981_);
  nor (_29989_, _23786_, _30869_);
  and (_29990_, _23786_, _30869_);
  or (_29991_, _29990_, _29989_);
  or (_29992_, _29991_, _29988_);
  and (_29993_, _09712_, _30901_);
  nor (_29995_, _09712_, _30901_);
  or (_29996_, _29995_, _29993_);
  or (_29997_, _29996_, _29992_);
  nor (_29998_, _24722_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_29999_, _24722_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_30000_, _23470_, _30884_);
  nor (_30001_, _23470_, _30884_);
  or (_30002_, _30001_, _30000_);
  nor (_30003_, _24417_, _30865_);
  and (_30004_, _24417_, _30865_);
  or (_30006_, _30004_, _30003_);
  or (_30007_, _30006_, _30002_);
  or (_30008_, _30007_, _29999_);
  or (_30009_, _30008_, _29998_);
  or (_30010_, _30009_, _29997_);
  or (_30011_, _30010_, _29980_);
  or (_30012_, _30011_, _29977_);
  or (_30013_, _30012_, _29976_);
  nor (_30014_, _21395_, _35051_);
  and (_30015_, _21395_, _35051_);
  or (_30017_, _30015_, _30014_);
  or (_30018_, _30017_, _30013_);
  or (_30019_, _30018_, _29975_);
  or (_30020_, _30019_, _29974_);
  and (_30021_, _22487_, _35063_);
  nor (_30022_, _21027_, _35047_);
  or (_30023_, _30022_, _30021_);
  nor (_30024_, _22487_, _35063_);
  and (_30025_, _21027_, _35047_);
  or (_30026_, _30025_, _30024_);
  or (_30028_, _30026_, _30023_);
  or (_30029_, _30028_, _30020_);
  nor (_30030_, _21767_, _35055_);
  and (_30031_, _21767_, _35055_);
  or (_30032_, _30031_, _30030_);
  or (_30033_, _30032_, _30029_);
  or (_30034_, _30033_, _29973_);
  or (_30035_, _30034_, _29971_);
  or (_30036_, _30035_, _29970_);
  or (_30037_, _30036_, _29969_);
  and (property_invalid_pc, _30037_, _28449_);
  buf (_35585_, _35583_);
  buf (_35599_, _35583_);
  buf (_35601_, _35583_);
  buf (_35603_, _35583_);
  buf (_35605_, _35583_);
  buf (_35607_, _35583_);
  buf (_35609_, _35583_);
  buf (_35611_, _35583_);
  buf (_35613_, _35583_);
  buf (_35587_, _35583_);
  buf (_35589_, _35583_);
  buf (_35591_, _35583_);
  buf (_35593_, _35583_);
  buf (_35595_, _35583_);
  buf (_35597_, _35583_);
  buf (_35798_[7], _35777_[7]);
  buf (_35799_[7], _35778_[7]);
  buf (_35810_[7], _35777_[7]);
  buf (_35811_[7], _35778_[7]);
  buf (_35798_[0], _35777_[0]);
  buf (_35798_[1], _35777_[1]);
  buf (_35798_[2], _35777_[2]);
  buf (_35798_[3], _35777_[3]);
  buf (_35798_[4], _35777_[4]);
  buf (_35798_[5], _35777_[5]);
  buf (_35798_[6], _35777_[6]);
  buf (_35799_[0], _35778_[0]);
  buf (_35799_[1], _35778_[1]);
  buf (_35799_[2], _35778_[2]);
  buf (_35799_[3], _35778_[3]);
  buf (_35799_[4], _35778_[4]);
  buf (_35799_[5], _35778_[5]);
  buf (_35799_[6], _35778_[6]);
  buf (_35810_[0], _35777_[0]);
  buf (_35810_[1], _35777_[1]);
  buf (_35810_[2], _35777_[2]);
  buf (_35810_[3], _35777_[3]);
  buf (_35810_[4], _35777_[4]);
  buf (_35810_[5], _35777_[5]);
  buf (_35810_[6], _35777_[6]);
  buf (_35811_[0], _35778_[0]);
  buf (_35811_[1], _35778_[1]);
  buf (_35811_[2], _35778_[2]);
  buf (_35811_[3], _35778_[3]);
  buf (_35811_[4], _35778_[4]);
  buf (_35811_[5], _35778_[5]);
  buf (_35811_[6], _35778_[6]);
  buf (_35964_, _35792_);
  buf (_35830_, _35792_);
  dff (p0in_reg[0], _00002_[0]);
  dff (p0in_reg[1], _00002_[1]);
  dff (p0in_reg[2], _00002_[2]);
  dff (p0in_reg[3], _00002_[3]);
  dff (p0in_reg[4], _00002_[4]);
  dff (p0in_reg[5], _00002_[5]);
  dff (p0in_reg[6], _00002_[6]);
  dff (p0in_reg[7], _00002_[7]);
  dff (p1in_reg[0], _00003_[0]);
  dff (p1in_reg[1], _00003_[1]);
  dff (p1in_reg[2], _00003_[2]);
  dff (p1in_reg[3], _00003_[3]);
  dff (p1in_reg[4], _00003_[4]);
  dff (p1in_reg[5], _00003_[5]);
  dff (p1in_reg[6], _00003_[6]);
  dff (p1in_reg[7], _00003_[7]);
  dff (p2in_reg[0], _00004_[0]);
  dff (p2in_reg[1], _00004_[1]);
  dff (p2in_reg[2], _00004_[2]);
  dff (p2in_reg[3], _00004_[3]);
  dff (p2in_reg[4], _00004_[4]);
  dff (p2in_reg[5], _00004_[5]);
  dff (p2in_reg[6], _00004_[6]);
  dff (p2in_reg[7], _00004_[7]);
  dff (p3in_reg[0], _00005_[0]);
  dff (p3in_reg[1], _00005_[1]);
  dff (p3in_reg[2], _00005_[2]);
  dff (p3in_reg[3], _00005_[3]);
  dff (p3in_reg[4], _00005_[4]);
  dff (p3in_reg[5], _00005_[5]);
  dff (p3in_reg[6], _00005_[6]);
  dff (p3in_reg[7], _00005_[7]);
  dff (op0_cnst, _00001_);
  dff (inst_finished_r, _00000_);
  dff (property_invalid_psw_1_r, _00006_);
  dff (property_invalid_sp_1_r, _00007_);
  dff (\oc8051_gm_cxrom_1.cell0.data [0], _35582_[0]);
  dff (\oc8051_gm_cxrom_1.cell0.data [1], _35582_[1]);
  dff (\oc8051_gm_cxrom_1.cell0.data [2], _35582_[2]);
  dff (\oc8051_gm_cxrom_1.cell0.data [3], _35582_[3]);
  dff (\oc8051_gm_cxrom_1.cell0.data [4], _35582_[4]);
  dff (\oc8051_gm_cxrom_1.cell0.data [5], _35582_[5]);
  dff (\oc8051_gm_cxrom_1.cell0.data [6], _35582_[6]);
  dff (\oc8051_gm_cxrom_1.cell0.data [7], _35582_[7]);
  dff (\oc8051_gm_cxrom_1.cell0.valid , _35583_);
  dff (\oc8051_gm_cxrom_1.cell1.data [0], _35584_[0]);
  dff (\oc8051_gm_cxrom_1.cell1.data [1], _35584_[1]);
  dff (\oc8051_gm_cxrom_1.cell1.data [2], _35584_[2]);
  dff (\oc8051_gm_cxrom_1.cell1.data [3], _35584_[3]);
  dff (\oc8051_gm_cxrom_1.cell1.data [4], _35584_[4]);
  dff (\oc8051_gm_cxrom_1.cell1.data [5], _35584_[5]);
  dff (\oc8051_gm_cxrom_1.cell1.data [6], _35584_[6]);
  dff (\oc8051_gm_cxrom_1.cell1.data [7], _35584_[7]);
  dff (\oc8051_gm_cxrom_1.cell1.valid , _35585_);
  dff (\oc8051_gm_cxrom_1.cell10.data [0], _35586_[0]);
  dff (\oc8051_gm_cxrom_1.cell10.data [1], _35586_[1]);
  dff (\oc8051_gm_cxrom_1.cell10.data [2], _35586_[2]);
  dff (\oc8051_gm_cxrom_1.cell10.data [3], _35586_[3]);
  dff (\oc8051_gm_cxrom_1.cell10.data [4], _35586_[4]);
  dff (\oc8051_gm_cxrom_1.cell10.data [5], _35586_[5]);
  dff (\oc8051_gm_cxrom_1.cell10.data [6], _35586_[6]);
  dff (\oc8051_gm_cxrom_1.cell10.data [7], _35586_[7]);
  dff (\oc8051_gm_cxrom_1.cell10.valid , _35587_);
  dff (\oc8051_gm_cxrom_1.cell11.data [0], _35588_[0]);
  dff (\oc8051_gm_cxrom_1.cell11.data [1], _35588_[1]);
  dff (\oc8051_gm_cxrom_1.cell11.data [2], _35588_[2]);
  dff (\oc8051_gm_cxrom_1.cell11.data [3], _35588_[3]);
  dff (\oc8051_gm_cxrom_1.cell11.data [4], _35588_[4]);
  dff (\oc8051_gm_cxrom_1.cell11.data [5], _35588_[5]);
  dff (\oc8051_gm_cxrom_1.cell11.data [6], _35588_[6]);
  dff (\oc8051_gm_cxrom_1.cell11.data [7], _35588_[7]);
  dff (\oc8051_gm_cxrom_1.cell11.valid , _35589_);
  dff (\oc8051_gm_cxrom_1.cell12.data [0], _35590_[0]);
  dff (\oc8051_gm_cxrom_1.cell12.data [1], _35590_[1]);
  dff (\oc8051_gm_cxrom_1.cell12.data [2], _35590_[2]);
  dff (\oc8051_gm_cxrom_1.cell12.data [3], _35590_[3]);
  dff (\oc8051_gm_cxrom_1.cell12.data [4], _35590_[4]);
  dff (\oc8051_gm_cxrom_1.cell12.data [5], _35590_[5]);
  dff (\oc8051_gm_cxrom_1.cell12.data [6], _35590_[6]);
  dff (\oc8051_gm_cxrom_1.cell12.data [7], _35590_[7]);
  dff (\oc8051_gm_cxrom_1.cell12.valid , _35591_);
  dff (\oc8051_gm_cxrom_1.cell13.data [0], _35592_[0]);
  dff (\oc8051_gm_cxrom_1.cell13.data [1], _35592_[1]);
  dff (\oc8051_gm_cxrom_1.cell13.data [2], _35592_[2]);
  dff (\oc8051_gm_cxrom_1.cell13.data [3], _35592_[3]);
  dff (\oc8051_gm_cxrom_1.cell13.data [4], _35592_[4]);
  dff (\oc8051_gm_cxrom_1.cell13.data [5], _35592_[5]);
  dff (\oc8051_gm_cxrom_1.cell13.data [6], _35592_[6]);
  dff (\oc8051_gm_cxrom_1.cell13.data [7], _35592_[7]);
  dff (\oc8051_gm_cxrom_1.cell13.valid , _35593_);
  dff (\oc8051_gm_cxrom_1.cell14.data [0], _35594_[0]);
  dff (\oc8051_gm_cxrom_1.cell14.data [1], _35594_[1]);
  dff (\oc8051_gm_cxrom_1.cell14.data [2], _35594_[2]);
  dff (\oc8051_gm_cxrom_1.cell14.data [3], _35594_[3]);
  dff (\oc8051_gm_cxrom_1.cell14.data [4], _35594_[4]);
  dff (\oc8051_gm_cxrom_1.cell14.data [5], _35594_[5]);
  dff (\oc8051_gm_cxrom_1.cell14.data [6], _35594_[6]);
  dff (\oc8051_gm_cxrom_1.cell14.data [7], _35594_[7]);
  dff (\oc8051_gm_cxrom_1.cell14.valid , _35595_);
  dff (\oc8051_gm_cxrom_1.cell15.data [0], _35596_[0]);
  dff (\oc8051_gm_cxrom_1.cell15.data [1], _35596_[1]);
  dff (\oc8051_gm_cxrom_1.cell15.data [2], _35596_[2]);
  dff (\oc8051_gm_cxrom_1.cell15.data [3], _35596_[3]);
  dff (\oc8051_gm_cxrom_1.cell15.data [4], _35596_[4]);
  dff (\oc8051_gm_cxrom_1.cell15.data [5], _35596_[5]);
  dff (\oc8051_gm_cxrom_1.cell15.data [6], _35596_[6]);
  dff (\oc8051_gm_cxrom_1.cell15.data [7], _35596_[7]);
  dff (\oc8051_gm_cxrom_1.cell15.valid , _35597_);
  dff (\oc8051_gm_cxrom_1.cell2.data [0], _35598_[0]);
  dff (\oc8051_gm_cxrom_1.cell2.data [1], _35598_[1]);
  dff (\oc8051_gm_cxrom_1.cell2.data [2], _35598_[2]);
  dff (\oc8051_gm_cxrom_1.cell2.data [3], _35598_[3]);
  dff (\oc8051_gm_cxrom_1.cell2.data [4], _35598_[4]);
  dff (\oc8051_gm_cxrom_1.cell2.data [5], _35598_[5]);
  dff (\oc8051_gm_cxrom_1.cell2.data [6], _35598_[6]);
  dff (\oc8051_gm_cxrom_1.cell2.data [7], _35598_[7]);
  dff (\oc8051_gm_cxrom_1.cell2.valid , _35599_);
  dff (\oc8051_gm_cxrom_1.cell3.data [0], _35600_[0]);
  dff (\oc8051_gm_cxrom_1.cell3.data [1], _35600_[1]);
  dff (\oc8051_gm_cxrom_1.cell3.data [2], _35600_[2]);
  dff (\oc8051_gm_cxrom_1.cell3.data [3], _35600_[3]);
  dff (\oc8051_gm_cxrom_1.cell3.data [4], _35600_[4]);
  dff (\oc8051_gm_cxrom_1.cell3.data [5], _35600_[5]);
  dff (\oc8051_gm_cxrom_1.cell3.data [6], _35600_[6]);
  dff (\oc8051_gm_cxrom_1.cell3.data [7], _35600_[7]);
  dff (\oc8051_gm_cxrom_1.cell3.valid , _35601_);
  dff (\oc8051_gm_cxrom_1.cell4.data [0], _35602_[0]);
  dff (\oc8051_gm_cxrom_1.cell4.data [1], _35602_[1]);
  dff (\oc8051_gm_cxrom_1.cell4.data [2], _35602_[2]);
  dff (\oc8051_gm_cxrom_1.cell4.data [3], _35602_[3]);
  dff (\oc8051_gm_cxrom_1.cell4.data [4], _35602_[4]);
  dff (\oc8051_gm_cxrom_1.cell4.data [5], _35602_[5]);
  dff (\oc8051_gm_cxrom_1.cell4.data [6], _35602_[6]);
  dff (\oc8051_gm_cxrom_1.cell4.data [7], _35602_[7]);
  dff (\oc8051_gm_cxrom_1.cell4.valid , _35603_);
  dff (\oc8051_gm_cxrom_1.cell5.data [0], _35604_[0]);
  dff (\oc8051_gm_cxrom_1.cell5.data [1], _35604_[1]);
  dff (\oc8051_gm_cxrom_1.cell5.data [2], _35604_[2]);
  dff (\oc8051_gm_cxrom_1.cell5.data [3], _35604_[3]);
  dff (\oc8051_gm_cxrom_1.cell5.data [4], _35604_[4]);
  dff (\oc8051_gm_cxrom_1.cell5.data [5], _35604_[5]);
  dff (\oc8051_gm_cxrom_1.cell5.data [6], _35604_[6]);
  dff (\oc8051_gm_cxrom_1.cell5.data [7], _35604_[7]);
  dff (\oc8051_gm_cxrom_1.cell5.valid , _35605_);
  dff (\oc8051_gm_cxrom_1.cell6.data [0], _35606_[0]);
  dff (\oc8051_gm_cxrom_1.cell6.data [1], _35606_[1]);
  dff (\oc8051_gm_cxrom_1.cell6.data [2], _35606_[2]);
  dff (\oc8051_gm_cxrom_1.cell6.data [3], _35606_[3]);
  dff (\oc8051_gm_cxrom_1.cell6.data [4], _35606_[4]);
  dff (\oc8051_gm_cxrom_1.cell6.data [5], _35606_[5]);
  dff (\oc8051_gm_cxrom_1.cell6.data [6], _35606_[6]);
  dff (\oc8051_gm_cxrom_1.cell6.data [7], _35606_[7]);
  dff (\oc8051_gm_cxrom_1.cell6.valid , _35607_);
  dff (\oc8051_gm_cxrom_1.cell7.data [0], _35608_[0]);
  dff (\oc8051_gm_cxrom_1.cell7.data [1], _35608_[1]);
  dff (\oc8051_gm_cxrom_1.cell7.data [2], _35608_[2]);
  dff (\oc8051_gm_cxrom_1.cell7.data [3], _35608_[3]);
  dff (\oc8051_gm_cxrom_1.cell7.data [4], _35608_[4]);
  dff (\oc8051_gm_cxrom_1.cell7.data [5], _35608_[5]);
  dff (\oc8051_gm_cxrom_1.cell7.data [6], _35608_[6]);
  dff (\oc8051_gm_cxrom_1.cell7.data [7], _35608_[7]);
  dff (\oc8051_gm_cxrom_1.cell7.valid , _35609_);
  dff (\oc8051_gm_cxrom_1.cell8.data [0], _35610_[0]);
  dff (\oc8051_gm_cxrom_1.cell8.data [1], _35610_[1]);
  dff (\oc8051_gm_cxrom_1.cell8.data [2], _35610_[2]);
  dff (\oc8051_gm_cxrom_1.cell8.data [3], _35610_[3]);
  dff (\oc8051_gm_cxrom_1.cell8.data [4], _35610_[4]);
  dff (\oc8051_gm_cxrom_1.cell8.data [5], _35610_[5]);
  dff (\oc8051_gm_cxrom_1.cell8.data [6], _35610_[6]);
  dff (\oc8051_gm_cxrom_1.cell8.data [7], _35610_[7]);
  dff (\oc8051_gm_cxrom_1.cell8.valid , _35611_);
  dff (\oc8051_gm_cxrom_1.cell9.data [0], _35612_[0]);
  dff (\oc8051_gm_cxrom_1.cell9.data [1], _35612_[1]);
  dff (\oc8051_gm_cxrom_1.cell9.data [2], _35612_[2]);
  dff (\oc8051_gm_cxrom_1.cell9.data [3], _35612_[3]);
  dff (\oc8051_gm_cxrom_1.cell9.data [4], _35612_[4]);
  dff (\oc8051_gm_cxrom_1.cell9.data [5], _35612_[5]);
  dff (\oc8051_gm_cxrom_1.cell9.data [6], _35612_[6]);
  dff (\oc8051_gm_cxrom_1.cell9.data [7], _35612_[7]);
  dff (\oc8051_gm_cxrom_1.cell9.valid , _35613_);
  dff (\oc8051_golden_model_1.IRAM[15] [0], _35691_);
  dff (\oc8051_golden_model_1.IRAM[15] [1], _35692_);
  dff (\oc8051_golden_model_1.IRAM[15] [2], _35693_);
  dff (\oc8051_golden_model_1.IRAM[15] [3], _35694_);
  dff (\oc8051_golden_model_1.IRAM[15] [4], _35695_);
  dff (\oc8051_golden_model_1.IRAM[15] [5], _35696_);
  dff (\oc8051_golden_model_1.IRAM[15] [6], _35697_);
  dff (\oc8051_golden_model_1.IRAM[15] [7], _35698_);
  dff (\oc8051_golden_model_1.IRAM[14] [0], _35683_);
  dff (\oc8051_golden_model_1.IRAM[14] [1], _35684_);
  dff (\oc8051_golden_model_1.IRAM[14] [2], _35685_);
  dff (\oc8051_golden_model_1.IRAM[14] [3], _35686_);
  dff (\oc8051_golden_model_1.IRAM[14] [4], _35687_);
  dff (\oc8051_golden_model_1.IRAM[14] [5], _35688_);
  dff (\oc8051_golden_model_1.IRAM[14] [6], _35689_);
  dff (\oc8051_golden_model_1.IRAM[14] [7], _35690_);
  dff (\oc8051_golden_model_1.IRAM[13] [0], _35675_);
  dff (\oc8051_golden_model_1.IRAM[13] [1], _35676_);
  dff (\oc8051_golden_model_1.IRAM[13] [2], _35677_);
  dff (\oc8051_golden_model_1.IRAM[13] [3], _35678_);
  dff (\oc8051_golden_model_1.IRAM[13] [4], _35679_);
  dff (\oc8051_golden_model_1.IRAM[13] [5], _35680_);
  dff (\oc8051_golden_model_1.IRAM[13] [6], _35681_);
  dff (\oc8051_golden_model_1.IRAM[13] [7], _35682_);
  dff (\oc8051_golden_model_1.IRAM[12] [0], _35667_);
  dff (\oc8051_golden_model_1.IRAM[12] [1], _35668_);
  dff (\oc8051_golden_model_1.IRAM[12] [2], _35669_);
  dff (\oc8051_golden_model_1.IRAM[12] [3], _35670_);
  dff (\oc8051_golden_model_1.IRAM[12] [4], _35671_);
  dff (\oc8051_golden_model_1.IRAM[12] [5], _35672_);
  dff (\oc8051_golden_model_1.IRAM[12] [6], _35673_);
  dff (\oc8051_golden_model_1.IRAM[12] [7], _35674_);
  dff (\oc8051_golden_model_1.IRAM[11] [0], _35659_);
  dff (\oc8051_golden_model_1.IRAM[11] [1], _35660_);
  dff (\oc8051_golden_model_1.IRAM[11] [2], _35661_);
  dff (\oc8051_golden_model_1.IRAM[11] [3], _35662_);
  dff (\oc8051_golden_model_1.IRAM[11] [4], _35663_);
  dff (\oc8051_golden_model_1.IRAM[11] [5], _35664_);
  dff (\oc8051_golden_model_1.IRAM[11] [6], _35665_);
  dff (\oc8051_golden_model_1.IRAM[11] [7], _35666_);
  dff (\oc8051_golden_model_1.IRAM[10] [0], _35651_);
  dff (\oc8051_golden_model_1.IRAM[10] [1], _35652_);
  dff (\oc8051_golden_model_1.IRAM[10] [2], _35653_);
  dff (\oc8051_golden_model_1.IRAM[10] [3], _35654_);
  dff (\oc8051_golden_model_1.IRAM[10] [4], _35655_);
  dff (\oc8051_golden_model_1.IRAM[10] [5], _35656_);
  dff (\oc8051_golden_model_1.IRAM[10] [6], _35657_);
  dff (\oc8051_golden_model_1.IRAM[10] [7], _35658_);
  dff (\oc8051_golden_model_1.IRAM[9] [0], _35763_);
  dff (\oc8051_golden_model_1.IRAM[9] [1], _35764_);
  dff (\oc8051_golden_model_1.IRAM[9] [2], _35765_);
  dff (\oc8051_golden_model_1.IRAM[9] [3], _35766_);
  dff (\oc8051_golden_model_1.IRAM[9] [4], _35767_);
  dff (\oc8051_golden_model_1.IRAM[9] [5], _35768_);
  dff (\oc8051_golden_model_1.IRAM[9] [6], _35769_);
  dff (\oc8051_golden_model_1.IRAM[9] [7], _35770_);
  dff (\oc8051_golden_model_1.IRAM[8] [0], _35755_);
  dff (\oc8051_golden_model_1.IRAM[8] [1], _35756_);
  dff (\oc8051_golden_model_1.IRAM[8] [2], _35757_);
  dff (\oc8051_golden_model_1.IRAM[8] [3], _35758_);
  dff (\oc8051_golden_model_1.IRAM[8] [4], _35759_);
  dff (\oc8051_golden_model_1.IRAM[8] [5], _35760_);
  dff (\oc8051_golden_model_1.IRAM[8] [6], _35761_);
  dff (\oc8051_golden_model_1.IRAM[8] [7], _35762_);
  dff (\oc8051_golden_model_1.IRAM[7] [0], _35747_);
  dff (\oc8051_golden_model_1.IRAM[7] [1], _35748_);
  dff (\oc8051_golden_model_1.IRAM[7] [2], _35749_);
  dff (\oc8051_golden_model_1.IRAM[7] [3], _35750_);
  dff (\oc8051_golden_model_1.IRAM[7] [4], _35751_);
  dff (\oc8051_golden_model_1.IRAM[7] [5], _35752_);
  dff (\oc8051_golden_model_1.IRAM[7] [6], _35753_);
  dff (\oc8051_golden_model_1.IRAM[7] [7], _35754_);
  dff (\oc8051_golden_model_1.IRAM[6] [0], _35739_);
  dff (\oc8051_golden_model_1.IRAM[6] [1], _35740_);
  dff (\oc8051_golden_model_1.IRAM[6] [2], _35741_);
  dff (\oc8051_golden_model_1.IRAM[6] [3], _35742_);
  dff (\oc8051_golden_model_1.IRAM[6] [4], _35743_);
  dff (\oc8051_golden_model_1.IRAM[6] [5], _35744_);
  dff (\oc8051_golden_model_1.IRAM[6] [6], _35745_);
  dff (\oc8051_golden_model_1.IRAM[6] [7], _35746_);
  dff (\oc8051_golden_model_1.IRAM[5] [0], _35731_);
  dff (\oc8051_golden_model_1.IRAM[5] [1], _35732_);
  dff (\oc8051_golden_model_1.IRAM[5] [2], _35733_);
  dff (\oc8051_golden_model_1.IRAM[5] [3], _35734_);
  dff (\oc8051_golden_model_1.IRAM[5] [4], _35735_);
  dff (\oc8051_golden_model_1.IRAM[5] [5], _35736_);
  dff (\oc8051_golden_model_1.IRAM[5] [6], _35737_);
  dff (\oc8051_golden_model_1.IRAM[5] [7], _35738_);
  dff (\oc8051_golden_model_1.IRAM[4] [0], _35723_);
  dff (\oc8051_golden_model_1.IRAM[4] [1], _35724_);
  dff (\oc8051_golden_model_1.IRAM[4] [2], _35725_);
  dff (\oc8051_golden_model_1.IRAM[4] [3], _35726_);
  dff (\oc8051_golden_model_1.IRAM[4] [4], _35727_);
  dff (\oc8051_golden_model_1.IRAM[4] [5], _35728_);
  dff (\oc8051_golden_model_1.IRAM[4] [6], _35729_);
  dff (\oc8051_golden_model_1.IRAM[4] [7], _35730_);
  dff (\oc8051_golden_model_1.IRAM[3] [0], _35715_);
  dff (\oc8051_golden_model_1.IRAM[3] [1], _35716_);
  dff (\oc8051_golden_model_1.IRAM[3] [2], _35717_);
  dff (\oc8051_golden_model_1.IRAM[3] [3], _35718_);
  dff (\oc8051_golden_model_1.IRAM[3] [4], _35719_);
  dff (\oc8051_golden_model_1.IRAM[3] [5], _35720_);
  dff (\oc8051_golden_model_1.IRAM[3] [6], _35721_);
  dff (\oc8051_golden_model_1.IRAM[3] [7], _35722_);
  dff (\oc8051_golden_model_1.IRAM[2] [0], _35707_);
  dff (\oc8051_golden_model_1.IRAM[2] [1], _35708_);
  dff (\oc8051_golden_model_1.IRAM[2] [2], _35709_);
  dff (\oc8051_golden_model_1.IRAM[2] [3], _35710_);
  dff (\oc8051_golden_model_1.IRAM[2] [4], _35711_);
  dff (\oc8051_golden_model_1.IRAM[2] [5], _35712_);
  dff (\oc8051_golden_model_1.IRAM[2] [6], _35713_);
  dff (\oc8051_golden_model_1.IRAM[2] [7], _35714_);
  dff (\oc8051_golden_model_1.IRAM[1] [0], _35699_);
  dff (\oc8051_golden_model_1.IRAM[1] [1], _35700_);
  dff (\oc8051_golden_model_1.IRAM[1] [2], _35701_);
  dff (\oc8051_golden_model_1.IRAM[1] [3], _35702_);
  dff (\oc8051_golden_model_1.IRAM[1] [4], _35703_);
  dff (\oc8051_golden_model_1.IRAM[1] [5], _35704_);
  dff (\oc8051_golden_model_1.IRAM[1] [6], _35705_);
  dff (\oc8051_golden_model_1.IRAM[1] [7], _35706_);
  dff (\oc8051_golden_model_1.IRAM[0] [0], _35643_);
  dff (\oc8051_golden_model_1.IRAM[0] [1], _35644_);
  dff (\oc8051_golden_model_1.IRAM[0] [2], _35645_);
  dff (\oc8051_golden_model_1.IRAM[0] [3], _35646_);
  dff (\oc8051_golden_model_1.IRAM[0] [4], _35647_);
  dff (\oc8051_golden_model_1.IRAM[0] [5], _35648_);
  dff (\oc8051_golden_model_1.IRAM[0] [6], _35649_);
  dff (\oc8051_golden_model_1.IRAM[0] [7], _35650_);
  dff (\oc8051_golden_model_1.B [0], _35615_[0]);
  dff (\oc8051_golden_model_1.B [1], _35615_[1]);
  dff (\oc8051_golden_model_1.B [2], _35615_[2]);
  dff (\oc8051_golden_model_1.B [3], _35615_[3]);
  dff (\oc8051_golden_model_1.B [4], _35615_[4]);
  dff (\oc8051_golden_model_1.B [5], _35615_[5]);
  dff (\oc8051_golden_model_1.B [6], _35615_[6]);
  dff (\oc8051_golden_model_1.B [7], _35615_[7]);
  dff (\oc8051_golden_model_1.ACC [0], _35614_[0]);
  dff (\oc8051_golden_model_1.ACC [1], _35614_[1]);
  dff (\oc8051_golden_model_1.ACC [2], _35614_[2]);
  dff (\oc8051_golden_model_1.ACC [3], _35614_[3]);
  dff (\oc8051_golden_model_1.ACC [4], _35614_[4]);
  dff (\oc8051_golden_model_1.ACC [5], _35614_[5]);
  dff (\oc8051_golden_model_1.ACC [6], _35614_[6]);
  dff (\oc8051_golden_model_1.ACC [7], _35614_[7]);
  dff (\oc8051_golden_model_1.DPL [0], _35617_[0]);
  dff (\oc8051_golden_model_1.DPL [1], _35617_[1]);
  dff (\oc8051_golden_model_1.DPL [2], _35617_[2]);
  dff (\oc8051_golden_model_1.DPL [3], _35617_[3]);
  dff (\oc8051_golden_model_1.DPL [4], _35617_[4]);
  dff (\oc8051_golden_model_1.DPL [5], _35617_[5]);
  dff (\oc8051_golden_model_1.DPL [6], _35617_[6]);
  dff (\oc8051_golden_model_1.DPL [7], _35617_[7]);
  dff (\oc8051_golden_model_1.DPH [0], _35616_[0]);
  dff (\oc8051_golden_model_1.DPH [1], _35616_[1]);
  dff (\oc8051_golden_model_1.DPH [2], _35616_[2]);
  dff (\oc8051_golden_model_1.DPH [3], _35616_[3]);
  dff (\oc8051_golden_model_1.DPH [4], _35616_[4]);
  dff (\oc8051_golden_model_1.DPH [5], _35616_[5]);
  dff (\oc8051_golden_model_1.DPH [6], _35616_[6]);
  dff (\oc8051_golden_model_1.DPH [7], _35616_[7]);
  dff (\oc8051_golden_model_1.IE [0], _35618_[0]);
  dff (\oc8051_golden_model_1.IE [1], _35618_[1]);
  dff (\oc8051_golden_model_1.IE [2], _35618_[2]);
  dff (\oc8051_golden_model_1.IE [3], _35618_[3]);
  dff (\oc8051_golden_model_1.IE [4], _35618_[4]);
  dff (\oc8051_golden_model_1.IE [5], _35618_[5]);
  dff (\oc8051_golden_model_1.IE [6], _35618_[6]);
  dff (\oc8051_golden_model_1.IE [7], _35618_[7]);
  dff (\oc8051_golden_model_1.IP [0], _35619_[0]);
  dff (\oc8051_golden_model_1.IP [1], _35619_[1]);
  dff (\oc8051_golden_model_1.IP [2], _35619_[2]);
  dff (\oc8051_golden_model_1.IP [3], _35619_[3]);
  dff (\oc8051_golden_model_1.IP [4], _35619_[4]);
  dff (\oc8051_golden_model_1.IP [5], _35619_[5]);
  dff (\oc8051_golden_model_1.IP [6], _35619_[6]);
  dff (\oc8051_golden_model_1.IP [7], _35619_[7]);
  dff (\oc8051_golden_model_1.P0 [0], _35621_[0]);
  dff (\oc8051_golden_model_1.P0 [1], _35621_[1]);
  dff (\oc8051_golden_model_1.P0 [2], _35621_[2]);
  dff (\oc8051_golden_model_1.P0 [3], _35621_[3]);
  dff (\oc8051_golden_model_1.P0 [4], _35621_[4]);
  dff (\oc8051_golden_model_1.P0 [5], _35621_[5]);
  dff (\oc8051_golden_model_1.P0 [6], _35621_[6]);
  dff (\oc8051_golden_model_1.P0 [7], _35621_[7]);
  dff (\oc8051_golden_model_1.P1 [0], _35623_[0]);
  dff (\oc8051_golden_model_1.P1 [1], _35623_[1]);
  dff (\oc8051_golden_model_1.P1 [2], _35623_[2]);
  dff (\oc8051_golden_model_1.P1 [3], _35623_[3]);
  dff (\oc8051_golden_model_1.P1 [4], _35623_[4]);
  dff (\oc8051_golden_model_1.P1 [5], _35623_[5]);
  dff (\oc8051_golden_model_1.P1 [6], _35623_[6]);
  dff (\oc8051_golden_model_1.P1 [7], _35623_[7]);
  dff (\oc8051_golden_model_1.P2 [0], _35625_[0]);
  dff (\oc8051_golden_model_1.P2 [1], _35625_[1]);
  dff (\oc8051_golden_model_1.P2 [2], _35625_[2]);
  dff (\oc8051_golden_model_1.P2 [3], _35625_[3]);
  dff (\oc8051_golden_model_1.P2 [4], _35625_[4]);
  dff (\oc8051_golden_model_1.P2 [5], _35625_[5]);
  dff (\oc8051_golden_model_1.P2 [6], _35625_[6]);
  dff (\oc8051_golden_model_1.P2 [7], _35625_[7]);
  dff (\oc8051_golden_model_1.P3 [0], _35627_[0]);
  dff (\oc8051_golden_model_1.P3 [1], _35627_[1]);
  dff (\oc8051_golden_model_1.P3 [2], _35627_[2]);
  dff (\oc8051_golden_model_1.P3 [3], _35627_[3]);
  dff (\oc8051_golden_model_1.P3 [4], _35627_[4]);
  dff (\oc8051_golden_model_1.P3 [5], _35627_[5]);
  dff (\oc8051_golden_model_1.P3 [6], _35627_[6]);
  dff (\oc8051_golden_model_1.P3 [7], _35627_[7]);
  dff (\oc8051_golden_model_1.PC [0], _35629_[0]);
  dff (\oc8051_golden_model_1.PC [1], _35629_[1]);
  dff (\oc8051_golden_model_1.PC [2], _35629_[2]);
  dff (\oc8051_golden_model_1.PC [3], _35629_[3]);
  dff (\oc8051_golden_model_1.PC [4], _35629_[4]);
  dff (\oc8051_golden_model_1.PC [5], _35629_[5]);
  dff (\oc8051_golden_model_1.PC [6], _35629_[6]);
  dff (\oc8051_golden_model_1.PC [7], _35629_[7]);
  dff (\oc8051_golden_model_1.PC [8], _35629_[8]);
  dff (\oc8051_golden_model_1.PC [9], _35629_[9]);
  dff (\oc8051_golden_model_1.PC [10], _35629_[10]);
  dff (\oc8051_golden_model_1.PC [11], _35629_[11]);
  dff (\oc8051_golden_model_1.PC [12], _35629_[12]);
  dff (\oc8051_golden_model_1.PC [13], _35629_[13]);
  dff (\oc8051_golden_model_1.PC [14], _35629_[14]);
  dff (\oc8051_golden_model_1.PC [15], _35629_[15]);
  dff (\oc8051_golden_model_1.PSW [0], _35630_[0]);
  dff (\oc8051_golden_model_1.PSW [1], _35630_[1]);
  dff (\oc8051_golden_model_1.PSW [2], _35630_[2]);
  dff (\oc8051_golden_model_1.PSW [3], _35630_[3]);
  dff (\oc8051_golden_model_1.PSW [4], _35630_[4]);
  dff (\oc8051_golden_model_1.PSW [5], _35630_[5]);
  dff (\oc8051_golden_model_1.PSW [6], _35630_[6]);
  dff (\oc8051_golden_model_1.PSW [7], _35630_[7]);
  dff (\oc8051_golden_model_1.PCON [0], _35628_[0]);
  dff (\oc8051_golden_model_1.PCON [1], _35628_[1]);
  dff (\oc8051_golden_model_1.PCON [2], _35628_[2]);
  dff (\oc8051_golden_model_1.PCON [3], _35628_[3]);
  dff (\oc8051_golden_model_1.PCON [4], _35628_[4]);
  dff (\oc8051_golden_model_1.PCON [5], _35628_[5]);
  dff (\oc8051_golden_model_1.PCON [6], _35628_[6]);
  dff (\oc8051_golden_model_1.PCON [7], _35628_[7]);
  dff (\oc8051_golden_model_1.SBUF [0], _35631_[0]);
  dff (\oc8051_golden_model_1.SBUF [1], _35631_[1]);
  dff (\oc8051_golden_model_1.SBUF [2], _35631_[2]);
  dff (\oc8051_golden_model_1.SBUF [3], _35631_[3]);
  dff (\oc8051_golden_model_1.SBUF [4], _35631_[4]);
  dff (\oc8051_golden_model_1.SBUF [5], _35631_[5]);
  dff (\oc8051_golden_model_1.SBUF [6], _35631_[6]);
  dff (\oc8051_golden_model_1.SBUF [7], _35631_[7]);
  dff (\oc8051_golden_model_1.SCON [0], _35632_[0]);
  dff (\oc8051_golden_model_1.SCON [1], _35632_[1]);
  dff (\oc8051_golden_model_1.SCON [2], _35632_[2]);
  dff (\oc8051_golden_model_1.SCON [3], _35632_[3]);
  dff (\oc8051_golden_model_1.SCON [4], _35632_[4]);
  dff (\oc8051_golden_model_1.SCON [5], _35632_[5]);
  dff (\oc8051_golden_model_1.SCON [6], _35632_[6]);
  dff (\oc8051_golden_model_1.SCON [7], _35632_[7]);
  dff (\oc8051_golden_model_1.SP [0], _35633_[0]);
  dff (\oc8051_golden_model_1.SP [1], _35633_[1]);
  dff (\oc8051_golden_model_1.SP [2], _35633_[2]);
  dff (\oc8051_golden_model_1.SP [3], _35633_[3]);
  dff (\oc8051_golden_model_1.SP [4], _35633_[4]);
  dff (\oc8051_golden_model_1.SP [5], _35633_[5]);
  dff (\oc8051_golden_model_1.SP [6], _35633_[6]);
  dff (\oc8051_golden_model_1.SP [7], _35633_[7]);
  dff (\oc8051_golden_model_1.TCON [0], _35634_[0]);
  dff (\oc8051_golden_model_1.TCON [1], _35634_[1]);
  dff (\oc8051_golden_model_1.TCON [2], _35634_[2]);
  dff (\oc8051_golden_model_1.TCON [3], _35634_[3]);
  dff (\oc8051_golden_model_1.TCON [4], _35634_[4]);
  dff (\oc8051_golden_model_1.TCON [5], _35634_[5]);
  dff (\oc8051_golden_model_1.TCON [6], _35634_[6]);
  dff (\oc8051_golden_model_1.TCON [7], _35634_[7]);
  dff (\oc8051_golden_model_1.TH0 [0], _35635_[0]);
  dff (\oc8051_golden_model_1.TH0 [1], _35635_[1]);
  dff (\oc8051_golden_model_1.TH0 [2], _35635_[2]);
  dff (\oc8051_golden_model_1.TH0 [3], _35635_[3]);
  dff (\oc8051_golden_model_1.TH0 [4], _35635_[4]);
  dff (\oc8051_golden_model_1.TH0 [5], _35635_[5]);
  dff (\oc8051_golden_model_1.TH0 [6], _35635_[6]);
  dff (\oc8051_golden_model_1.TH0 [7], _35635_[7]);
  dff (\oc8051_golden_model_1.TH1 [0], _35636_[0]);
  dff (\oc8051_golden_model_1.TH1 [1], _35636_[1]);
  dff (\oc8051_golden_model_1.TH1 [2], _35636_[2]);
  dff (\oc8051_golden_model_1.TH1 [3], _35636_[3]);
  dff (\oc8051_golden_model_1.TH1 [4], _35636_[4]);
  dff (\oc8051_golden_model_1.TH1 [5], _35636_[5]);
  dff (\oc8051_golden_model_1.TH1 [6], _35636_[6]);
  dff (\oc8051_golden_model_1.TH1 [7], _35636_[7]);
  dff (\oc8051_golden_model_1.TL0 [0], _35637_[0]);
  dff (\oc8051_golden_model_1.TL0 [1], _35637_[1]);
  dff (\oc8051_golden_model_1.TL0 [2], _35637_[2]);
  dff (\oc8051_golden_model_1.TL0 [3], _35637_[3]);
  dff (\oc8051_golden_model_1.TL0 [4], _35637_[4]);
  dff (\oc8051_golden_model_1.TL0 [5], _35637_[5]);
  dff (\oc8051_golden_model_1.TL0 [6], _35637_[6]);
  dff (\oc8051_golden_model_1.TL0 [7], _35637_[7]);
  dff (\oc8051_golden_model_1.TL1 [0], _35638_[0]);
  dff (\oc8051_golden_model_1.TL1 [1], _35638_[1]);
  dff (\oc8051_golden_model_1.TL1 [2], _35638_[2]);
  dff (\oc8051_golden_model_1.TL1 [3], _35638_[3]);
  dff (\oc8051_golden_model_1.TL1 [4], _35638_[4]);
  dff (\oc8051_golden_model_1.TL1 [5], _35638_[5]);
  dff (\oc8051_golden_model_1.TL1 [6], _35638_[6]);
  dff (\oc8051_golden_model_1.TL1 [7], _35638_[7]);
  dff (\oc8051_golden_model_1.TMOD [0], _35639_[0]);
  dff (\oc8051_golden_model_1.TMOD [1], _35639_[1]);
  dff (\oc8051_golden_model_1.TMOD [2], _35639_[2]);
  dff (\oc8051_golden_model_1.TMOD [3], _35639_[3]);
  dff (\oc8051_golden_model_1.TMOD [4], _35639_[4]);
  dff (\oc8051_golden_model_1.TMOD [5], _35639_[5]);
  dff (\oc8051_golden_model_1.TMOD [6], _35639_[6]);
  dff (\oc8051_golden_model_1.TMOD [7], _35639_[7]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [0], _35640_[0]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [1], _35640_[1]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [2], _35640_[2]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [3], _35640_[3]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [4], _35640_[4]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [5], _35640_[5]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [6], _35640_[6]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [7], _35640_[7]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [8], _35640_[8]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [9], _35640_[9]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [10], _35640_[10]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [11], _35640_[11]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [12], _35640_[12]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [13], _35640_[13]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [14], _35640_[14]);
  dff (\oc8051_golden_model_1.XRAM_ADDR [15], _35640_[15]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [0], _35642_[0]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [1], _35642_[1]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [2], _35642_[2]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [3], _35642_[3]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [4], _35642_[4]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [5], _35642_[5]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [6], _35642_[6]);
  dff (\oc8051_golden_model_1.XRAM_DATA_OUT [7], _35642_[7]);
  dff (\oc8051_golden_model_1.P0INREG [0], _35620_[0]);
  dff (\oc8051_golden_model_1.P0INREG [1], _35620_[1]);
  dff (\oc8051_golden_model_1.P0INREG [2], _35620_[2]);
  dff (\oc8051_golden_model_1.P0INREG [3], _35620_[3]);
  dff (\oc8051_golden_model_1.P0INREG [4], _35620_[4]);
  dff (\oc8051_golden_model_1.P0INREG [5], _35620_[5]);
  dff (\oc8051_golden_model_1.P0INREG [6], _35620_[6]);
  dff (\oc8051_golden_model_1.P0INREG [7], _35620_[7]);
  dff (\oc8051_golden_model_1.P1INREG [0], _35622_[0]);
  dff (\oc8051_golden_model_1.P1INREG [1], _35622_[1]);
  dff (\oc8051_golden_model_1.P1INREG [2], _35622_[2]);
  dff (\oc8051_golden_model_1.P1INREG [3], _35622_[3]);
  dff (\oc8051_golden_model_1.P1INREG [4], _35622_[4]);
  dff (\oc8051_golden_model_1.P1INREG [5], _35622_[5]);
  dff (\oc8051_golden_model_1.P1INREG [6], _35622_[6]);
  dff (\oc8051_golden_model_1.P1INREG [7], _35622_[7]);
  dff (\oc8051_golden_model_1.P2INREG [0], _35624_[0]);
  dff (\oc8051_golden_model_1.P2INREG [1], _35624_[1]);
  dff (\oc8051_golden_model_1.P2INREG [2], _35624_[2]);
  dff (\oc8051_golden_model_1.P2INREG [3], _35624_[3]);
  dff (\oc8051_golden_model_1.P2INREG [4], _35624_[4]);
  dff (\oc8051_golden_model_1.P2INREG [5], _35624_[5]);
  dff (\oc8051_golden_model_1.P2INREG [6], _35624_[6]);
  dff (\oc8051_golden_model_1.P2INREG [7], _35624_[7]);
  dff (\oc8051_golden_model_1.P3INREG [0], _35626_[0]);
  dff (\oc8051_golden_model_1.P3INREG [1], _35626_[1]);
  dff (\oc8051_golden_model_1.P3INREG [2], _35626_[2]);
  dff (\oc8051_golden_model_1.P3INREG [3], _35626_[3]);
  dff (\oc8051_golden_model_1.P3INREG [4], _35626_[4]);
  dff (\oc8051_golden_model_1.P3INREG [5], _35626_[5]);
  dff (\oc8051_golden_model_1.P3INREG [6], _35626_[6]);
  dff (\oc8051_golden_model_1.P3INREG [7], _35626_[7]);
  dff (\oc8051_golden_model_1.XRAM_DATA_IN [0], _35641_[0]);
  dff (\oc8051_golden_model_1.XRAM_DATA_IN [1], _35641_[1]);
  dff (\oc8051_golden_model_1.XRAM_DATA_IN [2], _35641_[2]);
  dff (\oc8051_golden_model_1.XRAM_DATA_IN [3], _35641_[3]);
  dff (\oc8051_golden_model_1.XRAM_DATA_IN [4], _35641_[4]);
  dff (\oc8051_golden_model_1.XRAM_DATA_IN [5], _35641_[5]);
  dff (\oc8051_golden_model_1.XRAM_DATA_IN [6], _35641_[6]);
  dff (\oc8051_golden_model_1.XRAM_DATA_IN [7], _35641_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _35772_[0]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _35772_[1]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _35772_[2]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _35772_[3]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _35772_[4]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _35772_[5]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _35771_[0]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _35771_[1]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _35773_[0]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _35773_[1]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _35773_[2]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _35773_[3]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _35773_[4]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _35773_[5]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _35773_[6]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _35773_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _35774_[0]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _35774_[1]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _35775_[0]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _35775_[1]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _35775_[2]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _35775_[3]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _35775_[4]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _35775_[5]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _35775_[6]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _35775_[7]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _35775_[8]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _35775_[9]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _35775_[10]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _35775_[11]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _35775_[12]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _35775_[13]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _35775_[14]);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _35775_[15]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _35776_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _35776_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _35776_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _35776_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _35776_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _35776_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _35776_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _35776_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _35777_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _35777_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _35777_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _35777_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _35777_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _35777_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _35777_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _35777_[7]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _35778_[0]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _35778_[1]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _35778_[2]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _35778_[3]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _35778_[4]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _35778_[5]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _35778_[6]);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _35778_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _35783_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _35784_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _35784_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _35785_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _35785_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _35786_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _35786_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _35786_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _35787_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _35787_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _35787_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _35788_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _35788_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _35789_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _35789_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _35789_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _35789_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _35790_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _35790_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _35791_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _35779_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _35779_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _35779_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _35780_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _35780_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _35780_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _35781_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _35781_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _35782_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _35782_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _35782_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _35782_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _35782_[4]);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _35782_[5]);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _35782_[6]);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _35782_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _35792_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _35793_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _35793_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _35793_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _35793_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _35793_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _35793_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _35793_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _35793_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _35793_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _35793_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _35793_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _35793_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _35793_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _35793_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _35793_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _35793_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _35794_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _35794_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _35794_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _35794_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _35794_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _35794_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _35794_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _35794_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _35794_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _35794_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _35794_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _35794_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _35794_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _35794_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _35794_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _35794_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _35817_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _35817_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _35817_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _35817_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _35817_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _35817_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _35817_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _35817_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _35817_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _35817_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _35817_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _35817_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _35817_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _35817_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _35817_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _35817_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _35817_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _35817_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _35817_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _35817_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _35817_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _35817_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _35817_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _35817_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _35817_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _35817_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _35817_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _35817_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _35817_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _35817_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _35817_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _35817_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _35795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _35796_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _35796_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _35796_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _35796_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _35796_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _35797_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _35797_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _35797_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _35797_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _35797_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _35797_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _35797_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _35797_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _35798_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _35798_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _35798_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _35798_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _35798_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _35798_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _35798_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _35798_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _35799_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _35799_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _35799_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _35799_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _35799_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _35799_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _35799_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _35799_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _35800_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _35801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _35802_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _35802_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _35802_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _35802_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _35802_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _35802_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _35802_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _35802_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _35803_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _35803_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _35803_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _35803_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _35803_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _35803_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _35803_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _35803_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _35803_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _35803_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _35803_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _35803_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _35803_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _35803_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _35803_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _35803_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _35804_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _35804_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _35804_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _35804_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _35804_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _35804_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _35804_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _35804_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _35804_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _35804_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _35804_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _35804_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _35804_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _35804_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _35804_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _35804_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _35805_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _35807_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _35806_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _35808_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _35808_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _35808_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _35808_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _35808_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _35808_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _35808_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _35808_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _35809_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _35809_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _35809_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _35810_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _35810_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _35810_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _35810_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _35810_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _35810_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _35810_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _35810_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _35811_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _35811_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _35811_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _35811_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _35811_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _35811_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _35811_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _35811_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _35812_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _35813_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _35813_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _35813_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _35813_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _35813_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _35813_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _35813_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _35813_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _35814_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _35815_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _35816_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _35816_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _35816_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _35816_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _35818_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _35818_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _35818_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _35818_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _35818_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _35818_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _35818_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _35818_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _35818_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _35818_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _35818_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _35818_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _35818_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _35818_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _35818_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _35818_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _35818_[16]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _35818_[17]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _35818_[18]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _35818_[19]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _35818_[20]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _35818_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _35818_[22]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _35818_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _35818_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _35818_[25]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _35818_[26]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _35818_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _35818_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _35818_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _35818_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _35818_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _35819_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _35819_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _35819_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _35819_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _35819_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _35819_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _35819_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _35819_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _35820_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _35821_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _35822_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _35822_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _35822_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _35822_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _35822_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _35822_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _35822_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _35822_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _35822_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _35822_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _35822_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _35822_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _35822_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _35822_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _35822_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _35822_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _35823_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _35824_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _35825_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _35826_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _35826_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _35826_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _35826_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _35826_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _35826_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _35826_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _35826_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _35826_[8]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _35826_[9]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _35826_[10]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _35826_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _35826_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _35826_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _35826_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _35826_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _35827_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _35828_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _35829_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _35829_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _35829_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _35829_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _35829_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _35829_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _35829_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _35829_[7]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _35830_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _35831_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _35831_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _35831_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _35832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _35833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _35834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _35835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _35836_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _35837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _35838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _35839_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _35944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _35945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _35946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _35947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _35948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _35949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _35950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _35951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _35888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _35889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _35890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _35891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _35892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _35893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _35894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _35895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _35936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _35937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _35938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _35939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _35940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _35941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _35942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _35943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _35928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _35929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _35930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _35931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _35932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _35933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _35934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _35935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _35920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _35921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _35922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _35923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _35924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _35925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _35926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _35927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _35912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _35913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _35914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _35915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _35916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _35917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _35918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _35919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _35904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _35905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _35906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _35907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _35908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _35909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _35910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _35911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _35896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _35897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _35898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _35899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _35900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _35901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _35902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _35903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _35952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _35953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _35954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _35955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _35956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _35957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _35958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _35959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _35872_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _35873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _35874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _35875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _35876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _35877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _35878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _35879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _35864_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _35865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _35866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _35867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _35868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _35869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _35870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _35871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _35856_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _35857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _35858_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _35859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _35860_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _35861_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _35862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _35863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _35848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _35849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _35850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _35851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _35852_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _35853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _35854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _35855_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _35840_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _35841_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _35842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _35843_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _35844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _35845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _35846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _35847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _35880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _35881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _35882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _35883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _35884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _35885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _35886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _35887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _35960_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _35960_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _35960_[2]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _35960_[3]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _35960_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _35960_[5]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _35960_[6]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _35960_[7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _35961_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _35962_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _35963_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _35963_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _35963_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _35963_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _35963_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _35963_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _35963_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _35963_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _35964_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _35965_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _35965_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _35965_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _35965_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _35965_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _35965_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _35965_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _35965_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _35966_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _35966_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _35966_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _35966_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _35966_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _35966_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _35966_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _35966_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _35967_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _35967_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _35967_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _35967_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _35967_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _35967_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _35967_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _35967_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _35968_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _35968_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _35968_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _35968_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _35968_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _35968_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _35968_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _35968_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _35969_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _35969_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _35969_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _35969_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _35969_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _35969_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _35969_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _35969_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _35970_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _35970_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _35970_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _35970_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _35970_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _35970_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _35970_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _35970_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _35971_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _35971_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _35971_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _35971_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _35971_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _35971_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _35971_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _35971_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _35972_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _35972_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _35972_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _35972_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _35972_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _35972_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _35972_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _35972_[7]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _35973_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _35973_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _35973_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _35973_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _35973_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _35973_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _35973_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _35974_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _35975_[0]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _35975_[1]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _35975_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _35975_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _35975_[4]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _35975_[5]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _35975_[6]);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _35975_[7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [1], \oc8051_top_1.oc8051_sfr1.psw_next [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [2], \oc8051_top_1.oc8051_sfr1.psw_next [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [3], \oc8051_top_1.oc8051_sfr1.psw_next [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [4], \oc8051_top_1.oc8051_sfr1.psw_next [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [5], \oc8051_top_1.oc8051_sfr1.psw_next [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [6], \oc8051_top_1.oc8051_sfr1.psw_next [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.psw_next_i [7], \oc8051_top_1.oc8051_sfr1.psw_next [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw_impl[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_next [0], psw_impl[0]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.SBUF_next [0], \oc8051_golden_model_1.SBUF [0]);
  buf(\oc8051_golden_model_1.SBUF_next [1], \oc8051_golden_model_1.SBUF [1]);
  buf(\oc8051_golden_model_1.SBUF_next [2], \oc8051_golden_model_1.SBUF [2]);
  buf(\oc8051_golden_model_1.SBUF_next [3], \oc8051_golden_model_1.SBUF [3]);
  buf(\oc8051_golden_model_1.SBUF_next [4], \oc8051_golden_model_1.SBUF [4]);
  buf(\oc8051_golden_model_1.SBUF_next [5], \oc8051_golden_model_1.SBUF [5]);
  buf(\oc8051_golden_model_1.SBUF_next [6], \oc8051_golden_model_1.SBUF [6]);
  buf(\oc8051_golden_model_1.SBUF_next [7], \oc8051_golden_model_1.SBUF [7]);
  buf(\oc8051_golden_model_1.SCON_next [0], \oc8051_golden_model_1.SCON [0]);
  buf(\oc8051_golden_model_1.SCON_next [1], \oc8051_golden_model_1.SCON [1]);
  buf(\oc8051_golden_model_1.SCON_next [2], \oc8051_golden_model_1.SCON [2]);
  buf(\oc8051_golden_model_1.SCON_next [3], \oc8051_golden_model_1.SCON [3]);
  buf(\oc8051_golden_model_1.SCON_next [4], \oc8051_golden_model_1.SCON [4]);
  buf(\oc8051_golden_model_1.SCON_next [5], \oc8051_golden_model_1.SCON [5]);
  buf(\oc8051_golden_model_1.SCON_next [6], \oc8051_golden_model_1.SCON [6]);
  buf(\oc8051_golden_model_1.SCON_next [7], \oc8051_golden_model_1.SCON [7]);
  buf(\oc8051_golden_model_1.PCON_next [0], \oc8051_golden_model_1.PCON [0]);
  buf(\oc8051_golden_model_1.PCON_next [1], \oc8051_golden_model_1.PCON [1]);
  buf(\oc8051_golden_model_1.PCON_next [2], \oc8051_golden_model_1.PCON [2]);
  buf(\oc8051_golden_model_1.PCON_next [3], \oc8051_golden_model_1.PCON [3]);
  buf(\oc8051_golden_model_1.PCON_next [4], \oc8051_golden_model_1.PCON [4]);
  buf(\oc8051_golden_model_1.PCON_next [5], \oc8051_golden_model_1.PCON [5]);
  buf(\oc8051_golden_model_1.PCON_next [6], \oc8051_golden_model_1.PCON [6]);
  buf(\oc8051_golden_model_1.PCON_next [7], \oc8051_golden_model_1.PCON [7]);
  buf(\oc8051_golden_model_1.TCON_next [0], \oc8051_golden_model_1.TCON [0]);
  buf(\oc8051_golden_model_1.TCON_next [1], \oc8051_golden_model_1.TCON [1]);
  buf(\oc8051_golden_model_1.TCON_next [2], \oc8051_golden_model_1.TCON [2]);
  buf(\oc8051_golden_model_1.TCON_next [3], \oc8051_golden_model_1.TCON [3]);
  buf(\oc8051_golden_model_1.TCON_next [4], \oc8051_golden_model_1.TCON [4]);
  buf(\oc8051_golden_model_1.TCON_next [5], \oc8051_golden_model_1.TCON [5]);
  buf(\oc8051_golden_model_1.TCON_next [6], \oc8051_golden_model_1.TCON [6]);
  buf(\oc8051_golden_model_1.TCON_next [7], \oc8051_golden_model_1.TCON [7]);
  buf(\oc8051_golden_model_1.TL0_next [0], \oc8051_golden_model_1.TL0 [0]);
  buf(\oc8051_golden_model_1.TL0_next [1], \oc8051_golden_model_1.TL0 [1]);
  buf(\oc8051_golden_model_1.TL0_next [2], \oc8051_golden_model_1.TL0 [2]);
  buf(\oc8051_golden_model_1.TL0_next [3], \oc8051_golden_model_1.TL0 [3]);
  buf(\oc8051_golden_model_1.TL0_next [4], \oc8051_golden_model_1.TL0 [4]);
  buf(\oc8051_golden_model_1.TL0_next [5], \oc8051_golden_model_1.TL0 [5]);
  buf(\oc8051_golden_model_1.TL0_next [6], \oc8051_golden_model_1.TL0 [6]);
  buf(\oc8051_golden_model_1.TL0_next [7], \oc8051_golden_model_1.TL0 [7]);
  buf(\oc8051_golden_model_1.TL1_next [0], \oc8051_golden_model_1.TL1 [0]);
  buf(\oc8051_golden_model_1.TL1_next [1], \oc8051_golden_model_1.TL1 [1]);
  buf(\oc8051_golden_model_1.TL1_next [2], \oc8051_golden_model_1.TL1 [2]);
  buf(\oc8051_golden_model_1.TL1_next [3], \oc8051_golden_model_1.TL1 [3]);
  buf(\oc8051_golden_model_1.TL1_next [4], \oc8051_golden_model_1.TL1 [4]);
  buf(\oc8051_golden_model_1.TL1_next [5], \oc8051_golden_model_1.TL1 [5]);
  buf(\oc8051_golden_model_1.TL1_next [6], \oc8051_golden_model_1.TL1 [6]);
  buf(\oc8051_golden_model_1.TL1_next [7], \oc8051_golden_model_1.TL1 [7]);
  buf(\oc8051_golden_model_1.TH0_next [0], \oc8051_golden_model_1.TH0 [0]);
  buf(\oc8051_golden_model_1.TH0_next [1], \oc8051_golden_model_1.TH0 [1]);
  buf(\oc8051_golden_model_1.TH0_next [2], \oc8051_golden_model_1.TH0 [2]);
  buf(\oc8051_golden_model_1.TH0_next [3], \oc8051_golden_model_1.TH0 [3]);
  buf(\oc8051_golden_model_1.TH0_next [4], \oc8051_golden_model_1.TH0 [4]);
  buf(\oc8051_golden_model_1.TH0_next [5], \oc8051_golden_model_1.TH0 [5]);
  buf(\oc8051_golden_model_1.TH0_next [6], \oc8051_golden_model_1.TH0 [6]);
  buf(\oc8051_golden_model_1.TH0_next [7], \oc8051_golden_model_1.TH0 [7]);
  buf(\oc8051_golden_model_1.TH1_next [0], \oc8051_golden_model_1.TH1 [0]);
  buf(\oc8051_golden_model_1.TH1_next [1], \oc8051_golden_model_1.TH1 [1]);
  buf(\oc8051_golden_model_1.TH1_next [2], \oc8051_golden_model_1.TH1 [2]);
  buf(\oc8051_golden_model_1.TH1_next [3], \oc8051_golden_model_1.TH1 [3]);
  buf(\oc8051_golden_model_1.TH1_next [4], \oc8051_golden_model_1.TH1 [4]);
  buf(\oc8051_golden_model_1.TH1_next [5], \oc8051_golden_model_1.TH1 [5]);
  buf(\oc8051_golden_model_1.TH1_next [6], \oc8051_golden_model_1.TH1 [6]);
  buf(\oc8051_golden_model_1.TH1_next [7], \oc8051_golden_model_1.TH1 [7]);
  buf(\oc8051_golden_model_1.TMOD_next [0], \oc8051_golden_model_1.TMOD [0]);
  buf(\oc8051_golden_model_1.TMOD_next [1], \oc8051_golden_model_1.TMOD [1]);
  buf(\oc8051_golden_model_1.TMOD_next [2], \oc8051_golden_model_1.TMOD [2]);
  buf(\oc8051_golden_model_1.TMOD_next [3], \oc8051_golden_model_1.TMOD [3]);
  buf(\oc8051_golden_model_1.TMOD_next [4], \oc8051_golden_model_1.TMOD [4]);
  buf(\oc8051_golden_model_1.TMOD_next [5], \oc8051_golden_model_1.TMOD [5]);
  buf(\oc8051_golden_model_1.TMOD_next [6], \oc8051_golden_model_1.TMOD [6]);
  buf(\oc8051_golden_model_1.TMOD_next [7], \oc8051_golden_model_1.TMOD [7]);
  buf(\oc8051_golden_model_1.IE_next [0], \oc8051_golden_model_1.IE [0]);
  buf(\oc8051_golden_model_1.IE_next [1], \oc8051_golden_model_1.IE [1]);
  buf(\oc8051_golden_model_1.IE_next [2], \oc8051_golden_model_1.IE [2]);
  buf(\oc8051_golden_model_1.IE_next [3], \oc8051_golden_model_1.IE [3]);
  buf(\oc8051_golden_model_1.IE_next [4], \oc8051_golden_model_1.IE [4]);
  buf(\oc8051_golden_model_1.IE_next [5], \oc8051_golden_model_1.IE [5]);
  buf(\oc8051_golden_model_1.IE_next [6], \oc8051_golden_model_1.IE [6]);
  buf(\oc8051_golden_model_1.IE_next [7], \oc8051_golden_model_1.IE [7]);
  buf(\oc8051_golden_model_1.IP_next [0], \oc8051_golden_model_1.IP [0]);
  buf(\oc8051_golden_model_1.IP_next [1], \oc8051_golden_model_1.IP [1]);
  buf(\oc8051_golden_model_1.IP_next [2], \oc8051_golden_model_1.IP [2]);
  buf(\oc8051_golden_model_1.IP_next [3], \oc8051_golden_model_1.IP [3]);
  buf(\oc8051_golden_model_1.IP_next [4], \oc8051_golden_model_1.IP [4]);
  buf(\oc8051_golden_model_1.IP_next [5], \oc8051_golden_model_1.IP [5]);
  buf(\oc8051_golden_model_1.IP_next [6], \oc8051_golden_model_1.IP [6]);
  buf(\oc8051_golden_model_1.IP_next [7], \oc8051_golden_model_1.IP [7]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e0 [0], \oc8051_golden_model_1.XRAM_DATA_IN [0]);
  buf(\oc8051_golden_model_1.ACC_e0 [1], \oc8051_golden_model_1.XRAM_DATA_IN [1]);
  buf(\oc8051_golden_model_1.ACC_e0 [2], \oc8051_golden_model_1.XRAM_DATA_IN [2]);
  buf(\oc8051_golden_model_1.ACC_e0 [3], \oc8051_golden_model_1.XRAM_DATA_IN [3]);
  buf(\oc8051_golden_model_1.ACC_e0 [4], \oc8051_golden_model_1.XRAM_DATA_IN [4]);
  buf(\oc8051_golden_model_1.ACC_e0 [5], \oc8051_golden_model_1.XRAM_DATA_IN [5]);
  buf(\oc8051_golden_model_1.ACC_e0 [6], \oc8051_golden_model_1.XRAM_DATA_IN [6]);
  buf(\oc8051_golden_model_1.ACC_e0 [7], \oc8051_golden_model_1.XRAM_DATA_IN [7]);
  buf(\oc8051_golden_model_1.ACC_e2 [0], \oc8051_golden_model_1.XRAM_DATA_IN [0]);
  buf(\oc8051_golden_model_1.ACC_e2 [1], \oc8051_golden_model_1.XRAM_DATA_IN [1]);
  buf(\oc8051_golden_model_1.ACC_e2 [2], \oc8051_golden_model_1.XRAM_DATA_IN [2]);
  buf(\oc8051_golden_model_1.ACC_e2 [3], \oc8051_golden_model_1.XRAM_DATA_IN [3]);
  buf(\oc8051_golden_model_1.ACC_e2 [4], \oc8051_golden_model_1.XRAM_DATA_IN [4]);
  buf(\oc8051_golden_model_1.ACC_e2 [5], \oc8051_golden_model_1.XRAM_DATA_IN [5]);
  buf(\oc8051_golden_model_1.ACC_e2 [6], \oc8051_golden_model_1.XRAM_DATA_IN [6]);
  buf(\oc8051_golden_model_1.ACC_e2 [7], \oc8051_golden_model_1.XRAM_DATA_IN [7]);
  buf(\oc8051_golden_model_1.ACC_e3 [0], \oc8051_golden_model_1.XRAM_DATA_IN [0]);
  buf(\oc8051_golden_model_1.ACC_e3 [1], \oc8051_golden_model_1.XRAM_DATA_IN [1]);
  buf(\oc8051_golden_model_1.ACC_e3 [2], \oc8051_golden_model_1.XRAM_DATA_IN [2]);
  buf(\oc8051_golden_model_1.ACC_e3 [3], \oc8051_golden_model_1.XRAM_DATA_IN [3]);
  buf(\oc8051_golden_model_1.ACC_e3 [4], \oc8051_golden_model_1.XRAM_DATA_IN [4]);
  buf(\oc8051_golden_model_1.ACC_e3 [5], \oc8051_golden_model_1.XRAM_DATA_IN [5]);
  buf(\oc8051_golden_model_1.ACC_e3 [6], \oc8051_golden_model_1.XRAM_DATA_IN [6]);
  buf(\oc8051_golden_model_1.ACC_e3 [7], \oc8051_golden_model_1.XRAM_DATA_IN [7]);
  buf(\oc8051_golden_model_1.ACC_e6 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.ACC_e6 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.ACC_e6 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.ACC_e6 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.ACC_e6 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.ACC_e6 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.ACC_e6 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.ACC_e6 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.ACC_e7 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.ACC_e7 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.ACC_e7 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.ACC_e7 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.ACC_e7 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.ACC_e7 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.ACC_e7 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.ACC_e7 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.PSW_00 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_00 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_00 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_00 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_00 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_00 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_00 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_00 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_01 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_01 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_01 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_01 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_01 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_01 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_01 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_01 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_02 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_02 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_02 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_02 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_02 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_02 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_02 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_02 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_03 [0], \oc8051_golden_model_1.n1041 [0]);
  buf(\oc8051_golden_model_1.PSW_03 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_03 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_03 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_03 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_03 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_03 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_03 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_04 [0], \oc8051_golden_model_1.n1058 [0]);
  buf(\oc8051_golden_model_1.PSW_04 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_04 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_04 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_04 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_04 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_04 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_04 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_06 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_06 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_06 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_06 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_06 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_06 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_06 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_06 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_07 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_07 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_07 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_07 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_07 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_07 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_07 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_07 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_08 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_08 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_08 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_08 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_08 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_08 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_08 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_08 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_09 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_09 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_09 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_09 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_09 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_09 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_09 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_09 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0a [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0b [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0c [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0d [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0e [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_0f [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_0f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_0f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_0f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_0f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_0f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_0f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_0f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_11 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_11 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_11 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_11 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_11 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_11 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_11 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_11 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_12 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_12 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_12 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_12 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_12 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_12 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_12 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_12 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.n1262 [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_14 [0], \oc8051_golden_model_1.n1279 [0]);
  buf(\oc8051_golden_model_1.PSW_14 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_14 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_14 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_14 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_14 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_14 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_14 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_16 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_16 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_16 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_16 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_16 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_16 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_16 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_16 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_17 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_17 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_17 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_17 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_17 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_17 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_17 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_17 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_18 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_18 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_18 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_18 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_18 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_18 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_18 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_18 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_19 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_19 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_19 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_19 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_19 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_19 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_19 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_19 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1a [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1b [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1c [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1d [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1e [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_1f [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_1f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_1f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_1f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_1f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_1f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_1f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_1f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_20 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_20 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_20 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_20 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_20 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_20 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_20 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_20 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_21 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_21 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_21 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_21 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_21 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_21 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_21 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_21 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_22 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_22 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_22 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_22 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_22 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_22 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_22 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_22 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_23 [0], \oc8051_golden_model_1.n1328 [0]);
  buf(\oc8051_golden_model_1.PSW_23 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_23 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_23 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_23 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_23 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_23 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_23 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.n1369 [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1369 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1369 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1369 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.n1425 [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1425 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1425 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1425 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.n1474 [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1461 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1461 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.n1474 [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1474 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1474 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.PSW_30 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_30 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_30 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_30 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_30 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_30 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_30 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_30 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_31 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_31 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_31 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_31 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_31 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_31 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_31 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_31 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_32 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_32 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_32 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_32 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_32 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_32 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_32 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_32 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.n1551 [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1587 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1587 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1587 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.n1620 [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1620 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1620 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1620 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.n1653 [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1653 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.n1653 [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1653 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.PSW_40 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_40 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_40 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_40 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_40 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_40 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_40 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_40 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_41 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_41 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_41 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_41 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_41 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_41 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_41 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_41 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_42 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_42 [1], \oc8051_golden_model_1.n1702 [1]);
  buf(\oc8051_golden_model_1.PSW_42 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.PSW_42 [3], \oc8051_golden_model_1.n1702 [3]);
  buf(\oc8051_golden_model_1.PSW_42 [4], \oc8051_golden_model_1.n1702 [4]);
  buf(\oc8051_golden_model_1.PSW_42 [5], \oc8051_golden_model_1.n1702 [5]);
  buf(\oc8051_golden_model_1.PSW_42 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.PSW_42 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.PSW_44 [0], \oc8051_golden_model_1.n1747 [0]);
  buf(\oc8051_golden_model_1.PSW_44 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_44 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_44 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_44 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_44 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_44 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_44 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_45 [0], \oc8051_golden_model_1.n1764 [0]);
  buf(\oc8051_golden_model_1.PSW_45 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_45 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_45 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_45 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_45 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_45 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_45 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_46 [0], \oc8051_golden_model_1.n1781 [0]);
  buf(\oc8051_golden_model_1.PSW_46 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_46 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_46 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_46 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_46 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_46 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_46 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_47 [0], \oc8051_golden_model_1.n1781 [0]);
  buf(\oc8051_golden_model_1.PSW_47 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_47 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_47 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_47 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_47 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_47 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_47 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_48 [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_48 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_48 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_48 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_48 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_48 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_48 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_48 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_49 [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_49 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_49 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_49 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_49 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_49 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_49 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_49 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4a [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4b [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4c [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4d [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4e [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_4f [0], \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.PSW_4f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_4f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_4f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_4f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_4f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_4f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_4f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_50 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_50 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_50 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_50 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_50 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_50 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_50 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_50 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_51 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_51 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_51 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_51 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_51 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_51 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_51 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_51 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_52 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_52 [1], \oc8051_golden_model_1.n1812 [1]);
  buf(\oc8051_golden_model_1.PSW_52 [2], \oc8051_golden_model_1.n1812 [2]);
  buf(\oc8051_golden_model_1.PSW_52 [3], \oc8051_golden_model_1.n1812 [3]);
  buf(\oc8051_golden_model_1.PSW_52 [4], \oc8051_golden_model_1.n1812 [4]);
  buf(\oc8051_golden_model_1.PSW_52 [5], \oc8051_golden_model_1.n1812 [5]);
  buf(\oc8051_golden_model_1.PSW_52 [6], \oc8051_golden_model_1.n1812 [6]);
  buf(\oc8051_golden_model_1.PSW_52 [7], \oc8051_golden_model_1.n1812 [7]);
  buf(\oc8051_golden_model_1.PSW_54 [0], \oc8051_golden_model_1.n1857 [0]);
  buf(\oc8051_golden_model_1.PSW_54 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_54 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_54 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_54 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_54 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_54 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_54 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_55 [0], \oc8051_golden_model_1.n1874 [0]);
  buf(\oc8051_golden_model_1.PSW_55 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_55 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_55 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_55 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_55 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_55 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_55 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_56 [0], \oc8051_golden_model_1.n1891 [0]);
  buf(\oc8051_golden_model_1.PSW_56 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_56 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_56 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_56 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_56 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_56 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_56 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_57 [0], \oc8051_golden_model_1.n1891 [0]);
  buf(\oc8051_golden_model_1.PSW_57 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_57 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_57 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_57 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_57 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_57 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_57 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_58 [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_58 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_58 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_58 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_58 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_58 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_58 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_58 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_59 [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_59 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_59 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_59 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_59 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_59 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_59 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_59 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5a [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5b [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5c [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5d [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5e [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_5f [0], \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.PSW_5f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_5f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_5f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_5f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_5f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_5f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_5f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_60 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_60 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_60 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_60 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_60 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_60 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_60 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_60 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_61 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_61 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_61 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_61 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_61 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_61 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_61 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_61 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_64 [0], \oc8051_golden_model_1.n1984 [0]);
  buf(\oc8051_golden_model_1.PSW_64 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_64 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_64 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_64 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_64 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_64 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_64 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_65 [0], \oc8051_golden_model_1.n2001 [0]);
  buf(\oc8051_golden_model_1.PSW_65 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_65 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_65 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_65 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_65 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_65 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_65 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_66 [0], \oc8051_golden_model_1.n2018 [0]);
  buf(\oc8051_golden_model_1.PSW_66 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_66 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_66 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_66 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_66 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_66 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_66 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_67 [0], \oc8051_golden_model_1.n2018 [0]);
  buf(\oc8051_golden_model_1.PSW_67 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_67 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_67 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_67 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_67 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_67 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_67 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_68 [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_68 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_68 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_68 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_68 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_68 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_68 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_68 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_69 [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_69 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_69 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_69 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_69 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_69 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_69 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_69 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6a [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6b [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6c [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6d [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6e [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_6f [0], \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.PSW_6f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_6f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_6f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_6f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_6f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_6f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_6f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_70 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_70 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_70 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_70 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_70 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_70 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_70 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_70 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_71 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_71 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_71 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_71 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_71 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_71 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_71 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_71 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n2043 [7]);
  buf(\oc8051_golden_model_1.PSW_73 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_73 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_73 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_73 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_73 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_73 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_73 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_73 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_74 [0], \oc8051_golden_model_1.n2059 [0]);
  buf(\oc8051_golden_model_1.PSW_74 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_74 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_74 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_74 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_74 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_74 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_74 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_76 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_76 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_76 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_76 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_76 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_76 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_76 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_76 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_77 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_77 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_77 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_77 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_77 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_77 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_77 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_77 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_78 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_78 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_78 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_78 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_78 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_78 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_78 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_78 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_79 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_79 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_79 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_79 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_79 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_79 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_79 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_79 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7a [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7a [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7a [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7a [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7b [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7b [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7b [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7b [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7c [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7c [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7c [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7c [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7d [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7d [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7d [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7d [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7e [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7e [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7e [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7e [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_7f [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_7f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_7f [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_7f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_7f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_7f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_7f [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_7f [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_80 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_80 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_80 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_80 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_80 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_80 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_80 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_80 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_81 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_81 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_81 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_81 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_81 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_81 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_81 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_81 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n2090 [7]);
  buf(\oc8051_golden_model_1.PSW_83 [0], \oc8051_golden_model_1.n2059 [0]);
  buf(\oc8051_golden_model_1.PSW_83 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_83 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_83 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_83 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_83 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_83 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_83 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.n2116 [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n2116 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_90 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_90 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_90 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_90 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_90 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_90 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_90 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_90 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_91 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_91 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_91 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_91 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_91 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_91 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_91 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_91 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_93 [0], \oc8051_golden_model_1.n2059 [0]);
  buf(\oc8051_golden_model_1.PSW_93 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_93 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_93 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_93 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_93 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_93 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_93 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.n2302 [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n2302 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n2302 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n2302 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.n2332 [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n2332 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n2332 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n2332 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.n2362 [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n2362 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n2362 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n2362 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.n2362 [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n2362 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n2362 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n2362 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n2397 [7]);
  buf(\oc8051_golden_model_1.PSW_a1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n2400 [7]);
  buf(\oc8051_golden_model_1.PSW_a3 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.n2428 [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n2428 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_a5 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a6 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a7 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a8 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_a9 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_a9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_aa [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_aa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_aa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_aa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_aa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_aa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_aa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_aa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ab [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ab [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ab [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ab [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ab [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ab [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ab [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ab [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ac [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ac [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ac [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ac [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ac [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ac [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ac [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ac [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ad [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ad [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ad [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ad [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ad [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ad [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ad [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ad [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ae [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ae [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ae [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ae [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ae [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ae [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ae [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ae [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_af [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_af [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_af [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_af [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_af [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_af [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_af [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_af [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n2433 [7]);
  buf(\oc8051_golden_model_1.PSW_b1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n2464 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n2472 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n2488 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n2488 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.PSW_c0 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_c0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_c1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_c4 [0], \oc8051_golden_model_1.n2537 [0]);
  buf(\oc8051_golden_model_1.PSW_c4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c6 [0], \oc8051_golden_model_1.n2579 [0]);
  buf(\oc8051_golden_model_1.PSW_c6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c7 [0], \oc8051_golden_model_1.n2579 [0]);
  buf(\oc8051_golden_model_1.PSW_c7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c8 [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_c8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_c9 [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_c9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ca [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ca [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ca [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ca [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ca [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ca [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ca [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ca [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cb [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_cb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cc [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_cc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cd [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_cd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ce [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ce [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ce [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ce [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ce [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ce [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ce [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ce [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_cf [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_cf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_cf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_cf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_cf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_cf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_cf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_cf [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_d1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.n2664 [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n2664 [7]);
  buf(\oc8051_golden_model_1.PSW_d6 [0], \oc8051_golden_model_1.n2686 [0]);
  buf(\oc8051_golden_model_1.PSW_d6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d7 [0], \oc8051_golden_model_1.n2686 [0]);
  buf(\oc8051_golden_model_1.PSW_d7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d8 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_d8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_d9 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_d9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_da [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_da [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_da [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_da [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_da [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_da [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_da [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_da [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_db [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_db [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_db [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_db [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_db [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_db [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_db [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_db [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dc [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_dc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_dd [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_dd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_dd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_dd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_dd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_dd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_dd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_dd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_de [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_de [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_de [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_de [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_de [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_de [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_de [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_de [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_df [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_df [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_df [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_df [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_df [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_df [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_df [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_df [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e0 [0], \oc8051_golden_model_1.n2705 [0]);
  buf(\oc8051_golden_model_1.PSW_e0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_e1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e2 [0], \oc8051_golden_model_1.n2705 [0]);
  buf(\oc8051_golden_model_1.PSW_e2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e2 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e3 [0], \oc8051_golden_model_1.n2705 [0]);
  buf(\oc8051_golden_model_1.PSW_e3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e4 [0], \oc8051_golden_model_1.n2722 [0]);
  buf(\oc8051_golden_model_1.PSW_e4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e5 [0], \oc8051_golden_model_1.n2723 [0]);
  buf(\oc8051_golden_model_1.PSW_e5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e5 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e6 [0], \oc8051_golden_model_1.n2579 [0]);
  buf(\oc8051_golden_model_1.PSW_e6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e7 [0], \oc8051_golden_model_1.n2579 [0]);
  buf(\oc8051_golden_model_1.PSW_e7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e8 [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_e8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_e9 [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_e9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_e9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_e9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_e9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_e9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_e9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_e9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ea [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ea [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ea [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ea [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ea [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ea [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ea [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ea [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_eb [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_eb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_eb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_eb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_eb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_eb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_eb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_eb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ec [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ec [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ec [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ec [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ec [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ec [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ec [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ec [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ed [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ed [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ed [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ed [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ed [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ed [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ed [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ed [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ee [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ee [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ee [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ee [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ee [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ee [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ee [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ee [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ef [0], \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.PSW_ef [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ef [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ef [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ef [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ef [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ef [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ef [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f0 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f0 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f1 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f1 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f1 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f1 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f1 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f1 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f1 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f1 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f2 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f2 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f3 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f3 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f4 [0], \oc8051_golden_model_1.n2740 [0]);
  buf(\oc8051_golden_model_1.PSW_f4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f4 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f5 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f5 [1], \oc8051_golden_model_1.n2741 [1]);
  buf(\oc8051_golden_model_1.PSW_f5 [2], \oc8051_golden_model_1.n2741 [2]);
  buf(\oc8051_golden_model_1.PSW_f5 [3], \oc8051_golden_model_1.n2741 [3]);
  buf(\oc8051_golden_model_1.PSW_f5 [4], \oc8051_golden_model_1.n2741 [4]);
  buf(\oc8051_golden_model_1.PSW_f5 [5], \oc8051_golden_model_1.n2741 [5]);
  buf(\oc8051_golden_model_1.PSW_f5 [6], \oc8051_golden_model_1.n2741 [6]);
  buf(\oc8051_golden_model_1.PSW_f5 [7], \oc8051_golden_model_1.n2741 [7]);
  buf(\oc8051_golden_model_1.PSW_f6 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f6 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f7 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f7 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f8 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f8 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_f9 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_f9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_f9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_f9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_f9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_f9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_f9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_f9 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fa [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_fa [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fa [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fa [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fa [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fa [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fa [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fa [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fb [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_fb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fb [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fc [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_fc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fc [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fd [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_fd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fd [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_fe [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_fe [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_fe [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_fe [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_fe [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_fe [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_fe [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_fe [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.PSW_ff [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.PSW_ff [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ff [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ff [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ff [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ff [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ff [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ff [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e0 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [8], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [9], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [10], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [11], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [12], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [13], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [14], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e2 [15], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [8], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [9], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [10], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [11], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [12], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [13], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [14], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_e3 [15], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f0 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [8], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [9], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [10], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [11], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [12], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [13], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [14], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f2 [15], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [8], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [9], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [10], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [11], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [12], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [13], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [14], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_ADDR_f3 [15], 1'b0);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f0 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f2 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.XRAM_DATA_OUT_f3 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0573 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n0573 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n0573 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n0573 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n0573 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.n0573 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.n0573 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.n0573 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n0606 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n0606 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n0606 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n0606 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n0606 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n0606 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n0606 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n0606 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n0713 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0713 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0713 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0713 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0713 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0713 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0713 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0713 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0713 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0713 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0745 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0745 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0745 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0745 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0745 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0745 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0745 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0745 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0745 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0745 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0745 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0745 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0745 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0745 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0745 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0745 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n1002 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1002 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1002 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1002 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1002 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1002 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1002 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1003 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1004 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1005 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1006 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1007 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1008 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1009 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1010 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1017 , \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n1018 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n1018 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1018 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1018 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1018 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1018 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1018 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1018 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1025 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1025 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1025 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1025 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1025 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1025 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1025 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1025 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1026 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1027 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1028 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1029 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1030 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1031 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1032 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1033 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1040 , \oc8051_golden_model_1.n1041 [0]);
  buf(\oc8051_golden_model_1.n1041 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1041 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1041 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1041 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1041 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1041 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1041 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1057 , \oc8051_golden_model_1.n1058 [0]);
  buf(\oc8051_golden_model_1.n1058 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1058 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1058 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1058 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1058 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1058 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1058 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1139 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n1139 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n1139 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n1139 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n1141 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1141 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1143 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1143 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1143 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1143 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1144 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1144 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1144 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1145 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1145 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1145 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1146 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1146 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1146 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1146 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1147 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1147 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1148 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1148 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1148 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1148 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1149 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1149 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1149 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1149 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1195 , \oc8051_golden_model_1.n2400 [7]);
  buf(\oc8051_golden_model_1.n1237 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1238 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1238 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1238 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1238 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1238 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1238 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1238 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1238 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1238 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1239 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1239 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1239 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1239 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1239 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1239 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1239 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1239 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1239 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1240 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1240 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1240 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1240 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1240 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1240 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1240 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1240 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1241 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1242 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1242 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1242 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1243 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1244 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1244 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1245 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1245 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1245 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1245 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1245 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1245 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1245 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1245 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1246 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1246 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1246 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1246 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1246 [6], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1247 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1248 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1249 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1251 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1252 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1253 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1254 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1261 , \oc8051_golden_model_1.n1262 [0]);
  buf(\oc8051_golden_model_1.n1262 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1262 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1262 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1262 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1262 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1262 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1262 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1278 , \oc8051_golden_model_1.n1279 [0]);
  buf(\oc8051_golden_model_1.n1279 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1279 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1279 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1279 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1279 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1279 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1279 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1310 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n1310 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n1310 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n1310 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n1310 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n1310 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n1310 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n1310 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n1310 [8], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n1310 [9], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n1310 [10], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n1310 [11], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n1310 [12], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.n1310 [13], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.n1310 [14], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.n1310 [15], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n1312 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1312 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1312 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1312 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1312 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1312 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1312 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1312 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1313 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1314 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1315 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1316 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1317 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1318 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1319 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1320 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1327 , \oc8051_golden_model_1.n1328 [0]);
  buf(\oc8051_golden_model_1.n1328 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1328 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1328 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1328 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1328 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1328 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1328 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1330 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1330 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1330 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1330 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1330 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1330 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1330 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1330 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1330 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1334 [8], \oc8051_golden_model_1.n1369 [7]);
  buf(\oc8051_golden_model_1.n1335 , \oc8051_golden_model_1.n1369 [7]);
  buf(\oc8051_golden_model_1.n1336 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1336 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1336 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1336 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1337 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1337 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1337 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1337 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1337 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.n1369 [6]);
  buf(\oc8051_golden_model_1.n1342 , \oc8051_golden_model_1.n1369 [6]);
  buf(\oc8051_golden_model_1.n1343 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1343 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1343 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1343 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1343 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1343 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1343 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1343 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1343 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1351 , \oc8051_golden_model_1.n1369 [2]);
  buf(\oc8051_golden_model_1.n1352 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1352 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1352 [2], \oc8051_golden_model_1.n1369 [2]);
  buf(\oc8051_golden_model_1.n1352 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1352 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1352 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1352 [6], \oc8051_golden_model_1.n1369 [6]);
  buf(\oc8051_golden_model_1.n1352 [7], \oc8051_golden_model_1.n1369 [7]);
  buf(\oc8051_golden_model_1.n1353 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1353 [1], \oc8051_golden_model_1.n1369 [2]);
  buf(\oc8051_golden_model_1.n1353 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1353 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1353 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1353 [5], \oc8051_golden_model_1.n1369 [6]);
  buf(\oc8051_golden_model_1.n1353 [6], \oc8051_golden_model_1.n1369 [7]);
  buf(\oc8051_golden_model_1.n1368 , \oc8051_golden_model_1.n1369 [0]);
  buf(\oc8051_golden_model_1.n1369 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1369 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1369 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1369 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1392 [8], \oc8051_golden_model_1.n1425 [7]);
  buf(\oc8051_golden_model_1.n1393 , \oc8051_golden_model_1.n1425 [7]);
  buf(\oc8051_golden_model_1.n1398 [4], \oc8051_golden_model_1.n1425 [6]);
  buf(\oc8051_golden_model_1.n1399 , \oc8051_golden_model_1.n1425 [6]);
  buf(\oc8051_golden_model_1.n1407 , \oc8051_golden_model_1.n1425 [2]);
  buf(\oc8051_golden_model_1.n1408 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1408 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1408 [2], \oc8051_golden_model_1.n1425 [2]);
  buf(\oc8051_golden_model_1.n1408 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1408 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1408 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1408 [6], \oc8051_golden_model_1.n1425 [6]);
  buf(\oc8051_golden_model_1.n1408 [7], \oc8051_golden_model_1.n1425 [7]);
  buf(\oc8051_golden_model_1.n1409 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1409 [1], \oc8051_golden_model_1.n1425 [2]);
  buf(\oc8051_golden_model_1.n1409 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1409 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1409 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1409 [5], \oc8051_golden_model_1.n1425 [6]);
  buf(\oc8051_golden_model_1.n1409 [6], \oc8051_golden_model_1.n1425 [7]);
  buf(\oc8051_golden_model_1.n1424 , \oc8051_golden_model_1.n1425 [0]);
  buf(\oc8051_golden_model_1.n1425 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1425 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1425 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1425 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1427 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n1427 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n1427 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n1427 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n1427 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n1427 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n1427 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n1427 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n1427 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1429 [8], \oc8051_golden_model_1.n1461 [7]);
  buf(\oc8051_golden_model_1.n1430 , \oc8051_golden_model_1.n1461 [7]);
  buf(\oc8051_golden_model_1.n1431 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n1431 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n1431 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n1431 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n1432 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n1432 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n1432 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n1432 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n1432 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1434 [4], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1435 , \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1436 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n1436 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n1436 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n1436 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n1436 [4], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n1436 [5], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n1436 [6], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n1436 [7], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n1436 [8], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n1443 , \oc8051_golden_model_1.n1461 [2]);
  buf(\oc8051_golden_model_1.n1444 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1444 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1444 [2], \oc8051_golden_model_1.n1461 [2]);
  buf(\oc8051_golden_model_1.n1444 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1444 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1444 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1444 [6], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1444 [7], \oc8051_golden_model_1.n1461 [7]);
  buf(\oc8051_golden_model_1.n1445 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1445 [1], \oc8051_golden_model_1.n1461 [2]);
  buf(\oc8051_golden_model_1.n1445 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1445 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1445 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1445 [5], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1445 [6], \oc8051_golden_model_1.n1461 [7]);
  buf(\oc8051_golden_model_1.n1460 , \oc8051_golden_model_1.n1474 [0]);
  buf(\oc8051_golden_model_1.n1461 [0], \oc8051_golden_model_1.n1474 [0]);
  buf(\oc8051_golden_model_1.n1461 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1461 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1461 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1461 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1461 [6], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1463 [8], \oc8051_golden_model_1.n1474 [7]);
  buf(\oc8051_golden_model_1.n1464 , \oc8051_golden_model_1.n1474 [7]);
  buf(\oc8051_golden_model_1.n1471 , \oc8051_golden_model_1.n1474 [2]);
  buf(\oc8051_golden_model_1.n1472 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1472 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1472 [2], \oc8051_golden_model_1.n1474 [2]);
  buf(\oc8051_golden_model_1.n1472 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1472 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1472 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1472 [6], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1472 [7], \oc8051_golden_model_1.n1474 [7]);
  buf(\oc8051_golden_model_1.n1473 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1473 [1], \oc8051_golden_model_1.n1474 [2]);
  buf(\oc8051_golden_model_1.n1473 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1473 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1473 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1473 [5], \oc8051_golden_model_1.n1474 [6]);
  buf(\oc8051_golden_model_1.n1473 [6], \oc8051_golden_model_1.n1474 [7]);
  buf(\oc8051_golden_model_1.n1474 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1474 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1474 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1474 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1476 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n1476 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n1476 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n1476 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n1476 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.n1476 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.n1476 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.n1476 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n1476 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1478 [8], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1479 , \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1480 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n1480 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n1480 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n1480 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n1480 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1482 [4], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1483 , \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1484 [0], \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n1484 [1], \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n1484 [2], \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n1484 [3], \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n1484 [4], \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.n1484 [5], \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.n1484 [6], \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.n1484 [7], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n1484 [8], \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n1491 , \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1492 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1492 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1492 [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1492 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1492 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1492 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1492 [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1492 [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1493 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1493 [1], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1493 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1493 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1493 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1493 [5], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1493 [6], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1508 , \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.n1509 [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.n1509 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1509 [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1509 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1509 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1509 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1509 [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1509 [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1511 [4], \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.n1512 , \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.n1513 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1513 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1513 [2], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1513 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1513 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1513 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1513 [6], \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.n1513 [7], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1514 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1514 [1], \oc8051_golden_model_1.n1515 [2]);
  buf(\oc8051_golden_model_1.n1514 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1514 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1514 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1514 [5], \oc8051_golden_model_1.n1515 [6]);
  buf(\oc8051_golden_model_1.n1514 [6], \oc8051_golden_model_1.n1515 [7]);
  buf(\oc8051_golden_model_1.n1515 [0], \oc8051_golden_model_1.n1528 [0]);
  buf(\oc8051_golden_model_1.n1515 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1515 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1515 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1515 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1517 [8], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1518 , \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1525 , \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1526 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1526 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1526 [2], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1526 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1526 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1526 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1526 [6], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1526 [7], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1527 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1527 [1], \oc8051_golden_model_1.n1528 [2]);
  buf(\oc8051_golden_model_1.n1527 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1527 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1527 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1527 [5], \oc8051_golden_model_1.n1528 [6]);
  buf(\oc8051_golden_model_1.n1527 [6], \oc8051_golden_model_1.n1528 [7]);
  buf(\oc8051_golden_model_1.n1528 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1528 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1528 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1528 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1531 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1531 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1531 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1531 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1531 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1531 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1531 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1531 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1531 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1532 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1532 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1532 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1532 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1532 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1532 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1532 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1532 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1532 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1533 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1533 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1533 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1533 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1533 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1533 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1533 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1533 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1534 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1534 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1534 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1534 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1534 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1534 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1534 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1534 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1535 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1535 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1535 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1535 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1535 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1535 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1535 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1536 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1537 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1538 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1539 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1540 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1541 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1542 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1543 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1550 , \oc8051_golden_model_1.n1551 [0]);
  buf(\oc8051_golden_model_1.n1551 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1551 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1551 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1551 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1551 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1551 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1551 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1552 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1552 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1552 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1555 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1555 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1557 [8], \oc8051_golden_model_1.n1587 [7]);
  buf(\oc8051_golden_model_1.n1558 , \oc8051_golden_model_1.n1587 [7]);
  buf(\oc8051_golden_model_1.n1559 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1559 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1559 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1559 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1559 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1561 [4], \oc8051_golden_model_1.n1587 [6]);
  buf(\oc8051_golden_model_1.n1562 , \oc8051_golden_model_1.n1587 [6]);
  buf(\oc8051_golden_model_1.n1569 , \oc8051_golden_model_1.n1587 [2]);
  buf(\oc8051_golden_model_1.n1570 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1570 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1570 [2], \oc8051_golden_model_1.n1587 [2]);
  buf(\oc8051_golden_model_1.n1570 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1570 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1570 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1570 [6], \oc8051_golden_model_1.n1587 [6]);
  buf(\oc8051_golden_model_1.n1570 [7], \oc8051_golden_model_1.n1587 [7]);
  buf(\oc8051_golden_model_1.n1571 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1571 [1], \oc8051_golden_model_1.n1587 [2]);
  buf(\oc8051_golden_model_1.n1571 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1571 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1571 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1571 [5], \oc8051_golden_model_1.n1587 [6]);
  buf(\oc8051_golden_model_1.n1571 [6], \oc8051_golden_model_1.n1587 [7]);
  buf(\oc8051_golden_model_1.n1586 , \oc8051_golden_model_1.n1587 [0]);
  buf(\oc8051_golden_model_1.n1587 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1587 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1587 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1587 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1591 [8], \oc8051_golden_model_1.n1620 [7]);
  buf(\oc8051_golden_model_1.n1592 , \oc8051_golden_model_1.n1620 [7]);
  buf(\oc8051_golden_model_1.n1594 [4], \oc8051_golden_model_1.n1620 [6]);
  buf(\oc8051_golden_model_1.n1595 , \oc8051_golden_model_1.n1620 [6]);
  buf(\oc8051_golden_model_1.n1602 , \oc8051_golden_model_1.n1620 [2]);
  buf(\oc8051_golden_model_1.n1603 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1603 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1603 [2], \oc8051_golden_model_1.n1620 [2]);
  buf(\oc8051_golden_model_1.n1603 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1603 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1603 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1603 [6], \oc8051_golden_model_1.n1620 [6]);
  buf(\oc8051_golden_model_1.n1603 [7], \oc8051_golden_model_1.n1620 [7]);
  buf(\oc8051_golden_model_1.n1604 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1604 [1], \oc8051_golden_model_1.n1620 [2]);
  buf(\oc8051_golden_model_1.n1604 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1604 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1604 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1604 [5], \oc8051_golden_model_1.n1620 [6]);
  buf(\oc8051_golden_model_1.n1604 [6], \oc8051_golden_model_1.n1620 [7]);
  buf(\oc8051_golden_model_1.n1619 , \oc8051_golden_model_1.n1620 [0]);
  buf(\oc8051_golden_model_1.n1620 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1620 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1620 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1620 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1624 [8], \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.n1625 , \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.n1627 [4], \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.n1628 , \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.n1635 , \oc8051_golden_model_1.n1653 [2]);
  buf(\oc8051_golden_model_1.n1636 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1636 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1636 [2], \oc8051_golden_model_1.n1653 [2]);
  buf(\oc8051_golden_model_1.n1636 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1636 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1636 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1636 [6], \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.n1636 [7], \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.n1637 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1637 [1], \oc8051_golden_model_1.n1653 [2]);
  buf(\oc8051_golden_model_1.n1637 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1637 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1637 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1637 [5], \oc8051_golden_model_1.n1653 [6]);
  buf(\oc8051_golden_model_1.n1637 [6], \oc8051_golden_model_1.n1653 [7]);
  buf(\oc8051_golden_model_1.n1652 , \oc8051_golden_model_1.n1653 [0]);
  buf(\oc8051_golden_model_1.n1653 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1653 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1653 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1653 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1657 [8], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.n1658 , \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.n1660 [4], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.n1661 , \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.n1668 , \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.n1669 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1669 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1669 [2], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.n1669 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1669 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1669 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1669 [6], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.n1669 [7], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.n1670 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1670 [1], \oc8051_golden_model_1.n1686 [2]);
  buf(\oc8051_golden_model_1.n1670 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1670 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1670 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1670 [5], \oc8051_golden_model_1.n1686 [6]);
  buf(\oc8051_golden_model_1.n1670 [6], \oc8051_golden_model_1.n1686 [7]);
  buf(\oc8051_golden_model_1.n1685 , \oc8051_golden_model_1.n1686 [0]);
  buf(\oc8051_golden_model_1.n1686 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1686 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1686 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1686 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1700 [1], \oc8051_golden_model_1.n1702 [1]);
  buf(\oc8051_golden_model_1.n1700 [2], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1700 [3], \oc8051_golden_model_1.n1702 [3]);
  buf(\oc8051_golden_model_1.n1700 [4], \oc8051_golden_model_1.n1702 [4]);
  buf(\oc8051_golden_model_1.n1700 [5], \oc8051_golden_model_1.n1702 [5]);
  buf(\oc8051_golden_model_1.n1700 [6], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1700 [7], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1701 [0], \oc8051_golden_model_1.n1702 [1]);
  buf(\oc8051_golden_model_1.n1701 [1], \oc8051_golden_model_1.n1702 [2]);
  buf(\oc8051_golden_model_1.n1701 [2], \oc8051_golden_model_1.n1702 [3]);
  buf(\oc8051_golden_model_1.n1701 [3], \oc8051_golden_model_1.n1702 [4]);
  buf(\oc8051_golden_model_1.n1701 [4], \oc8051_golden_model_1.n1702 [5]);
  buf(\oc8051_golden_model_1.n1701 [5], \oc8051_golden_model_1.n1702 [6]);
  buf(\oc8051_golden_model_1.n1701 [6], \oc8051_golden_model_1.n1702 [7]);
  buf(\oc8051_golden_model_1.n1702 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n1746 , \oc8051_golden_model_1.n1747 [0]);
  buf(\oc8051_golden_model_1.n1747 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1747 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1747 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1747 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1747 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1747 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1747 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1763 , \oc8051_golden_model_1.n1764 [0]);
  buf(\oc8051_golden_model_1.n1764 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1764 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1764 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1764 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1764 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1764 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1764 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1780 , \oc8051_golden_model_1.n1781 [0]);
  buf(\oc8051_golden_model_1.n1781 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1781 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1781 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1781 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1781 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1781 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1781 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1797 , \oc8051_golden_model_1.n1798 [0]);
  buf(\oc8051_golden_model_1.n1798 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1798 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1798 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1798 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1798 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1798 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1798 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1810 [1], \oc8051_golden_model_1.n1812 [1]);
  buf(\oc8051_golden_model_1.n1810 [2], \oc8051_golden_model_1.n1812 [2]);
  buf(\oc8051_golden_model_1.n1810 [3], \oc8051_golden_model_1.n1812 [3]);
  buf(\oc8051_golden_model_1.n1810 [4], \oc8051_golden_model_1.n1812 [4]);
  buf(\oc8051_golden_model_1.n1810 [5], \oc8051_golden_model_1.n1812 [5]);
  buf(\oc8051_golden_model_1.n1810 [6], \oc8051_golden_model_1.n1812 [6]);
  buf(\oc8051_golden_model_1.n1810 [7], \oc8051_golden_model_1.n1812 [7]);
  buf(\oc8051_golden_model_1.n1811 [0], \oc8051_golden_model_1.n1812 [1]);
  buf(\oc8051_golden_model_1.n1811 [1], \oc8051_golden_model_1.n1812 [2]);
  buf(\oc8051_golden_model_1.n1811 [2], \oc8051_golden_model_1.n1812 [3]);
  buf(\oc8051_golden_model_1.n1811 [3], \oc8051_golden_model_1.n1812 [4]);
  buf(\oc8051_golden_model_1.n1811 [4], \oc8051_golden_model_1.n1812 [5]);
  buf(\oc8051_golden_model_1.n1811 [5], \oc8051_golden_model_1.n1812 [6]);
  buf(\oc8051_golden_model_1.n1811 [6], \oc8051_golden_model_1.n1812 [7]);
  buf(\oc8051_golden_model_1.n1812 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n1856 , \oc8051_golden_model_1.n1857 [0]);
  buf(\oc8051_golden_model_1.n1857 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1857 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1857 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1857 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1857 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1857 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1857 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1873 , \oc8051_golden_model_1.n1874 [0]);
  buf(\oc8051_golden_model_1.n1874 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1874 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1874 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1874 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1874 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1874 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1874 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1890 , \oc8051_golden_model_1.n1891 [0]);
  buf(\oc8051_golden_model_1.n1891 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1891 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1891 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1891 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1891 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1891 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1891 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1907 , \oc8051_golden_model_1.n1908 [0]);
  buf(\oc8051_golden_model_1.n1908 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1908 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1908 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1908 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1908 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1908 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1908 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1983 , \oc8051_golden_model_1.n1984 [0]);
  buf(\oc8051_golden_model_1.n1984 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1984 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1984 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1984 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1984 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1984 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1984 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2000 , \oc8051_golden_model_1.n2001 [0]);
  buf(\oc8051_golden_model_1.n2001 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2001 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2001 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2001 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2001 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2001 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2001 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2017 , \oc8051_golden_model_1.n2018 [0]);
  buf(\oc8051_golden_model_1.n2018 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2018 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2018 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2018 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2018 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2018 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2018 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2034 , \oc8051_golden_model_1.n2035 [0]);
  buf(\oc8051_golden_model_1.n2035 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2035 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2035 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2035 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2035 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2039 , \oc8051_golden_model_1.n2043 [7]);
  buf(\oc8051_golden_model_1.n2040 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2040 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2040 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2040 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2040 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2040 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2040 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2041 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2041 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2041 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2041 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2041 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2041 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2041 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2041 [7], \oc8051_golden_model_1.n2043 [7]);
  buf(\oc8051_golden_model_1.n2042 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2042 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2042 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2042 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2042 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2042 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2042 [6], \oc8051_golden_model_1.n2043 [7]);
  buf(\oc8051_golden_model_1.n2043 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2043 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2043 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2043 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2043 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2043 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2043 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2058 , \oc8051_golden_model_1.n2059 [0]);
  buf(\oc8051_golden_model_1.n2059 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2059 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2059 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2059 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2059 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2059 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2059 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2087 , \oc8051_golden_model_1.n2090 [7]);
  buf(\oc8051_golden_model_1.n2088 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2088 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2088 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2088 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2088 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2088 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2088 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2088 [7], \oc8051_golden_model_1.n2090 [7]);
  buf(\oc8051_golden_model_1.n2089 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2089 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2089 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2089 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2089 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2089 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2089 [6], \oc8051_golden_model_1.n2090 [7]);
  buf(\oc8051_golden_model_1.n2090 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2090 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2090 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2090 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2090 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2090 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2090 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2097 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2097 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2097 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2097 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2098 , \oc8051_golden_model_1.n2116 [2]);
  buf(\oc8051_golden_model_1.n2099 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2099 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2099 [2], \oc8051_golden_model_1.n2116 [2]);
  buf(\oc8051_golden_model_1.n2099 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2099 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2099 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2099 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2099 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2100 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2100 [1], \oc8051_golden_model_1.n2116 [2]);
  buf(\oc8051_golden_model_1.n2100 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2100 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2100 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2100 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2100 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2115 , \oc8051_golden_model_1.n2116 [0]);
  buf(\oc8051_golden_model_1.n2116 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2116 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2116 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2116 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2116 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2116 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2273 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2273 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2276 , \oc8051_golden_model_1.n2302 [7]);
  buf(\oc8051_golden_model_1.n2278 , \oc8051_golden_model_1.n2302 [6]);
  buf(\oc8051_golden_model_1.n2284 , \oc8051_golden_model_1.n2302 [2]);
  buf(\oc8051_golden_model_1.n2285 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2285 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2285 [2], \oc8051_golden_model_1.n2302 [2]);
  buf(\oc8051_golden_model_1.n2285 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2285 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2285 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2285 [6], \oc8051_golden_model_1.n2302 [6]);
  buf(\oc8051_golden_model_1.n2285 [7], \oc8051_golden_model_1.n2302 [7]);
  buf(\oc8051_golden_model_1.n2286 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2286 [1], \oc8051_golden_model_1.n2302 [2]);
  buf(\oc8051_golden_model_1.n2286 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2286 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2286 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2286 [5], \oc8051_golden_model_1.n2302 [6]);
  buf(\oc8051_golden_model_1.n2286 [6], \oc8051_golden_model_1.n2302 [7]);
  buf(\oc8051_golden_model_1.n2301 , \oc8051_golden_model_1.n2302 [0]);
  buf(\oc8051_golden_model_1.n2302 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2302 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2302 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2302 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2306 , \oc8051_golden_model_1.n2332 [7]);
  buf(\oc8051_golden_model_1.n2308 , \oc8051_golden_model_1.n2332 [6]);
  buf(\oc8051_golden_model_1.n2314 , \oc8051_golden_model_1.n2332 [2]);
  buf(\oc8051_golden_model_1.n2315 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2315 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2315 [2], \oc8051_golden_model_1.n2332 [2]);
  buf(\oc8051_golden_model_1.n2315 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2315 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2315 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2315 [6], \oc8051_golden_model_1.n2332 [6]);
  buf(\oc8051_golden_model_1.n2315 [7], \oc8051_golden_model_1.n2332 [7]);
  buf(\oc8051_golden_model_1.n2316 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2316 [1], \oc8051_golden_model_1.n2332 [2]);
  buf(\oc8051_golden_model_1.n2316 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2316 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2316 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2316 [5], \oc8051_golden_model_1.n2332 [6]);
  buf(\oc8051_golden_model_1.n2316 [6], \oc8051_golden_model_1.n2332 [7]);
  buf(\oc8051_golden_model_1.n2331 , \oc8051_golden_model_1.n2332 [0]);
  buf(\oc8051_golden_model_1.n2332 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2332 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2332 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2332 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2336 , \oc8051_golden_model_1.n2362 [7]);
  buf(\oc8051_golden_model_1.n2338 , \oc8051_golden_model_1.n2362 [6]);
  buf(\oc8051_golden_model_1.n2344 , \oc8051_golden_model_1.n2362 [2]);
  buf(\oc8051_golden_model_1.n2345 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2345 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2345 [2], \oc8051_golden_model_1.n2362 [2]);
  buf(\oc8051_golden_model_1.n2345 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2345 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2345 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2345 [6], \oc8051_golden_model_1.n2362 [6]);
  buf(\oc8051_golden_model_1.n2345 [7], \oc8051_golden_model_1.n2362 [7]);
  buf(\oc8051_golden_model_1.n2346 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2346 [1], \oc8051_golden_model_1.n2362 [2]);
  buf(\oc8051_golden_model_1.n2346 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2346 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2346 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2346 [5], \oc8051_golden_model_1.n2362 [6]);
  buf(\oc8051_golden_model_1.n2346 [6], \oc8051_golden_model_1.n2362 [7]);
  buf(\oc8051_golden_model_1.n2361 , \oc8051_golden_model_1.n2362 [0]);
  buf(\oc8051_golden_model_1.n2362 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2362 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2362 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2362 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2366 , \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.n2368 , \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.n2374 , \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.n2375 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2375 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2375 [2], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.n2375 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2375 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2375 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2375 [6], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.n2375 [7], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.n2376 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2376 [1], \oc8051_golden_model_1.n2392 [2]);
  buf(\oc8051_golden_model_1.n2376 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2376 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2376 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2376 [5], \oc8051_golden_model_1.n2392 [6]);
  buf(\oc8051_golden_model_1.n2376 [6], \oc8051_golden_model_1.n2392 [7]);
  buf(\oc8051_golden_model_1.n2391 , \oc8051_golden_model_1.n2392 [0]);
  buf(\oc8051_golden_model_1.n2392 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2392 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2392 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2392 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2394 , \oc8051_golden_model_1.n2397 [7]);
  buf(\oc8051_golden_model_1.n2395 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2395 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2395 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2395 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2395 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2395 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2395 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2395 [7], \oc8051_golden_model_1.n2397 [7]);
  buf(\oc8051_golden_model_1.n2396 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2396 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2396 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2396 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2396 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2396 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2396 [6], \oc8051_golden_model_1.n2397 [7]);
  buf(\oc8051_golden_model_1.n2397 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2397 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2397 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2397 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2397 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2397 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2397 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2398 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2398 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2398 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2398 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2398 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2398 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2398 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2398 [7], \oc8051_golden_model_1.n2400 [7]);
  buf(\oc8051_golden_model_1.n2399 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2399 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2399 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2399 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2399 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2399 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2399 [6], \oc8051_golden_model_1.n2400 [7]);
  buf(\oc8051_golden_model_1.n2400 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2400 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2400 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2400 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2400 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2400 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2400 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2404 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n2404 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n2404 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n2404 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n2404 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n2404 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n2404 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n2404 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n2404 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2404 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2410 , \oc8051_golden_model_1.n2428 [2]);
  buf(\oc8051_golden_model_1.n2411 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2411 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2411 [2], \oc8051_golden_model_1.n2428 [2]);
  buf(\oc8051_golden_model_1.n2411 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2411 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2411 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2411 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2411 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2412 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2412 [1], \oc8051_golden_model_1.n2428 [2]);
  buf(\oc8051_golden_model_1.n2412 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2412 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2412 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2412 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2412 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2427 , \oc8051_golden_model_1.n2428 [0]);
  buf(\oc8051_golden_model_1.n2428 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2428 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2428 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2428 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2428 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2428 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2430 , \oc8051_golden_model_1.n2433 [7]);
  buf(\oc8051_golden_model_1.n2431 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2431 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2431 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2431 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2431 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2431 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2431 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2431 [7], \oc8051_golden_model_1.n2433 [7]);
  buf(\oc8051_golden_model_1.n2432 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2432 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2432 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2432 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2432 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2432 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2432 [6], \oc8051_golden_model_1.n2433 [7]);
  buf(\oc8051_golden_model_1.n2433 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2433 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2433 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2433 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2433 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2433 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2433 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2461 , \oc8051_golden_model_1.n2464 [7]);
  buf(\oc8051_golden_model_1.n2462 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2462 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2462 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2462 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2462 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2462 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2462 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2462 [7], \oc8051_golden_model_1.n2464 [7]);
  buf(\oc8051_golden_model_1.n2463 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2463 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2463 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2463 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2463 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2463 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2463 [6], \oc8051_golden_model_1.n2464 [7]);
  buf(\oc8051_golden_model_1.n2464 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2464 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2464 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2464 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2464 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2464 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2464 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2469 , \oc8051_golden_model_1.n2472 [7]);
  buf(\oc8051_golden_model_1.n2470 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2470 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2470 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2470 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2470 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2470 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2470 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2470 [7], \oc8051_golden_model_1.n2472 [7]);
  buf(\oc8051_golden_model_1.n2471 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2471 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2471 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2471 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2471 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2471 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2471 [6], \oc8051_golden_model_1.n2472 [7]);
  buf(\oc8051_golden_model_1.n2472 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2472 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2472 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2472 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2472 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2472 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2472 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2477 , \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2478 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2478 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2478 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2478 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2478 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2478 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2478 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2478 [7], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2479 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2479 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2479 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2479 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2479 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2479 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2479 [6], \oc8051_golden_model_1.n2480 [7]);
  buf(\oc8051_golden_model_1.n2480 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2480 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2480 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2480 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2480 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2480 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2480 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2485 , \oc8051_golden_model_1.n2488 [7]);
  buf(\oc8051_golden_model_1.n2486 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2486 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2486 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2486 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2486 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2486 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2486 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2486 [7], \oc8051_golden_model_1.n2488 [7]);
  buf(\oc8051_golden_model_1.n2487 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2487 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2487 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2487 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2487 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2487 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2487 [6], \oc8051_golden_model_1.n2488 [7]);
  buf(\oc8051_golden_model_1.n2488 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2488 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2488 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2488 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2488 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2488 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2488 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2493 , \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.n2494 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2494 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2494 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2494 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2494 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2494 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2494 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2494 [7], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.n2495 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2495 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2495 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2495 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2495 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2495 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2495 [6], \oc8051_golden_model_1.n2496 [7]);
  buf(\oc8051_golden_model_1.n2496 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2496 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2496 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2496 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2496 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2496 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2496 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2517 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2517 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2517 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2517 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2517 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2517 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2517 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2517 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2518 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2518 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2518 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2518 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2518 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2518 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2518 [6], 1'b0);
  buf(\oc8051_golden_model_1.n2519 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2519 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2519 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2519 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2519 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2519 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2519 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2519 [7], 1'b0);
  buf(\oc8051_golden_model_1.n2520 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2520 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2520 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2520 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2521 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2521 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2521 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2521 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2521 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2521 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2521 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2521 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2522 , \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2523 , \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2524 , \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2525 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2526 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2527 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2528 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2529 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2536 , \oc8051_golden_model_1.n2537 [0]);
  buf(\oc8051_golden_model_1.n2537 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2537 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2537 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2537 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2537 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2537 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2537 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2546 [1], \oc8051_golden_model_1.n2741 [1]);
  buf(\oc8051_golden_model_1.n2546 [2], \oc8051_golden_model_1.n2741 [2]);
  buf(\oc8051_golden_model_1.n2546 [3], \oc8051_golden_model_1.n2741 [3]);
  buf(\oc8051_golden_model_1.n2546 [4], \oc8051_golden_model_1.n2741 [4]);
  buf(\oc8051_golden_model_1.n2546 [5], \oc8051_golden_model_1.n2741 [5]);
  buf(\oc8051_golden_model_1.n2546 [6], \oc8051_golden_model_1.n2741 [6]);
  buf(\oc8051_golden_model_1.n2546 [7], \oc8051_golden_model_1.n2741 [7]);
  buf(\oc8051_golden_model_1.n2547 [0], \oc8051_golden_model_1.n2741 [1]);
  buf(\oc8051_golden_model_1.n2547 [1], \oc8051_golden_model_1.n2741 [2]);
  buf(\oc8051_golden_model_1.n2547 [2], \oc8051_golden_model_1.n2741 [3]);
  buf(\oc8051_golden_model_1.n2547 [3], \oc8051_golden_model_1.n2741 [4]);
  buf(\oc8051_golden_model_1.n2547 [4], \oc8051_golden_model_1.n2741 [5]);
  buf(\oc8051_golden_model_1.n2547 [5], \oc8051_golden_model_1.n2741 [6]);
  buf(\oc8051_golden_model_1.n2547 [6], \oc8051_golden_model_1.n2741 [7]);
  buf(\oc8051_golden_model_1.n2562 , \oc8051_golden_model_1.n2723 [0]);
  buf(\oc8051_golden_model_1.n2563 [0], \oc8051_golden_model_1.n2723 [0]);
  buf(\oc8051_golden_model_1.n2563 [1], \oc8051_golden_model_1.n2741 [1]);
  buf(\oc8051_golden_model_1.n2563 [2], \oc8051_golden_model_1.n2741 [2]);
  buf(\oc8051_golden_model_1.n2563 [3], \oc8051_golden_model_1.n2741 [3]);
  buf(\oc8051_golden_model_1.n2563 [4], \oc8051_golden_model_1.n2741 [4]);
  buf(\oc8051_golden_model_1.n2563 [5], \oc8051_golden_model_1.n2741 [5]);
  buf(\oc8051_golden_model_1.n2563 [6], \oc8051_golden_model_1.n2741 [6]);
  buf(\oc8051_golden_model_1.n2563 [7], \oc8051_golden_model_1.n2741 [7]);
  buf(\oc8051_golden_model_1.n2564 , \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n2565 , \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n2566 , \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n2567 , \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n2568 , \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n2569 , \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n2570 , \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n2571 , \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n2578 , \oc8051_golden_model_1.n2579 [0]);
  buf(\oc8051_golden_model_1.n2579 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2579 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2579 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2579 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2579 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2579 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2579 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2580 , \oc8051_golden_model_1.n2706 [7]);
  buf(\oc8051_golden_model_1.n2581 , \oc8051_golden_model_1.n2706 [6]);
  buf(\oc8051_golden_model_1.n2582 , \oc8051_golden_model_1.n2706 [5]);
  buf(\oc8051_golden_model_1.n2583 , \oc8051_golden_model_1.n2706 [4]);
  buf(\oc8051_golden_model_1.n2584 , \oc8051_golden_model_1.n2706 [3]);
  buf(\oc8051_golden_model_1.n2585 , \oc8051_golden_model_1.n2706 [2]);
  buf(\oc8051_golden_model_1.n2586 , \oc8051_golden_model_1.n2706 [1]);
  buf(\oc8051_golden_model_1.n2587 , \oc8051_golden_model_1.n2706 [0]);
  buf(\oc8051_golden_model_1.n2594 , \oc8051_golden_model_1.n2595 [0]);
  buf(\oc8051_golden_model_1.n2595 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2595 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2595 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2595 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2595 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2595 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2595 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2625 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2625 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2625 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2625 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2625 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2625 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2625 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2625 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2626 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2626 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2626 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2626 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2626 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2626 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2626 [6], 1'b1);
  buf(\oc8051_golden_model_1.n2627 [0], \oc8051_golden_model_1.n2741 [0]);
  buf(\oc8051_golden_model_1.n2627 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2627 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2627 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2627 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2627 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2627 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2627 [7], 1'b1);
  buf(\oc8051_golden_model_1.n2646 , \oc8051_golden_model_1.n2664 [7]);
  buf(\oc8051_golden_model_1.n2647 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n2647 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2647 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2647 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2647 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2647 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2647 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2647 [7], \oc8051_golden_model_1.n2664 [7]);
  buf(\oc8051_golden_model_1.n2648 [0], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2648 [1], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2648 [2], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2648 [3], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2648 [4], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2648 [5], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2648 [6], \oc8051_golden_model_1.n2664 [7]);
  buf(\oc8051_golden_model_1.n2663 , \oc8051_golden_model_1.n2664 [0]);
  buf(\oc8051_golden_model_1.n2664 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2664 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2664 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2664 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2664 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2664 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2668 [0], \oc8051_golden_model_1.n2678 );
  buf(\oc8051_golden_model_1.n2668 [1], \oc8051_golden_model_1.n2677 );
  buf(\oc8051_golden_model_1.n2668 [2], \oc8051_golden_model_1.n2676 );
  buf(\oc8051_golden_model_1.n2668 [3], \oc8051_golden_model_1.n2675 );
  buf(\oc8051_golden_model_1.n2668 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2668 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2668 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2668 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2669 [0], \oc8051_golden_model_1.n2670 [4]);
  buf(\oc8051_golden_model_1.n2669 [1], \oc8051_golden_model_1.n2670 [5]);
  buf(\oc8051_golden_model_1.n2669 [2], \oc8051_golden_model_1.n2670 [6]);
  buf(\oc8051_golden_model_1.n2669 [3], \oc8051_golden_model_1.n2670 [7]);
  buf(\oc8051_golden_model_1.n2670 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n2670 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n2670 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n2670 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n2671 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n2672 , \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n2673 , \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n2674 , \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n2685 , \oc8051_golden_model_1.n2686 [0]);
  buf(\oc8051_golden_model_1.n2686 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2686 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2686 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2686 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2686 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2686 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2686 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2690 , \oc8051_golden_model_1.XRAM_DATA_IN [7]);
  buf(\oc8051_golden_model_1.n2691 , \oc8051_golden_model_1.XRAM_DATA_IN [6]);
  buf(\oc8051_golden_model_1.n2692 , \oc8051_golden_model_1.XRAM_DATA_IN [5]);
  buf(\oc8051_golden_model_1.n2693 , \oc8051_golden_model_1.XRAM_DATA_IN [4]);
  buf(\oc8051_golden_model_1.n2694 , \oc8051_golden_model_1.XRAM_DATA_IN [3]);
  buf(\oc8051_golden_model_1.n2695 , \oc8051_golden_model_1.XRAM_DATA_IN [2]);
  buf(\oc8051_golden_model_1.n2696 , \oc8051_golden_model_1.XRAM_DATA_IN [1]);
  buf(\oc8051_golden_model_1.n2697 , \oc8051_golden_model_1.XRAM_DATA_IN [0]);
  buf(\oc8051_golden_model_1.n2704 , \oc8051_golden_model_1.n2705 [0]);
  buf(\oc8051_golden_model_1.n2705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2705 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2705 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2705 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2706 [8], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [9], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [10], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [11], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [12], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [13], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [14], 1'b0);
  buf(\oc8051_golden_model_1.n2706 [15], 1'b0);
  buf(\oc8051_golden_model_1.n2721 , \oc8051_golden_model_1.n2722 [0]);
  buf(\oc8051_golden_model_1.n2722 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2722 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2722 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2722 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2722 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2722 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2722 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2723 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2723 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2723 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2723 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2723 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2723 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2723 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n2739 , \oc8051_golden_model_1.n2740 [0]);
  buf(\oc8051_golden_model_1.n2740 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n2740 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n2740 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n2740 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n2740 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n2740 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n2740 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw_impl[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(TMOD_gm_next[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm_next[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm_next[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm_next[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm_next[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm_next[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm_next[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm_next[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TMOD_gm[0], \oc8051_golden_model_1.TMOD [0]);
  buf(TMOD_gm[1], \oc8051_golden_model_1.TMOD [1]);
  buf(TMOD_gm[2], \oc8051_golden_model_1.TMOD [2]);
  buf(TMOD_gm[3], \oc8051_golden_model_1.TMOD [3]);
  buf(TMOD_gm[4], \oc8051_golden_model_1.TMOD [4]);
  buf(TMOD_gm[5], \oc8051_golden_model_1.TMOD [5]);
  buf(TMOD_gm[6], \oc8051_golden_model_1.TMOD [6]);
  buf(TMOD_gm[7], \oc8051_golden_model_1.TMOD [7]);
  buf(TL1_gm_next[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm_next[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm_next[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm_next[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm_next[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm_next[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm_next[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm_next[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL1_gm[0], \oc8051_golden_model_1.TL1 [0]);
  buf(TL1_gm[1], \oc8051_golden_model_1.TL1 [1]);
  buf(TL1_gm[2], \oc8051_golden_model_1.TL1 [2]);
  buf(TL1_gm[3], \oc8051_golden_model_1.TL1 [3]);
  buf(TL1_gm[4], \oc8051_golden_model_1.TL1 [4]);
  buf(TL1_gm[5], \oc8051_golden_model_1.TL1 [5]);
  buf(TL1_gm[6], \oc8051_golden_model_1.TL1 [6]);
  buf(TL1_gm[7], \oc8051_golden_model_1.TL1 [7]);
  buf(TL0_gm_next[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm_next[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm_next[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm_next[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm_next[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm_next[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm_next[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm_next[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TL0_gm[0], \oc8051_golden_model_1.TL0 [0]);
  buf(TL0_gm[1], \oc8051_golden_model_1.TL0 [1]);
  buf(TL0_gm[2], \oc8051_golden_model_1.TL0 [2]);
  buf(TL0_gm[3], \oc8051_golden_model_1.TL0 [3]);
  buf(TL0_gm[4], \oc8051_golden_model_1.TL0 [4]);
  buf(TL0_gm[5], \oc8051_golden_model_1.TL0 [5]);
  buf(TL0_gm[6], \oc8051_golden_model_1.TL0 [6]);
  buf(TL0_gm[7], \oc8051_golden_model_1.TL0 [7]);
  buf(TH1_gm_next[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm_next[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm_next[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm_next[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm_next[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm_next[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm_next[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm_next[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH1_gm[0], \oc8051_golden_model_1.TH1 [0]);
  buf(TH1_gm[1], \oc8051_golden_model_1.TH1 [1]);
  buf(TH1_gm[2], \oc8051_golden_model_1.TH1 [2]);
  buf(TH1_gm[3], \oc8051_golden_model_1.TH1 [3]);
  buf(TH1_gm[4], \oc8051_golden_model_1.TH1 [4]);
  buf(TH1_gm[5], \oc8051_golden_model_1.TH1 [5]);
  buf(TH1_gm[6], \oc8051_golden_model_1.TH1 [6]);
  buf(TH1_gm[7], \oc8051_golden_model_1.TH1 [7]);
  buf(TH0_gm_next[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm_next[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm_next[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm_next[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm_next[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm_next[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm_next[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm_next[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TH0_gm[0], \oc8051_golden_model_1.TH0 [0]);
  buf(TH0_gm[1], \oc8051_golden_model_1.TH0 [1]);
  buf(TH0_gm[2], \oc8051_golden_model_1.TH0 [2]);
  buf(TH0_gm[3], \oc8051_golden_model_1.TH0 [3]);
  buf(TH0_gm[4], \oc8051_golden_model_1.TH0 [4]);
  buf(TH0_gm[5], \oc8051_golden_model_1.TH0 [5]);
  buf(TH0_gm[6], \oc8051_golden_model_1.TH0 [6]);
  buf(TH0_gm[7], \oc8051_golden_model_1.TH0 [7]);
  buf(TCON_gm_next[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm_next[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm_next[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm_next[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm_next[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm_next[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm_next[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm_next[7], \oc8051_golden_model_1.TCON [7]);
  buf(TCON_gm[0], \oc8051_golden_model_1.TCON [0]);
  buf(TCON_gm[1], \oc8051_golden_model_1.TCON [1]);
  buf(TCON_gm[2], \oc8051_golden_model_1.TCON [2]);
  buf(TCON_gm[3], \oc8051_golden_model_1.TCON [3]);
  buf(TCON_gm[4], \oc8051_golden_model_1.TCON [4]);
  buf(TCON_gm[5], \oc8051_golden_model_1.TCON [5]);
  buf(TCON_gm[6], \oc8051_golden_model_1.TCON [6]);
  buf(TCON_gm[7], \oc8051_golden_model_1.TCON [7]);
  buf(SP_gm[0], \oc8051_golden_model_1.SP [0]);
  buf(SP_gm[1], \oc8051_golden_model_1.SP [1]);
  buf(SP_gm[2], \oc8051_golden_model_1.SP [2]);
  buf(SP_gm[3], \oc8051_golden_model_1.SP [3]);
  buf(SP_gm[4], \oc8051_golden_model_1.SP [4]);
  buf(SP_gm[5], \oc8051_golden_model_1.SP [5]);
  buf(SP_gm[6], \oc8051_golden_model_1.SP [6]);
  buf(SP_gm[7], \oc8051_golden_model_1.SP [7]);
  buf(SCON_gm_next[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm_next[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm_next[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm_next[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm_next[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm_next[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm_next[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm_next[7], \oc8051_golden_model_1.SCON [7]);
  buf(SCON_gm[0], \oc8051_golden_model_1.SCON [0]);
  buf(SCON_gm[1], \oc8051_golden_model_1.SCON [1]);
  buf(SCON_gm[2], \oc8051_golden_model_1.SCON [2]);
  buf(SCON_gm[3], \oc8051_golden_model_1.SCON [3]);
  buf(SCON_gm[4], \oc8051_golden_model_1.SCON [4]);
  buf(SCON_gm[5], \oc8051_golden_model_1.SCON [5]);
  buf(SCON_gm[6], \oc8051_golden_model_1.SCON [6]);
  buf(SCON_gm[7], \oc8051_golden_model_1.SCON [7]);
  buf(SBUF_gm_next[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm_next[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm_next[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm_next[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm_next[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm_next[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm_next[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm_next[7], \oc8051_golden_model_1.SBUF [7]);
  buf(SBUF_gm[0], \oc8051_golden_model_1.SBUF [0]);
  buf(SBUF_gm[1], \oc8051_golden_model_1.SBUF [1]);
  buf(SBUF_gm[2], \oc8051_golden_model_1.SBUF [2]);
  buf(SBUF_gm[3], \oc8051_golden_model_1.SBUF [3]);
  buf(SBUF_gm[4], \oc8051_golden_model_1.SBUF [4]);
  buf(SBUF_gm[5], \oc8051_golden_model_1.SBUF [5]);
  buf(SBUF_gm[6], \oc8051_golden_model_1.SBUF [6]);
  buf(SBUF_gm[7], \oc8051_golden_model_1.SBUF [7]);
  buf(PSW_gm[0], \oc8051_golden_model_1.PSW [0]);
  buf(PSW_gm[1], \oc8051_golden_model_1.PSW [1]);
  buf(PSW_gm[2], \oc8051_golden_model_1.PSW [2]);
  buf(PSW_gm[3], \oc8051_golden_model_1.PSW [3]);
  buf(PSW_gm[4], \oc8051_golden_model_1.PSW [4]);
  buf(PSW_gm[5], \oc8051_golden_model_1.PSW [5]);
  buf(PSW_gm[6], \oc8051_golden_model_1.PSW [6]);
  buf(PSW_gm[7], \oc8051_golden_model_1.PSW [7]);
  buf(PCON_gm_next[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm_next[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm_next[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm_next[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm_next[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm_next[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm_next[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm_next[7], \oc8051_golden_model_1.PCON [7]);
  buf(PCON_gm[0], \oc8051_golden_model_1.PCON [0]);
  buf(PCON_gm[1], \oc8051_golden_model_1.PCON [1]);
  buf(PCON_gm[2], \oc8051_golden_model_1.PCON [2]);
  buf(PCON_gm[3], \oc8051_golden_model_1.PCON [3]);
  buf(PCON_gm[4], \oc8051_golden_model_1.PCON [4]);
  buf(PCON_gm[5], \oc8051_golden_model_1.PCON [5]);
  buf(PCON_gm[6], \oc8051_golden_model_1.PCON [6]);
  buf(PCON_gm[7], \oc8051_golden_model_1.PCON [7]);
  buf(P3_gm[0], \oc8051_golden_model_1.P3 [0]);
  buf(P3_gm[1], \oc8051_golden_model_1.P3 [1]);
  buf(P3_gm[2], \oc8051_golden_model_1.P3 [2]);
  buf(P3_gm[3], \oc8051_golden_model_1.P3 [3]);
  buf(P3_gm[4], \oc8051_golden_model_1.P3 [4]);
  buf(P3_gm[5], \oc8051_golden_model_1.P3 [5]);
  buf(P3_gm[6], \oc8051_golden_model_1.P3 [6]);
  buf(P3_gm[7], \oc8051_golden_model_1.P3 [7]);
  buf(P2_gm[0], \oc8051_golden_model_1.P2 [0]);
  buf(P2_gm[1], \oc8051_golden_model_1.P2 [1]);
  buf(P2_gm[2], \oc8051_golden_model_1.P2 [2]);
  buf(P2_gm[3], \oc8051_golden_model_1.P2 [3]);
  buf(P2_gm[4], \oc8051_golden_model_1.P2 [4]);
  buf(P2_gm[5], \oc8051_golden_model_1.P2 [5]);
  buf(P2_gm[6], \oc8051_golden_model_1.P2 [6]);
  buf(P2_gm[7], \oc8051_golden_model_1.P2 [7]);
  buf(P1_gm[0], \oc8051_golden_model_1.P1 [0]);
  buf(P1_gm[1], \oc8051_golden_model_1.P1 [1]);
  buf(P1_gm[2], \oc8051_golden_model_1.P1 [2]);
  buf(P1_gm[3], \oc8051_golden_model_1.P1 [3]);
  buf(P1_gm[4], \oc8051_golden_model_1.P1 [4]);
  buf(P1_gm[5], \oc8051_golden_model_1.P1 [5]);
  buf(P1_gm[6], \oc8051_golden_model_1.P1 [6]);
  buf(P1_gm[7], \oc8051_golden_model_1.P1 [7]);
  buf(P0_gm[0], \oc8051_golden_model_1.P0 [0]);
  buf(P0_gm[1], \oc8051_golden_model_1.P0 [1]);
  buf(P0_gm[2], \oc8051_golden_model_1.P0 [2]);
  buf(P0_gm[3], \oc8051_golden_model_1.P0 [3]);
  buf(P0_gm[4], \oc8051_golden_model_1.P0 [4]);
  buf(P0_gm[5], \oc8051_golden_model_1.P0 [5]);
  buf(P0_gm[6], \oc8051_golden_model_1.P0 [6]);
  buf(P0_gm[7], \oc8051_golden_model_1.P0 [7]);
  buf(IP_gm_next[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm_next[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm_next[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm_next[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm_next[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm_next[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm_next[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm_next[7], \oc8051_golden_model_1.IP [7]);
  buf(IP_gm[0], \oc8051_golden_model_1.IP [0]);
  buf(IP_gm[1], \oc8051_golden_model_1.IP [1]);
  buf(IP_gm[2], \oc8051_golden_model_1.IP [2]);
  buf(IP_gm[3], \oc8051_golden_model_1.IP [3]);
  buf(IP_gm[4], \oc8051_golden_model_1.IP [4]);
  buf(IP_gm[5], \oc8051_golden_model_1.IP [5]);
  buf(IP_gm[6], \oc8051_golden_model_1.IP [6]);
  buf(IP_gm[7], \oc8051_golden_model_1.IP [7]);
  buf(IE_gm_next[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm_next[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm_next[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm_next[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm_next[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm_next[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm_next[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm_next[7], \oc8051_golden_model_1.IE [7]);
  buf(IE_gm[0], \oc8051_golden_model_1.IE [0]);
  buf(IE_gm[1], \oc8051_golden_model_1.IE [1]);
  buf(IE_gm[2], \oc8051_golden_model_1.IE [2]);
  buf(IE_gm[3], \oc8051_golden_model_1.IE [3]);
  buf(IE_gm[4], \oc8051_golden_model_1.IE [4]);
  buf(IE_gm[5], \oc8051_golden_model_1.IE [5]);
  buf(IE_gm[6], \oc8051_golden_model_1.IE [6]);
  buf(IE_gm[7], \oc8051_golden_model_1.IE [7]);
  buf(DPH_gm[0], \oc8051_golden_model_1.DPH [0]);
  buf(DPH_gm[1], \oc8051_golden_model_1.DPH [1]);
  buf(DPH_gm[2], \oc8051_golden_model_1.DPH [2]);
  buf(DPH_gm[3], \oc8051_golden_model_1.DPH [3]);
  buf(DPH_gm[4], \oc8051_golden_model_1.DPH [4]);
  buf(DPH_gm[5], \oc8051_golden_model_1.DPH [5]);
  buf(DPH_gm[6], \oc8051_golden_model_1.DPH [6]);
  buf(DPH_gm[7], \oc8051_golden_model_1.DPH [7]);
  buf(DPL_gm[0], \oc8051_golden_model_1.DPL [0]);
  buf(DPL_gm[1], \oc8051_golden_model_1.DPL [1]);
  buf(DPL_gm[2], \oc8051_golden_model_1.DPL [2]);
  buf(DPL_gm[3], \oc8051_golden_model_1.DPL [3]);
  buf(DPL_gm[4], \oc8051_golden_model_1.DPL [4]);
  buf(DPL_gm[5], \oc8051_golden_model_1.DPL [5]);
  buf(DPL_gm[6], \oc8051_golden_model_1.DPL [6]);
  buf(DPL_gm[7], \oc8051_golden_model_1.DPL [7]);
  buf(B_gm[0], \oc8051_golden_model_1.B [0]);
  buf(B_gm[1], \oc8051_golden_model_1.B [1]);
  buf(B_gm[2], \oc8051_golden_model_1.B [2]);
  buf(B_gm[3], \oc8051_golden_model_1.B [3]);
  buf(B_gm[4], \oc8051_golden_model_1.B [4]);
  buf(B_gm[5], \oc8051_golden_model_1.B [5]);
  buf(B_gm[6], \oc8051_golden_model_1.B [6]);
  buf(B_gm[7], \oc8051_golden_model_1.B [7]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(PC_gm[0], \oc8051_golden_model_1.PC [0]);
  buf(PC_gm[1], \oc8051_golden_model_1.PC [1]);
  buf(PC_gm[2], \oc8051_golden_model_1.PC [2]);
  buf(PC_gm[3], \oc8051_golden_model_1.PC [3]);
  buf(PC_gm[4], \oc8051_golden_model_1.PC [4]);
  buf(PC_gm[5], \oc8051_golden_model_1.PC [5]);
  buf(PC_gm[6], \oc8051_golden_model_1.PC [6]);
  buf(PC_gm[7], \oc8051_golden_model_1.PC [7]);
  buf(PC_gm[8], \oc8051_golden_model_1.PC [8]);
  buf(PC_gm[9], \oc8051_golden_model_1.PC [9]);
  buf(PC_gm[10], \oc8051_golden_model_1.PC [10]);
  buf(PC_gm[11], \oc8051_golden_model_1.PC [11]);
  buf(PC_gm[12], \oc8051_golden_model_1.PC [12]);
  buf(PC_gm[13], \oc8051_golden_model_1.PC [13]);
  buf(PC_gm[14], \oc8051_golden_model_1.PC [14]);
  buf(PC_gm[15], \oc8051_golden_model_1.PC [15]);
  buf(dptr_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(dptr_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(dptr_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(dptr_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(dptr_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(dptr_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(dptr_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(dptr_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(dptr_impl[8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(dptr_impl[9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(dptr_impl[10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(dptr_impl[11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(dptr_impl[12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(dptr_impl[13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(dptr_impl[14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(dptr_impl[15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(b_reg_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(b_reg_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(b_reg_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(b_reg_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(b_reg_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(b_reg_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(b_reg_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(b_reg_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(acc_impl[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw_impl[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw_impl[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw_impl[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw_impl[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw_impl[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw_impl[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw_impl[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc_impl[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc_impl[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc_impl[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc_impl[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc_impl[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc_impl[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc_impl[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc_impl[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc_impl[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc_impl[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc_impl[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc_impl[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc_impl[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc_impl[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc_impl[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc_impl[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(property_invalid_dec_rom_pc, 1'b0);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
