
module oc8051_xiommu_gm_top(clk, rst, proc_wr, proc_stb, proc_addr, proc_data_in, input_sha_func_0, input_sha_func_1, input_sha_func_2, input_sha_func_3, input_sha_func_4, input_sha_func_5, input_aes_func_6, input_aes_func_7, input_sha_func_8, input_sha_func_9, input_sha_func_10, input_sha_func_11, input_sha_func_12, input_sha_func_13, input_sha_func_14, input_sha_func_15, input_sha_func_16, input_sha_func_17, input_sha_func_18, input_sha_func_19, input_sha_func_20, input_sha_func_21, input_sha_func_22, input_aes_func_23, input_aes_func_24, input_sha_func_25, input_sha_func_26, input_sha_func_27, input_sha_func_28, input_sha_func_29, input_sha_func_30, input_sha_func_31, input_sha_func_32, input_sha_func_33, input_sha_func_34, input_sha_func_35, input_sha_func_36, input_aes_func_37, input_aes_func_38, input_sha_func_39, input_sha_func_40, input_sha_func_41, input_sha_func_42, input_sha_func_43, input_sha_func_44, input_sha_func_45, input_sha_func_46, input_sha_func_47, input_sha_func_48, input_sha_func_49, input_sha_func_50, input_aes_func_51, input_aes_func_52, input_sha_func_53, input_sha_func_54, input_sha_func_55, RD_xram_0, RD_xram_1, RD_xram_2, RD_xram_3, RD_xram_4, RD_xram_5, RD_xram_6, RD_xram_7, RD_xram_8, RD_xram_9, RD_xram_10, RD_xram_11, RD_xram_12, RD_xram_13, RD_xram_14, RD_xram_15, RD_xram_16, RD_xram_17, RD_xram_18, RD_xram_19, RD_xram_20, RD_xram_21, RD_xram_22, RD_xram_23, RD_xram_24, RD_xram_25, RD_xram_26, RD_xram_27, RD_xram_28, RD_xram_29, RD_xram_30, RD_xram_31, RD_xram_32, RD_xram_33, RD_xram_34, RD_xram_35, RD_xram_36, RD_xram_37, RD_xram_38, RD_xram_39, RD_xram_40, RD_xram_41, RD_xram_42, RD_xram_43, RD_xram_44, RD_xram_45, RD_xram_46, RD_xram_47, RD_xram_48, RD_xram_49, RD_xram_50, RD_xram_51, RD_xram_52, RD_xram_53, RD_xram_54, RD_xram_55, RD_xram_56, RD_xram_57, RD_xram_58, RD_xram_59, RD_xram_60, RD_xram_61, RD_xram_62, RD_xram_63, RD_xram_64, RD_xram_65, RD_xram_66, RD_xram_67, RD_xram_68, RD_xram_69, RD_xram_70, RD_xram_71, RD_xram_72, RD_xram_73, RD_xram_74, RD_xram_75, RD_xram_76, RD_xram_77, RD_xram_78, RD_xram_79, RD_xram_80, nondet_memwrite_choice_0, nondet_memwrite_choice_1, nondet_memwrite_choice_2, nondet_memwrite_choice_3, nondet_memwrite_choice_4, nondet_memwrite_choice_5, nondet_memwrite_choice_6, nondet_memwrite_choice_7, nondet_memwrite_choice_8, nondet_memwrite_choice_9, nondet_memwrite_choice_10, nondet_memwrite_choice_11, nondet_memwrite_choice_12, nondet_memwrite_choice_13, nondet_memwrite_choice_14, nondet_memwrite_choice_15, nondet_memwrite_choice_16, nondet_memwrite_choice_17, nondet_memwrite_choice_18, nondet_memwrite_choice_19, nondet_memwrite_choice_20, nondet_memwrite_choice_21, nondet_memwrite_choice_22, nondet_memwrite_choice_23, nondet_memwrite_choice_24, nondet_memwrite_choice_25, nondet_memwrite_choice_26, nondet_memwrite_choice_27, nondet_memwrite_choice_28, nondet_memwrite_choice_29, nondet_memwrite_choice_30, nondet_memwrite_choice_31, nondet_memwrite_choice_32, nondet_memwrite_choice_33, nondet_memwrite_choice_34, nondet_memwrite_choice_35, nondet_memwrite_choice_36, nondet_memwrite_choice_37, nondet_memwrite_choice_38, nondet_memwrite_choice_39, nondet_memwrite_choice_40, nondet_memwrite_choice_41, nondet_memwrite_choice_42, nondet_memwrite_choice_43, nondet_memwrite_choice_44, nondet_memwrite_choice_45, nondet_memwrite_choice_46, nondet_memwrite_choice_47, nondet_memwrite_choice_48, nondet_memwrite_choice_49, nondet_memwrite_choice_50, nondet_memwrite_choice_51, nondet_memwrite_choice_52, nondet_memwrite_choice_53, nondet_memwrite_choice_54, nondet_memwrite_choice_55, nondet_memwrite_choice_56, nondet_memwrite_choice_57, nondet_memwrite_choice_58, nondet_memwrite_choice_59, nondet_memwrite_choice_60, nondet_memwrite_choice_61, nondet_memwrite_choice_62, nondet_memwrite_choice_63, nondet_memwrite_choice_64, nondet_memwrite_choice_65, nondet_memwrite_choice_66, nondet_memwrite_choice_67, nondet_memwrite_choice_68, nondet_memwrite_choice_69, nondet_memwrite_choice_70, nondet_memwrite_choice_71, nondet_memwrite_choice_72, nondet_memwrite_choice_73, nondet_memwrite_choice_74, nondet_memwrite_choice_75, nondet_memwrite_choice_76, nondet_memwrite_choice_77, nondet_memwrite_choice_78, nondet_memwrite_choice_79, nondet_memwrite_choice_80, nondet_memwrite_choice_81, nondet_memwrite_choice_82, nondet_memwrite_choice_83, nondet_memwrite_choice_84, nondet_memwrite_choice_85, nondet_memwrite_choice_86, nondet_memwrite_choice_87, nondet_memwrite_choice_88, nondet_memwrite_choice_89, nondet_memwrite_choice_90, nondet_memwrite_choice_91, nondet_memwrite_choice_92, nondet_memwrite_choice_93, nondet_memwrite_choice_94, nondet_memwrite_choice_95, nondet_memwrite_choice_96, nondet_memwrite_choice_97, nondet_memwrite_choice_98, nondet_memwrite_choice_99, nondet_memwrite_choice_100, nondet_memwrite_choice_101, nondet_memwrite_choice_102, nondet_memwrite_choice_103, nondet_memwrite_choice_104, nondet_memwrite_choice_105, nondet_memwrite_choice_106, nondet_memwrite_choice_107, nondet_memwrite_choice_108, nondet_memwrite_choice_109, nondet_memwrite_choice_110, nondet_memwrite_choice_111, nondet_memwrite_choice_112, nondet_memwrite_choice_113, nondet_memwrite_choice_114, nondet_memwrite_choice_115, nondet_memwrite_choice_116, nondet_memwrite_choice_117, nondet_memwrite_choice_118, nondet_memwrite_choice_119, property_invalid_aes_len, ABINPUT, ABINPUT000);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire _0006_;
  wire _0007_;
  wire _0008_;
  wire _0009_;
  wire _0010_;
  wire _0011_;
  wire _0012_;
  wire _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire _0018_;
  wire _0019_;
  wire _0020_;
  wire _0021_;
  wire _0022_;
  wire _0023_;
  wire _0024_;
  wire _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire _0031_;
  wire _0032_;
  wire _0033_;
  wire _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire _0038_;
  wire _0039_;
  wire _0040_;
  wire _0041_;
  wire _0042_;
  wire _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire _0073_;
  wire _0074_;
  wire _0075_;
  wire _0076_;
  wire _0077_;
  wire _0078_;
  wire _0079_;
  wire _0080_;
  wire _0081_;
  wire _0082_;
  wire _0083_;
  wire _0084_;
  wire _0085_;
  wire _0086_;
  wire _0087_;
  wire _0088_;
  wire _0089_;
  wire _0090_;
  wire _0091_;
  wire _0092_;
  wire _0093_;
  wire _0094_;
  wire _0095_;
  wire _0096_;
  wire _0097_;
  wire _0098_;
  wire _0099_;
  wire _0100_;
  wire _0101_;
  wire _0102_;
  wire _0103_;
  wire _0104_;
  wire _0105_;
  wire _0106_;
  wire _0107_;
  wire _0108_;
  wire _0109_;
  wire _0110_;
  wire _0111_;
  wire _0112_;
  wire _0113_;
  wire _0114_;
  wire _0115_;
  wire _0116_;
  wire _0117_;
  wire _0118_;
  wire _0119_;
  wire _0120_;
  wire _0121_;
  wire _0122_;
  wire _0123_;
  wire _0124_;
  wire _0125_;
  wire _0126_;
  wire _0127_;
  wire _0128_;
  wire _0129_;
  wire _0130_;
  wire _0131_;
  wire _0132_;
  wire _0133_;
  wire _0134_;
  wire _0135_;
  wire _0136_;
  wire _0137_;
  wire _0138_;
  wire _0139_;
  wire _0140_;
  wire _0141_;
  wire _0142_;
  wire _0143_;
  wire _0144_;
  wire _0145_;
  wire _0146_;
  wire _0147_;
  wire _0148_;
  wire _0149_;
  wire _0150_;
  wire _0151_;
  wire _0152_;
  wire _0153_;
  wire _0154_;
  wire _0155_;
  wire _0156_;
  wire _0157_;
  wire _0158_;
  wire _0159_;
  wire _0160_;
  wire _0161_;
  wire _0162_;
  wire _0163_;
  wire _0164_;
  wire _0165_;
  wire _0166_;
  wire _0167_;
  wire _0168_;
  wire _0169_;
  wire _0170_;
  wire _0171_;
  wire _0172_;
  wire _0173_;
  wire _0174_;
  wire _0175_;
  wire _0176_;
  wire _0177_;
  wire _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire _0198_;
  wire _0199_;
  wire _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire _0211_;
  wire _0212_;
  wire _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire _0229_;
  wire _0230_;
  wire _0231_;
  wire _0232_;
  wire _0233_;
  wire _0234_;
  wire _0235_;
  wire _0236_;
  wire _0237_;
  wire _0238_;
  wire _0239_;
  wire _0240_;
  wire _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire _0441_;
  wire _0442_;
  wire _0443_;
  wire _0444_;
  wire _0445_;
  wire _0446_;
  wire _0447_;
  wire _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire _0463_;
  wire _0464_;
  wire _0465_;
  wire _0466_;
  wire _0467_;
  wire _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire _0473_;
  wire _0474_;
  wire _0475_;
  wire _0476_;
  wire _0477_;
  wire _0478_;
  wire _0479_;
  wire _0480_;
  wire _0481_;
  wire _0482_;
  wire _0483_;
  wire _0484_;
  wire _0485_;
  wire _0486_;
  wire _0487_;
  wire _0488_;
  wire _0489_;
  wire _0490_;
  wire _0491_;
  wire _0492_;
  wire _0493_;
  wire _0494_;
  wire _0495_;
  wire _0496_;
  wire _0497_;
  wire _0498_;
  wire _0499_;
  wire _0500_;
  wire _0501_;
  wire _0502_;
  wire _0503_;
  wire _0504_;
  wire _0505_;
  wire _0506_;
  wire _0507_;
  wire _0508_;
  wire _0509_;
  wire _0510_;
  wire _0511_;
  wire _0512_;
  wire _0513_;
  wire _0514_;
  wire _0515_;
  wire _0516_;
  wire _0517_;
  wire _0518_;
  wire _0519_;
  wire _0520_;
  wire _0521_;
  wire _0522_;
  wire _0523_;
  wire _0524_;
  wire _0525_;
  wire _0526_;
  wire _0527_;
  wire _0528_;
  wire _0529_;
  wire _0530_;
  wire _0531_;
  wire _0532_;
  wire _0533_;
  wire _0534_;
  wire _0535_;
  wire _0536_;
  wire _0537_;
  wire _0538_;
  wire _0539_;
  wire _0540_;
  wire _0541_;
  wire _0542_;
  wire _0543_;
  wire _0544_;
  wire _0545_;
  wire _0546_;
  wire _0547_;
  wire _0548_;
  wire _0549_;
  wire _0550_;
  wire _0551_;
  wire _0552_;
  wire _0553_;
  wire _0554_;
  wire _0555_;
  wire _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire _0560_;
  wire _0561_;
  wire _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire _0566_;
  wire _0567_;
  wire _0568_;
  wire _0569_;
  wire _0570_;
  wire _0571_;
  wire _0572_;
  wire _0573_;
  wire _0574_;
  wire _0575_;
  wire _0576_;
  wire _0577_;
  wire _0578_;
  wire _0579_;
  wire _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire _0624_;
  wire _0625_;
  wire _0626_;
  wire _0627_;
  wire _0628_;
  wire _0629_;
  wire _0630_;
  wire _0631_;
  wire _0632_;
  wire _0633_;
  wire _0634_;
  wire _0635_;
  wire _0636_;
  wire _0637_;
  wire _0638_;
  wire _0639_;
  wire _0640_;
  wire _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire _0646_;
  wire _0647_;
  wire _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire _0657_;
  wire _0658_;
  wire _0659_;
  wire _0660_;
  wire _0661_;
  wire _0662_;
  wire _0663_;
  wire _0664_;
  wire _0665_;
  wire _0666_;
  wire _0667_;
  wire _0668_;
  wire _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire _0683_;
  wire _0684_;
  wire _0685_;
  wire _0686_;
  wire _0687_;
  wire _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire _0692_;
  wire _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire _0698_;
  wire _0699_;
  wire _0700_;
  wire _0701_;
  wire _0702_;
  wire _0703_;
  wire _0704_;
  wire _0705_;
  wire _0706_;
  wire _0707_;
  wire _0708_;
  wire _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire _0746_;
  wire _0747_;
  wire _0748_;
  wire _0749_;
  wire _0750_;
  wire _0751_;
  wire _0752_;
  wire _0753_;
  wire _0754_;
  wire _0755_;
  wire _0756_;
  wire _0757_;
  wire _0758_;
  wire _0759_;
  wire _0760_;
  wire _0761_;
  wire _0762_;
  wire _0763_;
  wire _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire _0780_;
  wire _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire _0811_;
  wire _0812_;
  wire _0813_;
  wire _0814_;
  wire _0815_;
  wire _0816_;
  wire _0817_;
  wire _0818_;
  wire _0819_;
  wire _0820_;
  wire _0821_;
  wire _0822_;
  wire _0823_;
  wire _0824_;
  wire _0825_;
  wire _0826_;
  wire _0827_;
  wire _0828_;
  wire _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire _0834_;
  wire _0835_;
  wire _0836_;
  wire _0837_;
  wire _0838_;
  wire _0839_;
  wire _0840_;
  wire _0841_;
  wire _0842_;
  wire _0843_;
  wire _0844_;
  wire _0845_;
  wire _0846_;
  wire _0847_;
  wire _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire _0853_;
  wire _0854_;
  wire _0855_;
  wire _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire _0877_;
  wire _0878_;
  wire _0879_;
  wire _0880_;
  wire _0881_;
  wire _0882_;
  wire _0883_;
  wire _0884_;
  wire _0885_;
  wire _0886_;
  wire _0887_;
  wire _0888_;
  wire _0889_;
  wire _0890_;
  wire _0891_;
  wire _0892_;
  wire _0893_;
  wire _0894_;
  wire _0895_;
  wire _0896_;
  wire _0897_;
  wire _0898_;
  wire _0899_;
  wire _0900_;
  wire _0901_;
  wire _0902_;
  wire _0903_;
  wire _0904_;
  wire _0905_;
  wire _0906_;
  wire _0907_;
  wire _0908_;
  wire _0909_;
  wire _0910_;
  wire _0911_;
  wire _0912_;
  wire _0913_;
  wire _0914_;
  wire _0915_;
  wire _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire _1010_;
  wire _1011_;
  wire _1012_;
  wire _1013_;
  wire _1014_;
  wire _1015_;
  wire _1016_;
  wire _1017_;
  wire _1018_;
  wire _1019_;
  wire _1020_;
  wire _1021_;
  wire _1022_;
  wire _1023_;
  wire _1024_;
  wire _1025_;
  wire _1026_;
  wire _1027_;
  wire _1028_;
  wire _1029_;
  wire _1030_;
  wire _1031_;
  wire _1032_;
  wire _1033_;
  wire _1034_;
  wire _1035_;
  wire _1036_;
  wire _1037_;
  wire _1038_;
  wire _1039_;
  wire _1040_;
  wire _1041_;
  wire _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire _1055_;
  wire _1056_;
  wire _1057_;
  wire _1058_;
  wire _1059_;
  wire _1060_;
  wire _1061_;
  wire _1062_;
  wire _1063_;
  wire _1064_;
  wire _1065_;
  wire _1066_;
  wire _1067_;
  wire _1068_;
  wire _1069_;
  wire _1070_;
  wire _1071_;
  wire _1072_;
  wire _1073_;
  wire _1074_;
  wire _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire _1079_;
  wire _1080_;
  wire _1081_;
  wire _1082_;
  wire _1083_;
  wire _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire _1142_;
  wire _1143_;
  wire _1144_;
  wire _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire _1150_;
  wire _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire _1176_;
  wire _1177_;
  wire _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire _1182_;
  wire _1183_;
  wire _1184_;
  wire _1185_;
  wire _1186_;
  wire _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire _1196_;
  wire _1197_;
  wire _1198_;
  wire _1199_;
  wire _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire _1204_;
  wire _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire _1212_;
  wire _1213_;
  wire _1214_;
  wire _1215_;
  wire _1216_;
  wire _1217_;
  wire _1218_;
  wire _1219_;
  wire _1220_;
  wire _1221_;
  wire _1222_;
  wire _1223_;
  wire _1224_;
  wire _1225_;
  wire _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire _1235_;
  wire _1236_;
  wire _1237_;
  wire _1238_;
  wire _1239_;
  wire _1240_;
  wire _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire _1248_;
  wire _1249_;
  wire _1250_;
  wire _1251_;
  wire _1252_;
  wire _1253_;
  wire _1254_;
  wire _1255_;
  wire _1256_;
  wire _1257_;
  wire _1258_;
  wire _1259_;
  wire _1260_;
  wire _1261_;
  wire _1262_;
  wire _1263_;
  wire _1264_;
  wire _1265_;
  wire _1266_;
  wire _1267_;
  wire _1268_;
  wire _1269_;
  wire _1270_;
  wire _1271_;
  wire _1272_;
  wire _1273_;
  wire _1274_;
  wire _1275_;
  wire _1276_;
  wire _1277_;
  wire _1278_;
  wire _1279_;
  wire _1280_;
  wire _1281_;
  wire _1282_;
  wire _1283_;
  wire _1284_;
  wire _1285_;
  wire _1286_;
  wire _1287_;
  wire _1288_;
  wire _1289_;
  wire _1290_;
  wire _1291_;
  wire _1292_;
  wire _1293_;
  wire _1294_;
  wire _1295_;
  wire _1296_;
  wire _1297_;
  wire _1298_;
  wire _1299_;
  wire _1300_;
  wire _1301_;
  wire _1302_;
  wire _1303_;
  wire _1304_;
  wire _1305_;
  wire _1306_;
  wire _1307_;
  wire _1308_;
  wire _1309_;
  wire _1310_;
  wire _1311_;
  wire _1312_;
  wire _1313_;
  wire _1314_;
  wire _1315_;
  wire _1316_;
  wire _1317_;
  wire _1318_;
  wire _1319_;
  wire _1320_;
  wire _1321_;
  wire _1322_;
  wire _1323_;
  wire _1324_;
  wire _1325_;
  wire _1326_;
  wire _1327_;
  wire _1328_;
  wire _1329_;
  wire _1330_;
  wire _1331_;
  wire _1332_;
  wire _1333_;
  wire _1334_;
  wire _1335_;
  wire _1336_;
  wire _1337_;
  wire _1338_;
  wire _1339_;
  wire _1340_;
  wire _1341_;
  wire _1342_;
  wire _1343_;
  wire _1344_;
  wire _1345_;
  wire _1346_;
  wire _1347_;
  wire _1348_;
  wire _1349_;
  wire _1350_;
  wire _1351_;
  wire _1352_;
  wire _1353_;
  wire _1354_;
  wire _1355_;
  wire _1356_;
  wire _1357_;
  wire _1358_;
  wire _1359_;
  wire _1360_;
  wire _1361_;
  wire _1362_;
  wire _1363_;
  wire _1364_;
  wire _1365_;
  wire _1366_;
  wire _1367_;
  wire _1368_;
  wire _1369_;
  wire _1370_;
  wire _1371_;
  wire _1372_;
  wire _1373_;
  wire _1374_;
  wire _1375_;
  wire _1376_;
  wire _1377_;
  wire _1378_;
  wire _1379_;
  wire _1380_;
  wire _1381_;
  wire _1382_;
  wire _1383_;
  wire _1384_;
  wire _1385_;
  wire _1386_;
  wire _1387_;
  wire _1388_;
  wire _1389_;
  wire _1390_;
  wire _1391_;
  wire _1392_;
  wire _1393_;
  wire _1394_;
  wire _1395_;
  wire _1396_;
  wire _1397_;
  wire _1398_;
  wire _1399_;
  wire _1400_;
  wire _1401_;
  wire _1402_;
  wire _1403_;
  wire _1404_;
  wire _1405_;
  wire _1406_;
  wire _1407_;
  wire _1408_;
  wire _1409_;
  wire _1410_;
  wire _1411_;
  wire _1412_;
  wire _1413_;
  wire _1414_;
  wire _1415_;
  wire _1416_;
  wire _1417_;
  wire _1418_;
  wire _1419_;
  wire _1420_;
  wire _1421_;
  wire _1422_;
  wire _1423_;
  wire _1424_;
  wire _1425_;
  wire _1426_;
  wire _1427_;
  wire _1428_;
  wire _1429_;
  wire _1430_;
  wire _1431_;
  wire _1432_;
  wire _1433_;
  wire _1434_;
  wire _1435_;
  wire _1436_;
  wire _1437_;
  wire _1438_;
  wire _1439_;
  wire _1440_;
  wire _1441_;
  wire _1442_;
  wire _1443_;
  wire _1444_;
  wire _1445_;
  wire _1446_;
  wire _1447_;
  wire _1448_;
  wire _1449_;
  wire _1450_;
  wire _1451_;
  wire _1452_;
  wire _1453_;
  wire _1454_;
  wire _1455_;
  wire _1456_;
  wire _1457_;
  wire _1458_;
  wire _1459_;
  wire _1460_;
  wire _1461_;
  wire _1462_;
  wire _1463_;
  wire _1464_;
  wire _1465_;
  wire _1466_;
  wire _1467_;
  wire _1468_;
  wire _1469_;
  wire _1470_;
  wire _1471_;
  wire _1472_;
  wire _1473_;
  wire _1474_;
  wire _1475_;
  wire _1476_;
  wire _1477_;
  wire _1478_;
  wire _1479_;
  wire _1480_;
  wire _1481_;
  wire _1482_;
  wire _1483_;
  wire _1484_;
  wire _1485_;
  wire _1486_;
  wire _1487_;
  wire _1488_;
  wire _1489_;
  wire _1490_;
  wire _1491_;
  wire _1492_;
  wire _1493_;
  wire _1494_;
  wire _1495_;
  wire _1496_;
  wire _1497_;
  wire _1498_;
  wire _1499_;
  wire _1500_;
  wire _1501_;
  wire _1502_;
  wire _1503_;
  wire _1504_;
  wire _1505_;
  wire _1506_;
  wire _1507_;
  wire _1508_;
  wire _1509_;
  wire _1510_;
  wire _1511_;
  wire _1512_;
  wire _1513_;
  wire _1514_;
  wire _1515_;
  wire _1516_;
  wire _1517_;
  wire _1518_;
  wire _1519_;
  wire _1520_;
  wire _1521_;
  wire _1522_;
  wire _1523_;
  wire _1524_;
  wire _1525_;
  wire _1526_;
  wire _1527_;
  wire _1528_;
  wire _1529_;
  wire _1530_;
  wire _1531_;
  wire _1532_;
  wire _1533_;
  wire _1534_;
  wire _1535_;
  wire _1536_;
  wire _1537_;
  wire _1538_;
  wire _1539_;
  wire _1540_;
  wire _1541_;
  wire _1542_;
  wire _1543_;
  wire _1544_;
  wire _1545_;
  wire _1546_;
  wire _1547_;
  wire _1548_;
  wire _1549_;
  wire _1550_;
  wire _1551_;
  wire _1552_;
  wire _1553_;
  wire _1554_;
  wire _1555_;
  wire _1556_;
  wire _1557_;
  wire _1558_;
  wire _1559_;
  wire _1560_;
  wire _1561_;
  wire _1562_;
  wire _1563_;
  wire _1564_;
  wire _1565_;
  wire _1566_;
  wire _1567_;
  wire _1568_;
  wire _1569_;
  wire _1570_;
  wire _1571_;
  wire _1572_;
  wire _1573_;
  wire _1574_;
  wire _1575_;
  wire _1576_;
  wire _1577_;
  wire _1578_;
  wire _1579_;
  wire _1580_;
  wire _1581_;
  wire _1582_;
  wire _1583_;
  wire _1584_;
  wire _1585_;
  wire _1586_;
  wire _1587_;
  wire _1588_;
  wire _1589_;
  wire _1590_;
  wire _1591_;
  wire _1592_;
  wire _1593_;
  wire _1594_;
  wire _1595_;
  wire _1596_;
  wire _1597_;
  wire _1598_;
  wire _1599_;
  wire _1600_;
  wire _1601_;
  wire _1602_;
  wire _1603_;
  wire _1604_;
  wire _1605_;
  wire _1606_;
  wire _1607_;
  wire _1608_;
  wire _1609_;
  wire _1610_;
  wire _1611_;
  wire _1612_;
  wire _1613_;
  wire _1614_;
  wire _1615_;
  wire _1616_;
  wire _1617_;
  wire _1618_;
  wire _1619_;
  wire _1620_;
  wire _1621_;
  wire _1622_;
  wire _1623_;
  wire _1624_;
  wire _1625_;
  wire _1626_;
  wire _1627_;
  wire _1628_;
  wire _1629_;
  wire _1630_;
  wire _1631_;
  wire _1632_;
  wire _1633_;
  wire _1634_;
  wire _1635_;
  wire _1636_;
  wire _1637_;
  wire _1638_;
  wire _1639_;
  wire _1640_;
  wire _1641_;
  wire _1642_;
  wire _1643_;
  wire _1644_;
  wire _1645_;
  wire _1646_;
  wire _1647_;
  wire _1648_;
  wire _1649_;
  wire _1650_;
  wire _1651_;
  wire _1652_;
  wire _1653_;
  wire _1654_;
  wire _1655_;
  wire _1656_;
  wire _1657_;
  wire _1658_;
  wire _1659_;
  wire _1660_;
  wire _1661_;
  wire _1662_;
  wire _1663_;
  wire _1664_;
  wire _1665_;
  wire _1666_;
  wire _1667_;
  wire _1668_;
  wire _1669_;
  wire _1670_;
  wire _1671_;
  wire _1672_;
  wire _1673_;
  wire _1674_;
  wire _1675_;
  wire _1676_;
  wire _1677_;
  wire _1678_;
  wire _1679_;
  wire _1680_;
  wire _1681_;
  wire _1682_;
  wire _1683_;
  wire _1684_;
  wire _1685_;
  wire _1686_;
  wire _1687_;
  wire _1688_;
  wire _1689_;
  wire _1690_;
  wire _1691_;
  wire _1692_;
  wire _1693_;
  wire _1694_;
  wire _1695_;
  wire _1696_;
  wire _1697_;
  wire _1698_;
  wire _1699_;
  wire _1700_;
  wire _1701_;
  wire _1702_;
  wire _1703_;
  wire _1704_;
  wire _1705_;
  wire _1706_;
  wire _1707_;
  wire _1708_;
  wire _1709_;
  wire _1710_;
  wire _1711_;
  wire _1712_;
  wire _1713_;
  wire _1714_;
  wire _1715_;
  wire _1716_;
  wire _1717_;
  wire _1718_;
  wire _1719_;
  wire _1720_;
  wire _1721_;
  wire _1722_;
  wire _1723_;
  wire _1724_;
  wire _1725_;
  wire _1726_;
  wire _1727_;
  wire _1728_;
  wire _1729_;
  wire _1730_;
  wire _1731_;
  wire _1732_;
  wire _1733_;
  wire _1734_;
  wire _1735_;
  wire _1736_;
  wire _1737_;
  wire _1738_;
  wire _1739_;
  wire _1740_;
  wire _1741_;
  wire _1742_;
  wire _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  wire _1750_;
  wire _1751_;
  wire _1752_;
  wire _1753_;
  wire _1754_;
  wire _1755_;
  wire _1756_;
  wire _1757_;
  wire _1758_;
  wire _1759_;
  wire _1760_;
  wire _1761_;
  wire _1762_;
  wire _1763_;
  wire _1764_;
  wire _1765_;
  wire _1766_;
  wire _1767_;
  wire _1768_;
  wire _1769_;
  wire _1770_;
  wire _1771_;
  wire _1772_;
  wire _1773_;
  wire _1774_;
  wire _1775_;
  wire _1776_;
  wire _1777_;
  wire _1778_;
  wire _1779_;
  wire _1780_;
  wire _1781_;
  wire _1782_;
  wire _1783_;
  wire _1784_;
  wire _1785_;
  wire _1786_;
  wire _1787_;
  wire _1788_;
  wire _1789_;
  wire _1790_;
  wire _1791_;
  wire _1792_;
  wire _1793_;
  wire _1794_;
  wire _1795_;
  wire _1796_;
  wire _1797_;
  wire _1798_;
  wire _1799_;
  wire _1800_;
  wire _1801_;
  wire _1802_;
  wire _1803_;
  wire _1804_;
  wire _1805_;
  wire _1806_;
  wire _1807_;
  wire _1808_;
  wire _1809_;
  wire _1810_;
  wire _1811_;
  wire _1812_;
  wire _1813_;
  wire _1814_;
  wire _1815_;
  wire _1816_;
  wire _1817_;
  wire _1818_;
  wire _1819_;
  wire _1820_;
  wire _1821_;
  wire _1822_;
  wire _1823_;
  wire _1824_;
  wire _1825_;
  wire _1826_;
  wire _1827_;
  wire _1828_;
  wire _1829_;
  wire _1830_;
  wire _1831_;
  wire _1832_;
  wire _1833_;
  wire _1834_;
  wire _1835_;
  wire _1836_;
  wire _1837_;
  wire _1838_;
  wire _1839_;
  wire _1840_;
  wire _1841_;
  wire _1842_;
  wire _1843_;
  wire _1844_;
  wire _1845_;
  wire _1846_;
  wire _1847_;
  wire _1848_;
  wire _1849_;
  wire _1850_;
  wire _1851_;
  wire _1852_;
  wire _1853_;
  wire _1854_;
  wire _1855_;
  wire _1856_;
  wire _1857_;
  wire _1858_;
  wire _1859_;
  wire _1860_;
  wire _1861_;
  wire _1862_;
  wire _1863_;
  wire _1864_;
  wire _1865_;
  wire _1866_;
  wire _1867_;
  wire _1868_;
  wire _1869_;
  wire _1870_;
  wire _1871_;
  wire _1872_;
  wire _1873_;
  wire _1874_;
  wire _1875_;
  wire _1876_;
  wire _1877_;
  wire _1878_;
  wire _1879_;
  wire _1880_;
  wire _1881_;
  wire _1882_;
  wire _1883_;
  wire _1884_;
  wire _1885_;
  wire _1886_;
  wire _1887_;
  wire _1888_;
  wire _1889_;
  wire _1890_;
  wire _1891_;
  wire [15:0] _1892_;
  wire [15:0] _1893_;
  wire [7:0] _1894_;
  wire [15:0] _1895_;
  wire [15:0] _1896_;
  wire [7:0] _1897_;
  input [127:0] ABINPUT;
  input [161:0] ABINPUT000;
  input [7:0] RD_xram_0;
  input [7:0] RD_xram_1;
  input [7:0] RD_xram_10;
  input [7:0] RD_xram_11;
  input [7:0] RD_xram_12;
  input [7:0] RD_xram_13;
  input [7:0] RD_xram_14;
  input [7:0] RD_xram_15;
  input [7:0] RD_xram_16;
  input [7:0] RD_xram_17;
  input [7:0] RD_xram_18;
  input [7:0] RD_xram_19;
  input [7:0] RD_xram_2;
  input [7:0] RD_xram_20;
  input [7:0] RD_xram_21;
  input [7:0] RD_xram_22;
  input [7:0] RD_xram_23;
  input [7:0] RD_xram_24;
  input [7:0] RD_xram_25;
  input [7:0] RD_xram_26;
  input [7:0] RD_xram_27;
  input [7:0] RD_xram_28;
  input [7:0] RD_xram_29;
  input [7:0] RD_xram_3;
  input [7:0] RD_xram_30;
  input [7:0] RD_xram_31;
  input [7:0] RD_xram_32;
  input [7:0] RD_xram_33;
  input [7:0] RD_xram_34;
  input [7:0] RD_xram_35;
  input [7:0] RD_xram_36;
  input [7:0] RD_xram_37;
  input [7:0] RD_xram_38;
  input [7:0] RD_xram_39;
  input [7:0] RD_xram_4;
  input [7:0] RD_xram_40;
  input [7:0] RD_xram_41;
  input [7:0] RD_xram_42;
  input [7:0] RD_xram_43;
  input [7:0] RD_xram_44;
  input [7:0] RD_xram_45;
  input [7:0] RD_xram_46;
  input [7:0] RD_xram_47;
  input [7:0] RD_xram_48;
  input [7:0] RD_xram_49;
  input [7:0] RD_xram_5;
  input [7:0] RD_xram_50;
  input [7:0] RD_xram_51;
  input [7:0] RD_xram_52;
  input [7:0] RD_xram_53;
  input [7:0] RD_xram_54;
  input [7:0] RD_xram_55;
  input [7:0] RD_xram_56;
  input [7:0] RD_xram_57;
  input [7:0] RD_xram_58;
  input [7:0] RD_xram_59;
  input [7:0] RD_xram_6;
  input [7:0] RD_xram_60;
  input [7:0] RD_xram_61;
  input [7:0] RD_xram_62;
  input [7:0] RD_xram_63;
  input [7:0] RD_xram_64;
  input [7:0] RD_xram_65;
  input [7:0] RD_xram_66;
  input [7:0] RD_xram_67;
  input [7:0] RD_xram_68;
  input [7:0] RD_xram_69;
  input [7:0] RD_xram_7;
  input [7:0] RD_xram_70;
  input [7:0] RD_xram_71;
  input [7:0] RD_xram_72;
  input [7:0] RD_xram_73;
  input [7:0] RD_xram_74;
  input [7:0] RD_xram_75;
  input [7:0] RD_xram_76;
  input [7:0] RD_xram_77;
  input [7:0] RD_xram_78;
  input [7:0] RD_xram_79;
  input [7:0] RD_xram_8;
  input [7:0] RD_xram_80;
  input [7:0] RD_xram_9;
  wire [15:0] addrin;
  wire [15:0] aes_addr_gm;
  wire [15:0] aes_len_gm;
  wire [15:0] aes_len_impl;
  wire [7:0] aes_state_gm;
  wire [1:0] aes_state_impl;
  input clk;
  wire [7:0] datain;
  input [63:0] input_aes_func_23;
  input [63:0] input_aes_func_24;
  input [63:0] input_aes_func_37;
  input [63:0] input_aes_func_38;
  input [63:0] input_aes_func_51;
  input [63:0] input_aes_func_52;
  input [63:0] input_aes_func_6;
  input [63:0] input_aes_func_7;
  input [63:0] input_sha_func_0;
  input [63:0] input_sha_func_1;
  input [31:0] input_sha_func_10;
  input [63:0] input_sha_func_11;
  input [63:0] input_sha_func_12;
  input [31:0] input_sha_func_13;
  input [63:0] input_sha_func_14;
  input [63:0] input_sha_func_15;
  input [31:0] input_sha_func_16;
  input [63:0] input_sha_func_17;
  input [63:0] input_sha_func_18;
  input [31:0] input_sha_func_19;
  input [31:0] input_sha_func_2;
  input [63:0] input_sha_func_20;
  input [63:0] input_sha_func_21;
  input [31:0] input_sha_func_22;
  input [63:0] input_sha_func_25;
  input [63:0] input_sha_func_26;
  input [31:0] input_sha_func_27;
  input [63:0] input_sha_func_28;
  input [63:0] input_sha_func_29;
  input [63:0] input_sha_func_3;
  input [31:0] input_sha_func_30;
  input [63:0] input_sha_func_31;
  input [63:0] input_sha_func_32;
  input [31:0] input_sha_func_33;
  input [63:0] input_sha_func_34;
  input [63:0] input_sha_func_35;
  input [31:0] input_sha_func_36;
  input [63:0] input_sha_func_39;
  input [63:0] input_sha_func_4;
  input [63:0] input_sha_func_40;
  input [31:0] input_sha_func_41;
  input [63:0] input_sha_func_42;
  input [63:0] input_sha_func_43;
  input [31:0] input_sha_func_44;
  input [63:0] input_sha_func_45;
  input [63:0] input_sha_func_46;
  input [31:0] input_sha_func_47;
  input [63:0] input_sha_func_48;
  input [63:0] input_sha_func_49;
  input [31:0] input_sha_func_5;
  input [31:0] input_sha_func_50;
  input [63:0] input_sha_func_53;
  input [63:0] input_sha_func_54;
  input [31:0] input_sha_func_55;
  input [63:0] input_sha_func_8;
  input [63:0] input_sha_func_9;
  input nondet_memwrite_choice_0;
  input nondet_memwrite_choice_1;
  input nondet_memwrite_choice_10;
  input nondet_memwrite_choice_100;
  input nondet_memwrite_choice_101;
  input nondet_memwrite_choice_102;
  input nondet_memwrite_choice_103;
  input nondet_memwrite_choice_104;
  input nondet_memwrite_choice_105;
  input nondet_memwrite_choice_106;
  input nondet_memwrite_choice_107;
  input nondet_memwrite_choice_108;
  input nondet_memwrite_choice_109;
  input nondet_memwrite_choice_11;
  input nondet_memwrite_choice_110;
  input nondet_memwrite_choice_111;
  input nondet_memwrite_choice_112;
  input nondet_memwrite_choice_113;
  input nondet_memwrite_choice_114;
  input nondet_memwrite_choice_115;
  input nondet_memwrite_choice_116;
  input nondet_memwrite_choice_117;
  input nondet_memwrite_choice_118;
  input nondet_memwrite_choice_119;
  input nondet_memwrite_choice_12;
  input nondet_memwrite_choice_13;
  input nondet_memwrite_choice_14;
  input nondet_memwrite_choice_15;
  input nondet_memwrite_choice_16;
  input nondet_memwrite_choice_17;
  input nondet_memwrite_choice_18;
  input nondet_memwrite_choice_19;
  input nondet_memwrite_choice_2;
  input nondet_memwrite_choice_20;
  input nondet_memwrite_choice_21;
  input nondet_memwrite_choice_22;
  input nondet_memwrite_choice_23;
  input nondet_memwrite_choice_24;
  input nondet_memwrite_choice_25;
  input nondet_memwrite_choice_26;
  input nondet_memwrite_choice_27;
  input nondet_memwrite_choice_28;
  input nondet_memwrite_choice_29;
  input nondet_memwrite_choice_3;
  input nondet_memwrite_choice_30;
  input nondet_memwrite_choice_31;
  input nondet_memwrite_choice_32;
  input nondet_memwrite_choice_33;
  input nondet_memwrite_choice_34;
  input nondet_memwrite_choice_35;
  input nondet_memwrite_choice_36;
  input nondet_memwrite_choice_37;
  input nondet_memwrite_choice_38;
  input nondet_memwrite_choice_39;
  input nondet_memwrite_choice_4;
  input nondet_memwrite_choice_40;
  input nondet_memwrite_choice_41;
  input nondet_memwrite_choice_42;
  input nondet_memwrite_choice_43;
  input nondet_memwrite_choice_44;
  input nondet_memwrite_choice_45;
  input nondet_memwrite_choice_46;
  input nondet_memwrite_choice_47;
  input nondet_memwrite_choice_48;
  input nondet_memwrite_choice_49;
  input nondet_memwrite_choice_5;
  input nondet_memwrite_choice_50;
  input nondet_memwrite_choice_51;
  input nondet_memwrite_choice_52;
  input nondet_memwrite_choice_53;
  input nondet_memwrite_choice_54;
  input nondet_memwrite_choice_55;
  input nondet_memwrite_choice_56;
  input nondet_memwrite_choice_57;
  input nondet_memwrite_choice_58;
  input nondet_memwrite_choice_59;
  input nondet_memwrite_choice_6;
  input nondet_memwrite_choice_60;
  input nondet_memwrite_choice_61;
  input nondet_memwrite_choice_62;
  input nondet_memwrite_choice_63;
  input nondet_memwrite_choice_64;
  input nondet_memwrite_choice_65;
  input nondet_memwrite_choice_66;
  input nondet_memwrite_choice_67;
  input nondet_memwrite_choice_68;
  input nondet_memwrite_choice_69;
  input nondet_memwrite_choice_7;
  input nondet_memwrite_choice_70;
  input nondet_memwrite_choice_71;
  input nondet_memwrite_choice_72;
  input nondet_memwrite_choice_73;
  input nondet_memwrite_choice_74;
  input nondet_memwrite_choice_75;
  input nondet_memwrite_choice_76;
  input nondet_memwrite_choice_77;
  input nondet_memwrite_choice_78;
  input nondet_memwrite_choice_79;
  input nondet_memwrite_choice_8;
  input nondet_memwrite_choice_80;
  input nondet_memwrite_choice_81;
  input nondet_memwrite_choice_82;
  input nondet_memwrite_choice_83;
  input nondet_memwrite_choice_84;
  input nondet_memwrite_choice_85;
  input nondet_memwrite_choice_86;
  input nondet_memwrite_choice_87;
  input nondet_memwrite_choice_88;
  input nondet_memwrite_choice_89;
  input nondet_memwrite_choice_9;
  input nondet_memwrite_choice_90;
  input nondet_memwrite_choice_91;
  input nondet_memwrite_choice_92;
  input nondet_memwrite_choice_93;
  input nondet_memwrite_choice_94;
  input nondet_memwrite_choice_95;
  input nondet_memwrite_choice_96;
  input nondet_memwrite_choice_97;
  input nondet_memwrite_choice_98;
  input nondet_memwrite_choice_99;
  wire [127:0] \oc8051_xiommu_impl_1.ABINPUT ;
  wire [161:0] \oc8051_xiommu_impl_1.ABINPUT000 ;
  wire [15:0] \oc8051_xiommu_impl_1.aes_len ;
  wire [1:0] \oc8051_xiommu_impl_1.aes_state ;
  wire [127:0] \oc8051_xiommu_impl_1.aes_top_i.ABINPUT ;
  wire [15:0] \oc8051_xiommu_impl_1.aes_top_i.addr ;
  wire [15:0] \oc8051_xiommu_impl_1.aes_top_i.aes_len ;
  wire [127:0] \oc8051_xiommu_impl_1.aes_top_i.aes_out ;
  wire [3:0] \oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.addr ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.clk ;
  wire [7:0] \oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.data_in ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.rst ;
  wire [3:0] \oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.addr ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.clk ;
  wire [7:0] \oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.data_in ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.rst ;
  wire [3:0] \oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.addr ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.clk ;
  wire [7:0] \oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.data_in ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.rst ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.addr ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.clk ;
  wire [7:0] \oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.data_in ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.rst ;
  wire [15:0] \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.addr ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.clk ;
  wire [7:0] \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.data_in ;
  wire [15:0] \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out ;
  wire \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.rst ;
  wire [1:0] \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state ;
  wire [1:0] \oc8051_xiommu_impl_1.aes_top_i.aes_state ;
  wire [3:0] \oc8051_xiommu_impl_1.aes_top_i.byte_counter ;
  wire \oc8051_xiommu_impl_1.aes_top_i.clk ;
  wire [7:0] \oc8051_xiommu_impl_1.aes_top_i.data_in ;
  wire [15:0] \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count ;
  wire \oc8051_xiommu_impl_1.aes_top_i.rst ;
  wire \oc8051_xiommu_impl_1.clk ;
  wire [15:0] \oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A ;
  wire [1:0] \oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbit_holder ;
  wire \oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbiter_state ;
  wire \oc8051_xiommu_impl_1.oc8051_memarbiter_i.clk ;
  wire [7:0] \oc8051_xiommu_impl_1.oc8051_memarbiter_i.data_in_A ;
  wire \oc8051_xiommu_impl_1.oc8051_memarbiter_i.rst ;
  wire \oc8051_xiommu_impl_1.oc8051_xram_i.ackr ;
  wire \oc8051_xiommu_impl_1.oc8051_xram_i.ackw ;
  wire \oc8051_xiommu_impl_1.oc8051_xram_i.clk ;
  wire [2:0] \oc8051_xiommu_impl_1.oc8051_xram_i.cnt ;
  wire \oc8051_xiommu_impl_1.oc8051_xram_i.rst ;
  wire [15:0] \oc8051_xiommu_impl_1.proc_addr ;
  wire [7:0] \oc8051_xiommu_impl_1.proc_data_in ;
  wire \oc8051_xiommu_impl_1.proc_stb ;
  wire \oc8051_xiommu_impl_1.proc_wr ;
  wire \oc8051_xiommu_impl_1.rst ;
  wire [15:0] \oc8051_xiommu_impl_1.sha_len ;
  wire [1:0] \oc8051_xiommu_impl_1.sha_state ;
  wire [161:0] \oc8051_xiommu_impl_1.sha_top_i.ABINPUT ;
  wire [15:0] \oc8051_xiommu_impl_1.sha_top_i.addr ;
  wire [5:0] \oc8051_xiommu_impl_1.sha_top_i.byte_counter ;
  wire \oc8051_xiommu_impl_1.sha_top_i.clk ;
  wire [7:0] \oc8051_xiommu_impl_1.sha_top_i.data_in ;
  wire [7:0] \oc8051_xiommu_impl_1.sha_top_i.data_out_state ;
  wire [15:0] \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read ;
  wire \oc8051_xiommu_impl_1.sha_top_i.rst ;
  wire [159:0] \oc8051_xiommu_impl_1.sha_top_i.sha_core_digest ;
  wire \oc8051_xiommu_impl_1.sha_top_i.sha_core_digest_valid ;
  wire \oc8051_xiommu_impl_1.sha_top_i.sha_core_ready ;
  wire [15:0] \oc8051_xiommu_impl_1.sha_top_i.sha_len ;
  wire [15:0] \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len ;
  wire \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.addr ;
  wire \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.clk ;
  wire [7:0] \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.data_in ;
  wire [15:0] \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out ;
  wire \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.rst ;
  wire \oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.addr ;
  wire \oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.clk ;
  wire [7:0] \oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.data_in ;
  wire \oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.rst ;
  wire [1:0] \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state ;
  wire \oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.addr ;
  wire \oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.clk ;
  wire [7:0] \oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.data_in ;
  wire \oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.rst ;
  wire [1:0] \oc8051_xiommu_impl_1.sha_top_i.sha_state ;
  input [15:0] proc_addr;
  input [7:0] proc_data_in;
  input proc_stb;
  wire proc_stb_r;
  wire proc_stb_valid;
  input proc_wr;
  output property_invalid_aes_len;
  input rst;
  wire [15:0] sha_len_gm;
  wire [15:0] sha_len_impl;
  wire [15:0] sha_rdaddr_gm;
  wire [7:0] sha_state_gm;
  wire [1:0] sha_state_impl;
  wire [15:0] sha_wraddr_gm;
  wire [7:0] \xm8051_golden_model_1.RD_xram_0 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_1 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_10 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_11 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_12 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_13 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_14 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_15 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_16 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_17 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_18 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_19 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_2 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_20 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_21 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_22 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_23 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_24 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_25 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_26 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_27 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_28 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_29 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_3 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_30 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_31 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_32 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_33 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_34 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_35 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_36 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_37 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_38 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_39 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_4 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_40 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_41 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_42 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_43 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_44 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_45 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_46 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_47 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_48 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_49 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_5 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_50 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_51 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_52 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_53 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_54 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_55 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_56 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_57 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_58 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_59 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_6 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_60 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_61 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_62 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_63 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_64 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_65 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_66 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_67 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_68 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_69 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_7 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_70 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_71 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_72 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_73 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_74 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_75 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_76 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_77 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_78 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_79 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_8 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_80 ;
  wire [7:0] \xm8051_golden_model_1.RD_xram_9 ;
  wire [15:0] \xm8051_golden_model_1.WR_XRAM_ADDR_00 ;
  wire [15:0] \xm8051_golden_model_1.WR_XRAM_ADDR_01 ;
  wire [15:0] \xm8051_golden_model_1.WR_XRAM_ADDR_02 ;
  wire [15:0] \xm8051_golden_model_1.WR_XRAM_ADDR_04 ;
  wire [15:0] \xm8051_golden_model_1.WR_XRAM_ADDR_05 ;
  wire [15:0] \xm8051_golden_model_1.WR_XRAM_ADDR_06 ;
  wire [15:0] \xm8051_golden_model_1.WR_XRAM_ADDR_08 ;
  wire [15:0] \xm8051_golden_model_1.WR_XRAM_ADDR_09 ;
  wire [15:0] \xm8051_golden_model_1.WR_XRAM_ADDR_0a ;
  wire [15:0] \xm8051_golden_model_1.WR_XRAM_ADDR_0c ;
  wire [15:0] \xm8051_golden_model_1.WR_XRAM_ADDR_0e ;
  wire [15:0] \xm8051_golden_model_1.addrin ;
  wire [15:0] \xm8051_golden_model_1.aes_bytes_processed ;
  wire [15:0] \xm8051_golden_model_1.aes_bytes_processed_03 ;
  wire [15:0] \xm8051_golden_model_1.aes_bytes_processed_07 ;
  wire [15:0] \xm8051_golden_model_1.aes_bytes_processed_0b ;
  wire [15:0] \xm8051_golden_model_1.aes_bytes_processed_0f ;
  wire [15:0] \xm8051_golden_model_1.aes_len ;
  wire [7:0] \xm8051_golden_model_1.aes_state ;
  wire \xm8051_golden_model_1.clk ;
  wire [7:0] \xm8051_golden_model_1.datain ;
  wire [63:0] \xm8051_golden_model_1.input_aes_func_23 ;
  wire [63:0] \xm8051_golden_model_1.input_aes_func_24 ;
  wire [63:0] \xm8051_golden_model_1.input_aes_func_37 ;
  wire [63:0] \xm8051_golden_model_1.input_aes_func_38 ;
  wire [63:0] \xm8051_golden_model_1.input_aes_func_51 ;
  wire [63:0] \xm8051_golden_model_1.input_aes_func_52 ;
  wire [63:0] \xm8051_golden_model_1.input_aes_func_6 ;
  wire [63:0] \xm8051_golden_model_1.input_aes_func_7 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_0 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_1 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_10 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_11 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_12 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_13 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_14 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_15 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_16 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_17 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_18 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_19 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_2 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_20 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_21 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_22 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_25 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_26 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_27 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_28 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_29 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_3 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_30 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_31 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_32 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_33 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_34 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_35 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_36 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_39 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_4 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_40 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_41 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_42 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_43 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_44 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_45 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_46 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_47 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_48 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_49 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_5 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_50 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_53 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_54 ;
  wire [31:0] \xm8051_golden_model_1.input_sha_func_55 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_8 ;
  wire [63:0] \xm8051_golden_model_1.input_sha_func_9 ;
  wire [1:0] \xm8051_golden_model_1.n0001 ;
  wire [1:0] \xm8051_golden_model_1.n0002 ;
  wire [3:0] \xm8051_golden_model_1.n0003 ;
  wire [15:0] \xm8051_golden_model_1.n0037 ;
  wire [15:0] \xm8051_golden_model_1.n0055 ;
  wire [15:0] \xm8051_golden_model_1.n0064 ;
  wire [15:0] \xm8051_golden_model_1.n0077 ;
  wire [15:0] \xm8051_golden_model_1.n0086 ;
  wire [15:0] \xm8051_golden_model_1.n0099 ;
  wire [15:0] \xm8051_golden_model_1.n0108 ;
  wire [15:0] \xm8051_golden_model_1.n0121 ;
  wire [15:0] \xm8051_golden_model_1.n0130 ;
  wire [15:0] \xm8051_golden_model_1.n0143 ;
  wire [15:0] \xm8051_golden_model_1.n0152 ;
  wire [15:0] \xm8051_golden_model_1.n0165 ;
  wire [15:0] \xm8051_golden_model_1.n0174 ;
  wire [15:0] \xm8051_golden_model_1.n0187 ;
  wire [15:0] \xm8051_golden_model_1.n0196 ;
  wire [15:0] \xm8051_golden_model_1.n0209 ;
  wire [15:0] \xm8051_golden_model_1.n0218 ;
  wire [15:0] \xm8051_golden_model_1.n0233 ;
  wire [15:0] \xm8051_golden_model_1.n0245 ;
  wire [15:0] \xm8051_golden_model_1.n0257 ;
  wire [15:0] \xm8051_golden_model_1.n0269 ;
  wire [15:0] \xm8051_golden_model_1.n0281 ;
  wire [15:0] \xm8051_golden_model_1.n0293 ;
  wire [15:0] \xm8051_golden_model_1.n0305 ;
  wire [15:0] \xm8051_golden_model_1.n0317 ;
  wire [15:0] \xm8051_golden_model_1.n0329 ;
  wire [15:0] \xm8051_golden_model_1.n0341 ;
  wire [15:0] \xm8051_golden_model_1.n0353 ;
  wire [15:0] \xm8051_golden_model_1.n0365 ;
  wire [15:0] \xm8051_golden_model_1.n0377 ;
  wire [15:0] \xm8051_golden_model_1.n0389 ;
  wire [15:0] \xm8051_golden_model_1.n0401 ;
  wire [15:0] \xm8051_golden_model_1.n0413 ;
  wire [15:0] \xm8051_golden_model_1.n0423 ;
  wire [15:0] \xm8051_golden_model_1.n0433 ;
  wire [15:0] \xm8051_golden_model_1.n0443 ;
  wire [15:0] \xm8051_golden_model_1.n0453 ;
  wire [15:0] \xm8051_golden_model_1.n0463 ;
  wire [15:0] \xm8051_golden_model_1.n0473 ;
  wire [15:0] \xm8051_golden_model_1.n0483 ;
  wire [15:0] \xm8051_golden_model_1.n0493 ;
  wire [14:0] \xm8051_golden_model_1.n0510 ;
  wire [15:0] \xm8051_golden_model_1.n0512 ;
  wire \xm8051_golden_model_1.n0515 ;
  wire [7:0] \xm8051_golden_model_1.n0523 ;
  wire [7:0] \xm8051_golden_model_1.n0524 ;
  wire [11:0] \xm8051_golden_model_1.n0527 ;
  wire [15:0] \xm8051_golden_model_1.n0529 ;
  wire [3:0] \xm8051_golden_model_1.n0532 ;
  wire [7:0] \xm8051_golden_model_1.n0690 ;
  wire [7:0] \xm8051_golden_model_1.n0691 ;
  wire [15:0] \xm8051_golden_model_1.n0703 ;
  wire [15:0] \xm8051_golden_model_1.n0704 ;
  wire [15:0] \xm8051_golden_model_1.n0710 ;
  wire [15:0] \xm8051_golden_model_1.n0711 ;
  wire [127:0] \xm8051_golden_model_1.n0716 ;
  wire [111:0] \xm8051_golden_model_1.n0717 ;
  wire [127:0] \xm8051_golden_model_1.n0718 ;
  wire [103:0] \xm8051_golden_model_1.n0719 ;
  wire [15:0] \xm8051_golden_model_1.n0720 ;
  wire [127:0] \xm8051_golden_model_1.n0721 ;
  wire [95:0] \xm8051_golden_model_1.n0722 ;
  wire [23:0] \xm8051_golden_model_1.n0723 ;
  wire [127:0] \xm8051_golden_model_1.n0724 ;
  wire [87:0] \xm8051_golden_model_1.n0725 ;
  wire [31:0] \xm8051_golden_model_1.n0726 ;
  wire [127:0] \xm8051_golden_model_1.n0727 ;
  wire [79:0] \xm8051_golden_model_1.n0728 ;
  wire [39:0] \xm8051_golden_model_1.n0729 ;
  wire [127:0] \xm8051_golden_model_1.n0730 ;
  wire [71:0] \xm8051_golden_model_1.n0731 ;
  wire [47:0] \xm8051_golden_model_1.n0732 ;
  wire [127:0] \xm8051_golden_model_1.n0733 ;
  wire [63:0] \xm8051_golden_model_1.n0734 ;
  wire [55:0] \xm8051_golden_model_1.n0735 ;
  wire [127:0] \xm8051_golden_model_1.n0736 ;
  wire [55:0] \xm8051_golden_model_1.n0737 ;
  wire [63:0] \xm8051_golden_model_1.n0738 ;
  wire [127:0] \xm8051_golden_model_1.n0739 ;
  wire [47:0] \xm8051_golden_model_1.n0740 ;
  wire [71:0] \xm8051_golden_model_1.n0741 ;
  wire [127:0] \xm8051_golden_model_1.n0742 ;
  wire [39:0] \xm8051_golden_model_1.n0743 ;
  wire [79:0] \xm8051_golden_model_1.n0744 ;
  wire [127:0] \xm8051_golden_model_1.n0745 ;
  wire [31:0] \xm8051_golden_model_1.n0746 ;
  wire [87:0] \xm8051_golden_model_1.n0747 ;
  wire [127:0] \xm8051_golden_model_1.n0748 ;
  wire [23:0] \xm8051_golden_model_1.n0749 ;
  wire [95:0] \xm8051_golden_model_1.n0750 ;
  wire [127:0] \xm8051_golden_model_1.n0751 ;
  wire [15:0] \xm8051_golden_model_1.n0752 ;
  wire [103:0] \xm8051_golden_model_1.n0753 ;
  wire [127:0] \xm8051_golden_model_1.n0754 ;
  wire [111:0] \xm8051_golden_model_1.n0755 ;
  wire [127:0] \xm8051_golden_model_1.n0756 ;
  wire [119:0] \xm8051_golden_model_1.n0757 ;
  wire [127:0] \xm8051_golden_model_1.n0758 ;
  wire [127:0] \xm8051_golden_model_1.n0759 ;
  wire [127:0] \xm8051_golden_model_1.n0760 ;
  wire [127:0] \xm8051_golden_model_1.n0761 ;
  wire [127:0] \xm8051_golden_model_1.n0762 ;
  wire [127:0] \xm8051_golden_model_1.n0763 ;
  wire [127:0] \xm8051_golden_model_1.n0764 ;
  wire [127:0] \xm8051_golden_model_1.n0765 ;
  wire [127:0] \xm8051_golden_model_1.n0766 ;
  wire [127:0] \xm8051_golden_model_1.n0767 ;
  wire [127:0] \xm8051_golden_model_1.n0768 ;
  wire [127:0] \xm8051_golden_model_1.n0769 ;
  wire [127:0] \xm8051_golden_model_1.n0770 ;
  wire [127:0] \xm8051_golden_model_1.n0771 ;
  wire [127:0] \xm8051_golden_model_1.n0772 ;
  wire \xm8051_golden_model_1.n0775 ;
  wire [15:0] \xm8051_golden_model_1.n0782 ;
  wire [15:0] \xm8051_golden_model_1.n0783 ;
  wire [127:0] \xm8051_golden_model_1.n0788 ;
  wire [111:0] \xm8051_golden_model_1.n0789 ;
  wire [127:0] \xm8051_golden_model_1.n0790 ;
  wire [103:0] \xm8051_golden_model_1.n0791 ;
  wire [15:0] \xm8051_golden_model_1.n0792 ;
  wire [127:0] \xm8051_golden_model_1.n0793 ;
  wire [95:0] \xm8051_golden_model_1.n0794 ;
  wire [23:0] \xm8051_golden_model_1.n0795 ;
  wire [127:0] \xm8051_golden_model_1.n0796 ;
  wire [87:0] \xm8051_golden_model_1.n0797 ;
  wire [31:0] \xm8051_golden_model_1.n0798 ;
  wire [127:0] \xm8051_golden_model_1.n0799 ;
  wire [79:0] \xm8051_golden_model_1.n0800 ;
  wire [39:0] \xm8051_golden_model_1.n0801 ;
  wire [127:0] \xm8051_golden_model_1.n0802 ;
  wire [71:0] \xm8051_golden_model_1.n0803 ;
  wire [47:0] \xm8051_golden_model_1.n0804 ;
  wire [127:0] \xm8051_golden_model_1.n0805 ;
  wire [63:0] \xm8051_golden_model_1.n0806 ;
  wire [55:0] \xm8051_golden_model_1.n0807 ;
  wire [127:0] \xm8051_golden_model_1.n0808 ;
  wire [55:0] \xm8051_golden_model_1.n0809 ;
  wire [63:0] \xm8051_golden_model_1.n0810 ;
  wire [127:0] \xm8051_golden_model_1.n0811 ;
  wire [47:0] \xm8051_golden_model_1.n0812 ;
  wire [71:0] \xm8051_golden_model_1.n0813 ;
  wire [127:0] \xm8051_golden_model_1.n0814 ;
  wire [39:0] \xm8051_golden_model_1.n0815 ;
  wire [79:0] \xm8051_golden_model_1.n0816 ;
  wire [127:0] \xm8051_golden_model_1.n0817 ;
  wire [31:0] \xm8051_golden_model_1.n0818 ;
  wire [87:0] \xm8051_golden_model_1.n0819 ;
  wire [127:0] \xm8051_golden_model_1.n0820 ;
  wire [23:0] \xm8051_golden_model_1.n0821 ;
  wire [95:0] \xm8051_golden_model_1.n0822 ;
  wire [127:0] \xm8051_golden_model_1.n0823 ;
  wire [15:0] \xm8051_golden_model_1.n0824 ;
  wire [103:0] \xm8051_golden_model_1.n0825 ;
  wire [127:0] \xm8051_golden_model_1.n0826 ;
  wire [111:0] \xm8051_golden_model_1.n0827 ;
  wire [127:0] \xm8051_golden_model_1.n0828 ;
  wire [119:0] \xm8051_golden_model_1.n0829 ;
  wire [127:0] \xm8051_golden_model_1.n0830 ;
  wire [127:0] \xm8051_golden_model_1.n0831 ;
  wire [127:0] \xm8051_golden_model_1.n0832 ;
  wire [127:0] \xm8051_golden_model_1.n0833 ;
  wire [127:0] \xm8051_golden_model_1.n0834 ;
  wire [127:0] \xm8051_golden_model_1.n0835 ;
  wire [127:0] \xm8051_golden_model_1.n0836 ;
  wire [127:0] \xm8051_golden_model_1.n0837 ;
  wire [127:0] \xm8051_golden_model_1.n0838 ;
  wire [127:0] \xm8051_golden_model_1.n0839 ;
  wire [127:0] \xm8051_golden_model_1.n0840 ;
  wire [127:0] \xm8051_golden_model_1.n0841 ;
  wire [127:0] \xm8051_golden_model_1.n0842 ;
  wire [127:0] \xm8051_golden_model_1.n0843 ;
  wire [127:0] \xm8051_golden_model_1.n0844 ;
  wire [127:0] \xm8051_golden_model_1.n0849 ;
  wire [111:0] \xm8051_golden_model_1.n0850 ;
  wire [127:0] \xm8051_golden_model_1.n0851 ;
  wire [103:0] \xm8051_golden_model_1.n0852 ;
  wire [15:0] \xm8051_golden_model_1.n0853 ;
  wire [127:0] \xm8051_golden_model_1.n0854 ;
  wire [95:0] \xm8051_golden_model_1.n0855 ;
  wire [23:0] \xm8051_golden_model_1.n0856 ;
  wire [127:0] \xm8051_golden_model_1.n0857 ;
  wire [87:0] \xm8051_golden_model_1.n0858 ;
  wire [31:0] \xm8051_golden_model_1.n0859 ;
  wire [127:0] \xm8051_golden_model_1.n0860 ;
  wire [79:0] \xm8051_golden_model_1.n0861 ;
  wire [39:0] \xm8051_golden_model_1.n0862 ;
  wire [127:0] \xm8051_golden_model_1.n0863 ;
  wire [71:0] \xm8051_golden_model_1.n0864 ;
  wire [47:0] \xm8051_golden_model_1.n0865 ;
  wire [127:0] \xm8051_golden_model_1.n0866 ;
  wire [63:0] \xm8051_golden_model_1.n0867 ;
  wire [55:0] \xm8051_golden_model_1.n0868 ;
  wire [127:0] \xm8051_golden_model_1.n0869 ;
  wire [55:0] \xm8051_golden_model_1.n0870 ;
  wire [63:0] \xm8051_golden_model_1.n0871 ;
  wire [127:0] \xm8051_golden_model_1.n0872 ;
  wire [47:0] \xm8051_golden_model_1.n0873 ;
  wire [71:0] \xm8051_golden_model_1.n0874 ;
  wire [127:0] \xm8051_golden_model_1.n0875 ;
  wire [39:0] \xm8051_golden_model_1.n0876 ;
  wire [79:0] \xm8051_golden_model_1.n0877 ;
  wire [127:0] \xm8051_golden_model_1.n0878 ;
  wire [31:0] \xm8051_golden_model_1.n0879 ;
  wire [87:0] \xm8051_golden_model_1.n0880 ;
  wire [127:0] \xm8051_golden_model_1.n0881 ;
  wire [127:0] \xm8051_golden_model_1.n0884 ;
  wire [15:0] \xm8051_golden_model_1.n0885 ;
  wire [103:0] \xm8051_golden_model_1.n0886 ;
  wire [127:0] \xm8051_golden_model_1.n0887 ;
  wire [111:0] \xm8051_golden_model_1.n0888 ;
  wire [127:0] \xm8051_golden_model_1.n0889 ;
  wire [119:0] \xm8051_golden_model_1.n0890 ;
  wire [127:0] \xm8051_golden_model_1.n0891 ;
  wire [127:0] \xm8051_golden_model_1.n0892 ;
  wire [127:0] \xm8051_golden_model_1.n0893 ;
  wire [127:0] \xm8051_golden_model_1.n0894 ;
  wire [127:0] \xm8051_golden_model_1.n0895 ;
  wire [127:0] \xm8051_golden_model_1.n0896 ;
  wire [127:0] \xm8051_golden_model_1.n0897 ;
  wire [127:0] \xm8051_golden_model_1.n0898 ;
  wire [127:0] \xm8051_golden_model_1.n0899 ;
  wire [127:0] \xm8051_golden_model_1.n0900 ;
  wire [127:0] \xm8051_golden_model_1.n0901 ;
  wire [127:0] \xm8051_golden_model_1.n0902 ;
  wire [127:0] \xm8051_golden_model_1.n0903 ;
  wire [127:0] \xm8051_golden_model_1.n0904 ;
  wire [127:0] \xm8051_golden_model_1.n0905 ;
  wire [15:0] \xm8051_golden_model_1.n0909 ;
  wire [15:0] \xm8051_golden_model_1.n0910 ;
  wire [15:0] \xm8051_golden_model_1.n0920 ;
  wire [15:0] \xm8051_golden_model_1.n0921 ;
  wire [159:0] \xm8051_golden_model_1.n0931 ;
  wire [127:0] \xm8051_golden_model_1.n0956 ;
  wire [159:0] \xm8051_golden_model_1.n0958 ;
  wire [127:0] \xm8051_golden_model_1.n0966 ;
  wire [159:0] \xm8051_golden_model_1.n0968 ;
  wire [15:0] \xm8051_golden_model_1.n0972 ;
  wire [15:0] \xm8051_golden_model_1.n0973 ;
  wire [159:0] \xm8051_golden_model_1.n0983 ;
  wire [159:0] \xm8051_golden_model_1.n1236 ;
  wire [511:0] \xm8051_golden_model_1.n1240 ;
  wire [159:0] \xm8051_golden_model_1.n1244 ;
  wire [511:0] \xm8051_golden_model_1.n1248 ;
  wire [159:0] \xm8051_golden_model_1.n1250 ;
  wire [127:0] \xm8051_golden_model_1.n1254 ;
  wire [159:0] \xm8051_golden_model_1.n1256 ;
  wire [15:0] \xm8051_golden_model_1.n1262 ;
  wire [15:0] \xm8051_golden_model_1.n1263 ;
  wire [159:0] \xm8051_golden_model_1.n1267 ;
  wire [159:0] \xm8051_golden_model_1.n1271 ;
  wire [159:0] \xm8051_golden_model_1.n1275 ;
  wire [127:0] \xm8051_golden_model_1.n1279 ;
  wire [159:0] \xm8051_golden_model_1.n1281 ;
  wire [159:0] \xm8051_golden_model_1.n1285 ;
  wire [127:0] \xm8051_golden_model_1.n1290 ;
  wire [159:0] \xm8051_golden_model_1.n1295 ;
  wire [159:0] \xm8051_golden_model_1.n1299 ;
  wire [127:0] \xm8051_golden_model_1.n1303 ;
  wire [159:0] \xm8051_golden_model_1.n1305 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_0 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_1 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_10 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_100 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_101 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_102 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_103 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_104 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_105 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_106 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_107 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_108 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_109 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_11 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_110 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_111 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_112 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_113 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_114 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_115 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_116 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_117 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_118 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_119 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_12 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_13 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_14 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_15 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_16 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_17 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_18 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_19 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_2 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_20 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_21 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_22 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_23 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_24 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_25 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_26 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_27 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_28 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_29 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_3 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_30 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_31 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_32 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_33 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_34 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_35 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_36 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_37 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_38 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_39 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_4 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_40 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_41 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_42 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_43 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_44 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_45 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_46 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_47 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_48 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_49 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_5 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_50 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_51 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_52 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_53 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_54 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_55 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_56 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_57 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_58 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_59 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_6 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_60 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_61 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_62 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_63 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_64 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_65 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_66 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_67 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_68 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_69 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_7 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_70 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_71 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_72 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_73 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_74 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_75 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_76 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_77 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_78 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_79 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_8 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_80 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_81 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_82 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_83 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_84 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_85 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_86 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_87 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_88 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_89 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_9 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_90 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_91 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_92 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_93 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_94 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_95 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_96 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_97 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_98 ;
  wire \xm8051_golden_model_1.nondet_memwrite_choice_99 ;
  wire \xm8051_golden_model_1.rst ;
  wire [15:0] \xm8051_golden_model_1.sha_bytes_processed ;
  wire [15:0] \xm8051_golden_model_1.sha_bytes_processed_08 ;
  wire [15:0] \xm8051_golden_model_1.sha_bytes_processed_09 ;
  wire [15:0] \xm8051_golden_model_1.sha_bytes_processed_0a ;
  wire [15:0] \xm8051_golden_model_1.sha_bytes_processed_0b ;
  wire [15:0] \xm8051_golden_model_1.sha_len ;
  wire [7:0] \xm8051_golden_model_1.sha_state ;
  not (_1270_, proc_stb);
  not (_1271_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [0]);
  nor (_1272_, proc_addr[6], proc_addr[7]);
  not (_1273_, _1272_);
  and (_1274_, proc_addr[12], proc_addr[14]);
  and (_1275_, proc_addr[15], proc_addr[13]);
  and (_1276_, _1275_, _1274_);
  and (_1277_, proc_addr[11], proc_addr[10]);
  and (_1278_, proc_addr[9], proc_addr[8]);
  and (_1279_, _1278_, _1277_);
  nand (_1280_, _1279_, _1276_);
  or (_1281_, _1280_, _1273_);
  and (_1282_, _1281_, proc_stb);
  nor (_1283_, proc_addr[5], proc_addr[4]);
  and (_1284_, _1283_, _1272_);
  not (_1285_, proc_addr[8]);
  and (_1286_, proc_addr[9], _1285_);
  and (_1287_, _1286_, _1277_);
  and (_1288_, _1287_, _1276_);
  nand (_1289_, _1288_, _1284_);
  nand (_1290_, _1289_, _1282_);
  and (_1291_, _1290_, _1271_);
  and (_1292_, _1291_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0]);
  or (_1293_, _1292_, \oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbiter_state );
  not (_1294_, \oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbiter_state );
  nor (_1295_, \oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbit_holder [1], _1294_);
  not (_1296_, _1295_);
  and (_1297_, _1296_, _1293_);
  not (_1298_, _1297_);
  nor (_1299_, \oc8051_xiommu_impl_1.oc8051_xram_i.ackr , \oc8051_xiommu_impl_1.oc8051_xram_i.ackw );
  not (_1300_, _1299_);
  and (_1301_, \oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbiter_state , \oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbit_holder [0]);
  and (_1302_, _1290_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [0]);
  and (_1303_, _1302_, _1294_);
  nor (_1304_, _1303_, _1301_);
  and (_1305_, _1304_, _1300_);
  and (_1306_, _1305_, _1298_);
  nor (_1307_, _1281_, _1270_);
  and (_1308_, _1284_, _1287_);
  and (_1309_, _1308_, _1276_);
  and (_1310_, _1309_, proc_stb);
  or (_1311_, _1310_, _1307_);
  nor (_1312_, _1311_, _1306_);
  nor (_1313_, _1312_, _1270_);
  and (_1314_, _1313_, proc_wr);
  or (_1315_, \xm8051_golden_model_1.sha_state [6], \xm8051_golden_model_1.sha_state [7]);
  or (_1316_, \xm8051_golden_model_1.sha_state [2], \xm8051_golden_model_1.sha_state [4]);
  or (_1317_, _1316_, _1315_);
  nor (_1318_, \xm8051_golden_model_1.sha_state [1], \xm8051_golden_model_1.sha_state [0]);
  not (_1319_, _1318_);
  or (_1320_, \xm8051_golden_model_1.sha_state [5], \xm8051_golden_model_1.sha_state [3]);
  or (_1321_, _1320_, _1319_);
  nor (_1322_, _1321_, _1317_);
  nor (_1323_, proc_addr[1], proc_addr[2]);
  nor (_1324_, proc_addr[3], proc_addr[0]);
  and (_1325_, _1324_, _1323_);
  and (_1326_, _1325_, proc_data_in[0]);
  and (_1327_, _1326_, _1309_);
  and (_1328_, _1327_, _1322_);
  nand (_1329_, _1328_, _1314_);
  not (_1330_, rst);
  and (_1331_, \xm8051_golden_model_1.sha_bytes_processed [1], _1330_);
  and (_1895_[1], _1331_, _1329_);
  not (_1332_, proc_addr[0]);
  nor (_1333_, \xm8051_golden_model_1.aes_state [2], \xm8051_golden_model_1.aes_state [3]);
  nor (_1334_, \xm8051_golden_model_1.aes_state [7], \xm8051_golden_model_1.aes_state [6]);
  and (_1335_, _1334_, _1333_);
  nor (_1336_, \xm8051_golden_model_1.aes_state [1], \xm8051_golden_model_1.aes_state [0]);
  nor (_1337_, \xm8051_golden_model_1.aes_state [5], \xm8051_golden_model_1.aes_state [4]);
  and (_1338_, _1337_, _1336_);
  and (_1339_, _1338_, _1335_);
  and (_1340_, _1339_, _1314_);
  not (_1341_, proc_addr[1]);
  not (_1342_, proc_addr[3]);
  and (_1343_, _1342_, proc_addr[2]);
  and (_1344_, _1343_, _1341_);
  not (_1345_, _1280_);
  and (_1346_, _1284_, _1345_);
  and (_1347_, _1346_, _1344_);
  and (_1348_, _1347_, _1340_);
  and (_1349_, _1348_, _1332_);
  and (_1350_, _1349_, proc_data_in[4]);
  not (_1351_, \xm8051_golden_model_1.aes_len [4]);
  nor (_1352_, _1349_, _1351_);
  or (_1353_, _1352_, _1350_);
  and (_1893_[4], _1353_, _1330_);
  not (_1354_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [13]);
  nor (_1355_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [1], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [0]);
  and (_1356_, _1355_, proc_wr);
  and (_1357_, _1356_, _1307_);
  and (_1358_, _1357_, _1347_);
  and (_1359_, _1358_, proc_addr[0]);
  nor (_1360_, _1359_, _1354_);
  and (_1361_, _1359_, proc_data_in[5]);
  or (_1362_, _1361_, _1360_);
  and (_0508_, _1362_, _1330_);
  and (_1363_, _1348_, proc_addr[0]);
  and (_1364_, _1363_, proc_data_in[4]);
  not (_1365_, \xm8051_golden_model_1.aes_len [12]);
  nor (_1366_, _1363_, _1365_);
  or (_1367_, _1366_, _1364_);
  and (_1893_[12], _1367_, _1330_);
  not (_1368_, \xm8051_golden_model_1.sha_bytes_processed [8]);
  not (_1369_, \xm8051_golden_model_1.sha_state [0]);
  and (_1370_, \xm8051_golden_model_1.sha_state [1], _1369_);
  nor (_1371_, _1370_, _1368_);
  not (_1372_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0]);
  and (_1373_, _1372_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [1]);
  and (_1374_, _1373_, ABINPUT000[161]);
  nor (_1375_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [1]);
  and (_1376_, _1375_, proc_wr);
  and (_1377_, _1376_, _1310_);
  and (_1378_, _1377_, _1327_);
  nor (_1379_, _1378_, _1374_);
  not (_1380_, _1379_);
  not (_1381_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [1]);
  and (_1382_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0], _1381_);
  and (_1383_, _1305_, _1297_);
  and (_1384_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [0], \oc8051_xiommu_impl_1.sha_top_i.byte_counter [1]);
  and (_1385_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [3], \oc8051_xiommu_impl_1.sha_top_i.byte_counter [2]);
  and (_1386_, _1385_, _1384_);
  and (_1387_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [4], \oc8051_xiommu_impl_1.sha_top_i.byte_counter [5]);
  and (_1388_, _1387_, _1386_);
  not (_1389_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [0]);
  and (_1390_, _1383_, _1382_);
  or (_1391_, _1390_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [0]);
  and (_1392_, _1390_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [0]);
  nor (_1393_, _1375_, _1392_);
  and (_1394_, _1393_, _1391_);
  or (_1395_, _1394_, _1389_);
  nand (_1396_, _1394_, _1389_);
  and (_1397_, _1396_, _1395_);
  not (_1398_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [1]);
  or (_1399_, _1392_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [1]);
  and (_1400_, _1392_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [1]);
  nor (_1401_, _1375_, _1400_);
  and (_1402_, _1401_, _1399_);
  or (_1403_, _1402_, _1398_);
  and (_1404_, _1403_, _1397_);
  nand (_1405_, _1402_, _1398_);
  and (_1406_, _1405_, _1404_);
  not (_1407_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [3]);
  not (_1408_, _1375_);
  and (_1409_, _1400_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [2]);
  nand (_1410_, _1409_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [3]);
  or (_1411_, _1409_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [3]);
  and (_1412_, _1411_, _1410_);
  and (_1413_, _1412_, _1408_);
  or (_1414_, _1413_, _1407_);
  nand (_1415_, _1413_, _1407_);
  and (_1416_, _1415_, _1414_);
  not (_1417_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [2]);
  or (_1418_, _1400_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [2]);
  nor (_1419_, _1375_, _1409_);
  and (_1420_, _1419_, _1418_);
  or (_1421_, _1420_, _1417_);
  nand (_1422_, _1420_, _1417_);
  and (_1423_, _1422_, _1421_);
  and (_1424_, _1423_, _1416_);
  and (_1425_, _1424_, _1406_);
  not (_1426_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [4]);
  not (_1427_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [4]);
  or (_1428_, _1410_, _1427_);
  nand (_1429_, _1410_, _1427_);
  and (_1430_, _1429_, _1408_);
  and (_1431_, _1430_, _1428_);
  or (_1432_, _1431_, _1426_);
  nand (_1433_, _1431_, _1426_);
  and (_1434_, _1433_, _1432_);
  not (_1435_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [5]);
  not (_1436_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [5]);
  nand (_1437_, _1428_, _1436_);
  and (_1438_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [2], \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [3]);
  and (_1439_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [4], \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [5]);
  and (_1440_, _1439_, _1438_);
  and (_1441_, _1440_, _1400_);
  nor (_1442_, _1441_, _1375_);
  and (_1443_, _1442_, _1437_);
  or (_1444_, _1443_, _1435_);
  nand (_1445_, _1443_, _1435_);
  and (_1446_, _1445_, _1444_);
  and (_1447_, _1446_, _1434_);
  not (_1448_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [7]);
  nand (_1449_, _1441_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [6]);
  or (_1450_, _1449_, _1448_);
  nand (_1451_, _1449_, _1448_);
  and (_1452_, _1451_, _1450_);
  and (_1453_, _1452_, _1408_);
  nor (_1454_, _1453_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [7]);
  and (_1455_, _1453_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [7]);
  or (_1456_, _1455_, _1454_);
  not (_1457_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [6]);
  or (_1458_, _1441_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [6]);
  and (_1459_, _1449_, _1408_);
  and (_1460_, _1459_, _1458_);
  nand (_1461_, _1460_, _1457_);
  or (_1462_, _1460_, _1457_);
  and (_1463_, _1462_, _1461_);
  and (_1464_, _1463_, _1456_);
  and (_1465_, _1464_, _1447_);
  and (_1466_, _1465_, _1425_);
  not (_1467_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [9]);
  not (_1468_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [9]);
  and (_1469_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [1], \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [0]);
  and (_1470_, _1438_, _1469_);
  and (_1471_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [6], \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [7]);
  and (_1472_, _1471_, _1439_);
  and (_1473_, _1472_, _1470_);
  and (_1474_, _1473_, _1390_);
  nand (_1475_, _1474_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [8]);
  or (_1476_, _1475_, _1468_);
  nand (_1477_, _1475_, _1468_);
  and (_1478_, _1477_, _1476_);
  and (_1479_, _1478_, _1408_);
  nand (_1480_, _1479_, _1467_);
  or (_1481_, _1479_, _1467_);
  and (_1482_, _1481_, _1480_);
  not (_1483_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [8]);
  or (_1484_, _1474_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [8]);
  and (_1485_, _1475_, _1408_);
  and (_1486_, _1485_, _1484_);
  nand (_1487_, _1486_, _1483_);
  or (_1488_, _1486_, _1483_);
  and (_1489_, _1488_, _1487_);
  and (_1490_, _1489_, _1482_);
  not (_1491_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [11]);
  not (_1492_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [11]);
  not (_1493_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [10]);
  or (_1494_, _1476_, _1493_);
  or (_1495_, _1494_, _1492_);
  nand (_1496_, _1494_, _1492_);
  and (_1498_, _1496_, _1408_);
  and (_1499_, _1498_, _1495_);
  nand (_1501_, _1499_, _1491_);
  or (_1502_, _1499_, _1491_);
  and (_1503_, _1502_, _1501_);
  not (_1504_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [10]);
  nand (_1505_, _1476_, _1493_);
  and (_1506_, _1505_, _1408_);
  and (_1507_, _1506_, _1494_);
  or (_1508_, _1507_, _1504_);
  nand (_1509_, _1507_, _1504_);
  and (_1510_, _1509_, _1508_);
  and (_1511_, _1510_, _1503_);
  and (_1512_, _1511_, _1490_);
  not (_1513_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [13]);
  not (_1514_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [12]);
  and (_1515_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [8], \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [9]);
  and (_1516_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [10], \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [11]);
  and (_1517_, _1516_, _1515_);
  nand (_1518_, _1517_, _1474_);
  or (_1519_, _1518_, _1514_);
  nand (_1520_, _1519_, _1513_);
  and (_1521_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [12], \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [13]);
  not (_1522_, _1521_);
  or (_1523_, _1522_, _1518_);
  and (_1524_, _1523_, _1408_);
  and (_1525_, _1524_, _1520_);
  nor (_1526_, _1525_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [13]);
  and (_1527_, _1525_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [13]);
  or (_1528_, _1527_, _1526_);
  not (_1529_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [12]);
  nand (_1530_, _1518_, _1514_);
  and (_1531_, _1519_, _1408_);
  and (_1532_, _1531_, _1530_);
  or (_1533_, _1532_, _1529_);
  nand (_1534_, _1532_, _1529_);
  and (_1535_, _1534_, _1533_);
  and (_1536_, _1535_, _1528_);
  not (_1537_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [15]);
  not (_1538_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [14]);
  or (_1539_, _1523_, _1538_);
  and (_1540_, _1539_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [15]);
  nor (_1541_, _1539_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [15]);
  or (_1542_, _1541_, _1540_);
  and (_1543_, _1542_, _1408_);
  nand (_1544_, _1543_, _1537_);
  or (_1545_, _1543_, _1537_);
  and (_1546_, _1545_, _1544_);
  not (_1547_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [14]);
  and (_1548_, _1523_, _1538_);
  nor (_1549_, _1548_, _1375_);
  and (_1550_, _1549_, _1539_);
  or (_1552_, _1550_, _1547_);
  nand (_1553_, _1550_, _1547_);
  and (_1555_, _1553_, _1552_);
  and (_1556_, _1555_, _1546_);
  and (_1557_, _1556_, _1536_);
  and (_1558_, _1557_, _1512_);
  and (_1559_, _1558_, _1466_);
  or (_1560_, _1559_, _1388_);
  nand (_1561_, _1560_, _1383_);
  nand (_1562_, _1561_, _1382_);
  not (_1563_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [2]);
  and (_1564_, _1384_, _1383_);
  and (_1565_, _1564_, _1563_);
  nor (_1566_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [3], \oc8051_xiommu_impl_1.sha_top_i.byte_counter [5]);
  and (_1567_, _1566_, _1565_);
  and (_1568_, _1567_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [4]);
  and (_1569_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [1]);
  not (_1570_, _1569_);
  nor (_1571_, _1570_, _1568_);
  nor (_1572_, _1571_, _1380_);
  nand (_1573_, _1572_, _1562_);
  nor (_1574_, _1573_, _1372_);
  or (_1575_, _1574_, _1380_);
  and (_1576_, \xm8051_golden_model_1.sha_bytes_processed [7], \xm8051_golden_model_1.sha_bytes_processed [6]);
  nand (_1577_, _1576_, _1575_);
  nor (_1578_, _1577_, _1368_);
  and (_1579_, _1577_, _1368_);
  nor (_1580_, _1579_, _1578_);
  and (_1581_, _1580_, _1370_);
  or (_1582_, _1581_, _1371_);
  and (_1583_, _1582_, _1319_);
  and (_1584_, _1318_, \xm8051_golden_model_1.sha_bytes_processed [8]);
  and (_1585_, _1584_, _1329_);
  or (_1586_, _1585_, _1583_);
  and (_1895_[8], _1586_, _1330_);
  and (_1587_, \xm8051_golden_model_1.sha_bytes_processed [0], _1330_);
  and (_1895_[0], _1587_, _1329_);
  not (_1589_, _1326_);
  or (_1590_, _1589_, _1289_);
  or (_1591_, _1320_, _1317_);
  or (_1592_, _1591_, _1590_);
  nor (_1593_, _1592_, _1319_);
  nand (_1594_, _1593_, _1314_);
  and (_1595_, \xm8051_golden_model_1.aes_state [1], \xm8051_golden_model_1.aes_state [0]);
  and (_1596_, _1595_, _1318_);
  not (_1597_, _1596_);
  or (_1598_, _1597_, _1594_);
  and (_1599_, _1598_, \xm8051_golden_model_1.sha_bytes_processed [14]);
  not (_1600_, _1370_);
  not (_1601_, \xm8051_golden_model_1.sha_bytes_processed [13]);
  not (_1602_, \xm8051_golden_model_1.sha_bytes_processed [12]);
  and (_1603_, \xm8051_golden_model_1.sha_bytes_processed [8], \xm8051_golden_model_1.sha_bytes_processed [9]);
  and (_1604_, _1603_, _1576_);
  and (_1605_, _1604_, _1575_);
  and (_1606_, _1605_, \xm8051_golden_model_1.sha_bytes_processed [10]);
  nand (_1607_, _1606_, \xm8051_golden_model_1.sha_bytes_processed [11]);
  or (_1608_, _1607_, _1602_);
  or (_1609_, _1608_, _1601_);
  nor (_1610_, _1609_, _1600_);
  or (_1611_, _1610_, _1599_);
  not (_1612_, \xm8051_golden_model_1.sha_bytes_processed [14]);
  or (_1613_, _1609_, _1612_);
  or (_1614_, _1613_, _1600_);
  and (_1615_, _1614_, _1611_);
  not (_1616_, _1595_);
  and (_1617_, _1616_, _1318_);
  or (_1618_, _1617_, _1615_);
  nand (_1619_, _1329_, \xm8051_golden_model_1.sha_bytes_processed [14]);
  nand (_1620_, _1617_, _1619_);
  and (_1621_, _1620_, _1330_);
  and (_1895_[14], _1621_, _1618_);
  or (_1622_, _1304_, _1297_);
  nand (_1623_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [1], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [0]);
  nor (_1624_, _1623_, _1622_);
  not (_1625_, _1624_);
  nor (_1626_, _1301_, _1290_);
  and (_1627_, _1626_, _1298_);
  and (_1628_, _1627_, proc_wr);
  and (_1629_, _1297_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0]);
  and (_1630_, _1629_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [1]);
  nor (_1631_, _1630_, _1628_);
  and (_1632_, _1631_, _1625_);
  not (_1633_, _1632_);
  not (_1634_, \oc8051_xiommu_impl_1.oc8051_xram_i.cnt [2]);
  nor (_1635_, \oc8051_xiommu_impl_1.oc8051_xram_i.cnt [0], \oc8051_xiommu_impl_1.oc8051_xram_i.cnt [1]);
  and (_1636_, _1635_, _1634_);
  and (_1637_, _1636_, _1330_);
  and (_1497_, _1637_, _1633_);
  not (_1638_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [1]);
  and (_1639_, _1358_, _1332_);
  nor (_1640_, _1639_, _1638_);
  and (_1641_, _1639_, proc_data_in[1]);
  or (_1642_, _1641_, _1640_);
  and (_1500_, _1642_, _1330_);
  or (_1643_, _1622_, _1299_);
  not (_1644_, \oc8051_xiommu_impl_1.aes_top_i.byte_counter [3]);
  and (_1645_, \oc8051_xiommu_impl_1.aes_top_i.byte_counter [1], \oc8051_xiommu_impl_1.aes_top_i.byte_counter [0]);
  nand (_1646_, _1645_, \oc8051_xiommu_impl_1.aes_top_i.byte_counter [2]);
  nor (_1647_, _1646_, _1644_);
  not (_1648_, _1647_);
  or (_1649_, _1648_, _1643_);
  or (_1650_, _1649_, _1623_);
  and (_1651_, _1650_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [10]);
  not (_1652_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [10]);
  and (_1653_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [4], \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [5]);
  and (_1654_, _1653_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [6]);
  and (_1655_, _1654_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [7]);
  and (_1657_, _1655_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [8]);
  and (_1658_, _1657_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [9]);
  and (_1659_, _1658_, _1652_);
  nor (_1660_, _1658_, _1652_);
  nor (_1661_, _1660_, _1659_);
  nor (_1662_, _1661_, _1650_);
  or (_1663_, _1662_, _1651_);
  and (_1664_, _1346_, _1326_);
  and (_1665_, _1664_, _1357_);
  nor (_1666_, _1665_, rst);
  and (_1551_, _1666_, _1663_);
  and (_1668_, _1650_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [14]);
  nor (_1669_, _1649_, _1623_);
  not (_1670_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [14]);
  and (_1671_, _1658_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [10]);
  and (_1672_, _1671_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [11]);
  and (_1673_, _1672_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [12]);
  and (_1674_, _1673_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [13]);
  nand (_1675_, _1674_, _1670_);
  or (_1676_, _1674_, _1670_);
  nand (_1677_, _1676_, _1675_);
  and (_1678_, _1677_, _1669_);
  or (_1679_, _1678_, _1668_);
  and (_1554_, _1679_, _1666_);
  not (_1680_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [2]);
  nor (_1681_, _1639_, _1680_);
  and (_1682_, _1639_, proc_data_in[2]);
  or (_1683_, _1682_, _1681_);
  and (_1588_, _1683_, _1330_);
  not (_1685_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [3]);
  nor (_1686_, _1639_, _1685_);
  and (_1687_, _1639_, proc_data_in[3]);
  or (_1688_, _1687_, _1686_);
  and (_1656_, _1688_, _1330_);
  not (_1689_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [15]);
  nor (_1690_, _1359_, _1689_);
  and (_1691_, _1359_, proc_data_in[7]);
  or (_1692_, _1691_, _1690_);
  and (_1667_, _1692_, _1330_);
  and (_1684_, _1394_, _1330_);
  nor (_1693_, _1622_, _1271_);
  not (_1694_, _1693_);
  nor (_1695_, _1629_, _1627_);
  and (_1696_, _1695_, _1694_);
  not (_1697_, _1696_);
  and (_1698_, _1697_, _1632_);
  and (_1703_, _1698_, _1637_);
  nor (_1699_, _1646_, _1643_);
  not (_1700_, _1643_);
  and (_1701_, _1645_, _1700_);
  or (_1702_, _1701_, \oc8051_xiommu_impl_1.aes_top_i.byte_counter [2]);
  nand (_1704_, _1702_, _1666_);
  nor (_1709_, _1704_, _1699_);
  nor (_1705_, _1574_, _1380_);
  and (_1706_, \xm8051_golden_model_1.sha_bytes_processed [11], \xm8051_golden_model_1.sha_bytes_processed [10]);
  and (_1707_, _1706_, _1603_);
  and (_1708_, _1707_, _1576_);
  and (_1710_, _1708_, \xm8051_golden_model_1.sha_bytes_processed [12]);
  and (_1711_, _1710_, _1601_);
  nor (_1712_, _1710_, _1601_);
  nor (_1713_, _1712_, _1711_);
  nor (_1714_, _1713_, _1705_);
  and (_1715_, _1705_, \xm8051_golden_model_1.sha_bytes_processed [13]);
  or (_1716_, _1715_, _1714_);
  and (_1717_, _1716_, _1370_);
  and (_1718_, _1318_, \xm8051_golden_model_1.sha_bytes_processed [13]);
  and (_1719_, _1718_, _1329_);
  and (_1720_, \xm8051_golden_model_1.sha_state [0], \xm8051_golden_model_1.sha_bytes_processed [13]);
  or (_1721_, _1720_, _1719_);
  or (_1722_, _1721_, _1717_);
  and (_1895_[13], _1722_, _1330_);
  and (_1723_, \xm8051_golden_model_1.sha_bytes_processed [5], _1330_);
  and (_1895_[5], _1723_, _1329_);
  not (_1724_, proc_addr[7]);
  and (_1725_, proc_addr[6], _1724_);
  and (_1726_, _1725_, _1283_);
  nand (_1727_, _1726_, _1325_);
  and (_1728_, _1727_, _1273_);
  and (_1729_, _1728_, _1345_);
  nor (_1730_, _1727_, _1280_);
  nor (_1731_, _1730_, _1729_);
  and (_1732_, _1731_, _1345_);
  and (_1733_, _1732_, proc_stb);
  and (_1734_, _1733_, proc_wr);
  and (_1735_, _1734_, _1355_);
  and (_1736_, _1325_, _1284_);
  and (_1737_, _1736_, _1345_);
  and (_1738_, _1737_, proc_data_in[0]);
  nand (_1739_, _1738_, _1735_);
  not (_1740_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [5]);
  or (_1741_, _1669_, _1740_);
  and (_1742_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [4], _1740_);
  not (_1743_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [4]);
  and (_1744_, _1743_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [5]);
  nor (_1745_, _1744_, _1742_);
  or (_1746_, _1745_, _1650_);
  nand (_1747_, _1746_, _1741_);
  and (_1748_, _1747_, _1739_);
  and (_1834_, _1748_, _1330_);
  not (_1749_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [7]);
  or (_1750_, _1669_, _1749_);
  and (_1751_, _1654_, _1749_);
  nor (_1752_, _1654_, _1749_);
  nor (_1753_, _1752_, _1751_);
  or (_1754_, _1753_, _1650_);
  nand (_1755_, _1754_, _1750_);
  and (_1756_, _1755_, _1739_);
  and (_1837_, _1756_, _1330_);
  and (_1757_, _1336_, _1318_);
  and (_1758_, _1649_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [0]);
  not (_1759_, _1758_);
  nand (_1760_, _1679_, _1739_);
  nand (_1761_, _1760_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [14]);
  or (_1762_, _1760_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [14]);
  and (_1763_, _1762_, _1761_);
  and (_1764_, _1307_, proc_wr);
  and (_1765_, _1764_, _1355_);
  and (_1766_, _1664_, _1765_);
  not (_1767_, _1766_);
  and (_1768_, _1650_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [15]);
  not (_1769_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [15]);
  and (_1770_, _1674_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [14]);
  nand (_1771_, _1770_, _1769_);
  or (_1772_, _1770_, _1769_);
  nand (_1773_, _1772_, _1771_);
  and (_1774_, _1773_, _1669_);
  or (_1775_, _1774_, _1768_);
  and (_1776_, _1775_, _1767_);
  nand (_1777_, _1776_, _1689_);
  or (_1778_, _1776_, _1689_);
  and (_1779_, _1778_, _1777_);
  and (_1780_, _1779_, _1763_);
  and (_1781_, _1673_, _1669_);
  or (_1782_, _1781_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [13]);
  not (_1783_, _1665_);
  nand (_1784_, _1781_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [13]);
  and (_1785_, _1784_, _1783_);
  and (_1786_, _1785_, _1782_);
  or (_1787_, _1786_, _1354_);
  nand (_1788_, _1786_, _1354_);
  and (_1789_, _1788_, _1787_);
  not (_1790_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [12]);
  not (_1791_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [12]);
  nand (_1792_, _1672_, _1669_);
  nand (_1793_, _1792_, _1791_);
  or (_1794_, _1792_, _1791_);
  and (_1795_, _1794_, _1793_);
  nand (_1796_, _1795_, _1767_);
  nand (_1797_, _1796_, _1790_);
  or (_1798_, _1796_, _1790_);
  nand (_1799_, _1798_, _1797_);
  and (_1800_, _1799_, _1789_);
  and (_1801_, _1800_, _1780_);
  nand (_1802_, _1739_, _1663_);
  and (_1803_, _1802_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [10]);
  nor (_1804_, _1802_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [10]);
  nor (_1805_, _1804_, _1803_);
  not (_1806_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [11]);
  and (_1807_, _1650_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [11]);
  not (_1808_, _1671_);
  nor (_1809_, _1808_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [11]);
  and (_1810_, _1808_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [11]);
  nor (_1811_, _1810_, _1809_);
  nor (_1812_, _1811_, _1650_);
  or (_1813_, _1812_, _1807_);
  and (_1814_, _1813_, _1767_);
  nand (_1815_, _1814_, _1806_);
  or (_1816_, _1814_, _1806_);
  and (_1817_, _1816_, _1815_);
  and (_1818_, _1817_, _1805_);
  and (_1819_, _1650_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [8]);
  not (_1820_, _1655_);
  nor (_1821_, _1820_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [8]);
  and (_1822_, _1820_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [8]);
  nor (_1823_, _1822_, _1821_);
  nor (_1824_, _1823_, _1650_);
  or (_1825_, _1824_, _1819_);
  nand (_1826_, _1825_, _1767_);
  and (_1827_, _1826_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [8]);
  not (_1828_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [9]);
  and (_1829_, _1657_, _1669_);
  or (_1830_, _1829_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [9]);
  and (_1831_, _1658_, _1669_);
  nor (_1832_, _1665_, _1831_);
  and (_1833_, _1832_, _1830_);
  or (_1835_, _1833_, _1828_);
  nand (_1836_, _1833_, _1828_);
  and (_1838_, _1836_, _1835_);
  or (_1839_, _1826_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [8]);
  nand (_1840_, _1839_, _1838_);
  nor (_1841_, _1840_, _1827_);
  and (_1842_, _1841_, _1818_);
  and (_1843_, _1842_, _1801_);
  not (_1844_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [7]);
  or (_1845_, _1756_, _1844_);
  nand (_1846_, _1756_, _1844_);
  and (_1847_, _1846_, _1845_);
  and (_1848_, _1650_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [6]);
  not (_1849_, _1653_);
  nor (_1850_, _1849_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [6]);
  and (_1851_, _1849_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [6]);
  nor (_1852_, _1851_, _1850_);
  nor (_1853_, _1852_, _1650_);
  or (_1854_, _1853_, _1848_);
  nand (_1855_, _1854_, _1767_);
  and (_1856_, _1855_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [6]);
  nor (_1857_, _1855_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [6]);
  nor (_1858_, _1857_, _1856_);
  and (_1859_, _1858_, _1847_);
  not (_1860_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [4]);
  or (_1861_, _1669_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [4]);
  or (_1862_, _1650_, _1743_);
  and (_1863_, _1862_, _1783_);
  and (_1864_, _1863_, _1861_);
  or (_1865_, _1864_, _1860_);
  nand (_1866_, _1864_, _1860_);
  and (_1867_, _1866_, _1865_);
  or (_1868_, _1748_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [5]);
  not (_1869_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [5]);
  nand (_1870_, _1747_, _1739_);
  or (_1871_, _1870_, _1869_);
  nand (_1872_, _1871_, _1868_);
  and (_1873_, _1872_, _1867_);
  and (_1874_, _1873_, _1859_);
  and (_1875_, _1783_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [2]);
  nor (_1876_, _1875_, _1680_);
  not (_1877_, _1876_);
  and (_1878_, _1783_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [3]);
  and (_1879_, _1878_, _1685_);
  nor (_1880_, _1879_, _1877_);
  nor (_1881_, _1878_, _1685_);
  and (_1882_, _1875_, _1680_);
  not (_1883_, _1882_);
  nor (_1884_, _1879_, _1881_);
  and (_1885_, _1884_, _1877_);
  and (_1886_, _1885_, _1883_);
  not (_1887_, _1886_);
  and (_1888_, _1783_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [1]);
  nor (_1889_, _1888_, _1638_);
  and (_1890_, _1888_, _1638_);
  not (_1891_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [0]);
  and (_0002_, _1783_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [0]);
  and (_0003_, _0002_, _1891_);
  or (_0004_, _0003_, _1889_);
  nor (_0005_, _0004_, _1890_);
  nor (_0006_, _0005_, _1889_);
  nor (_0007_, _0006_, _1887_);
  or (_0008_, _0007_, _1881_);
  or (_0009_, _0008_, _1880_);
  nand (_0010_, _0009_, _1874_);
  or (_0011_, _1870_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [5]);
  or (_0012_, _1748_, _1869_);
  nand (_0013_, _1865_, _0012_);
  and (_0014_, _0013_, _0011_);
  nand (_0015_, _0014_, _1859_);
  nand (_0016_, _1856_, _1846_);
  and (_0017_, _0016_, _1845_);
  and (_0018_, _0017_, _0015_);
  nand (_0019_, _0018_, _0010_);
  nand (_0020_, _0019_, _1843_);
  nand (_0021_, _1836_, _1827_);
  nand (_0022_, _0021_, _1835_);
  nand (_0023_, _0022_, _1818_);
  nand (_0024_, _1803_, _1815_);
  and (_0025_, _0024_, _1816_);
  nand (_0026_, _0025_, _0023_);
  nand (_0027_, _0026_, _1801_);
  and (_0028_, _1796_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [12]);
  nand (_0029_, _1788_, _0028_);
  nand (_0030_, _0029_, _1787_);
  nand (_0031_, _0030_, _1780_);
  not (_0032_, _1761_);
  nand (_0033_, _0032_, _1777_);
  and (_0034_, _0033_, _1778_);
  and (_0035_, _0034_, _0031_);
  and (_0036_, _0035_, _0027_);
  nand (_0037_, _0036_, _0020_);
  nor (_0038_, _0002_, _1891_);
  nor (_0039_, _0038_, _1887_);
  and (_0040_, _0039_, _0005_);
  and (_0041_, _0040_, _1874_);
  nand (_0042_, _0041_, _1843_);
  and (_0043_, _0042_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [1]);
  nand (_0044_, _0043_, _0037_);
  and (_0045_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [1], _1271_);
  nor (_0046_, _0045_, _1665_);
  and (_0047_, _0046_, _1759_);
  nand (_0048_, _0047_, _0044_);
  or (_0049_, _0048_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [0]);
  and (_0050_, _0049_, _1759_);
  and (_0051_, \xm8051_golden_model_1.aes_bytes_processed [4], \xm8051_golden_model_1.aes_bytes_processed [5]);
  and (_0052_, _0051_, \xm8051_golden_model_1.aes_bytes_processed [6]);
  and (_0053_, _0052_, \xm8051_golden_model_1.aes_bytes_processed [7]);
  and (_0054_, _0053_, \xm8051_golden_model_1.aes_bytes_processed [8]);
  and (_0055_, _0054_, \xm8051_golden_model_1.aes_bytes_processed [9]);
  and (_0056_, _0055_, \xm8051_golden_model_1.aes_bytes_processed [10]);
  and (_0057_, _0056_, \xm8051_golden_model_1.aes_bytes_processed [11]);
  and (_0058_, _0057_, \xm8051_golden_model_1.aes_bytes_processed [12]);
  and (_0059_, _0058_, \xm8051_golden_model_1.aes_bytes_processed [13]);
  and (_0060_, _0059_, _0050_);
  nand (_0061_, _0060_, \xm8051_golden_model_1.aes_bytes_processed [14]);
  or (_0063_, _0060_, \xm8051_golden_model_1.aes_bytes_processed [14]);
  and (_0065_, _0063_, _0061_);
  or (_0066_, _0065_, _1616_);
  and (_0067_, _1664_, _1340_);
  not (_0068_, _0067_);
  and (_0069_, _0068_, \xm8051_golden_model_1.aes_bytes_processed [14]);
  nor (_0070_, \xm8051_golden_model_1.sha_state [1], _1369_);
  and (_0071_, _0070_, _1336_);
  and (_0072_, _0071_, _0069_);
  or (_0073_, _0072_, _1596_);
  not (_0074_, _0071_);
  and (_0075_, _1595_, _0070_);
  and (_0076_, _1370_, _1336_);
  and (_0077_, _0069_, _0076_);
  or (_0078_, _0077_, _0075_);
  not (_0079_, _0076_);
  and (_0080_, \xm8051_golden_model_1.sha_state [1], \xm8051_golden_model_1.sha_state [0]);
  and (_0081_, _0080_, _1336_);
  not (_0082_, _0081_);
  and (_0083_, _0080_, _1595_);
  or (_0084_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [14]);
  and (_0085_, _0084_, _0082_);
  and (_0086_, _1595_, _1370_);
  and (_0087_, _0081_, _0069_);
  or (_0088_, _0087_, _0086_);
  or (_0089_, _0088_, _0085_);
  and (_0090_, _0089_, _0079_);
  or (_0091_, _0090_, _0078_);
  and (_0092_, _0091_, _0074_);
  or (_0093_, _0092_, _0073_);
  and (_0094_, _0093_, _0066_);
  or (_0095_, _0094_, _1757_);
  not (_0096_, _1757_);
  or (_0097_, _0069_, _0096_);
  and (_0098_, _0097_, _1330_);
  and (_1892_[14], _0098_, _0095_);
  and (_0099_, _1363_, proc_data_in[2]);
  not (_0100_, \xm8051_golden_model_1.aes_len [10]);
  nor (_0101_, _1363_, _0100_);
  or (_0102_, _0101_, _0099_);
  and (_1893_[10], _0102_, _1330_);
  and (_0103_, _1291_, _1372_);
  nand (_0104_, _0103_, _1294_);
  and (_0105_, _1299_, _1330_);
  and (_0062_, _0105_, _0104_);
  not (_0106_, _0103_);
  and (_0107_, _1299_, _1294_);
  and (_0108_, _0107_, _0106_);
  and (_0109_, _0108_, _1292_);
  not (_0110_, _0108_);
  and (_0111_, _0110_, \oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbit_holder [1]);
  or (_0112_, _0111_, _0109_);
  and (_0064_, _0112_, _1330_);
  not (_0113_, \xm8051_golden_model_1.aes_bytes_processed [2]);
  or (_0114_, _0113_, rst);
  nor (_1892_[2], _0114_, _0067_);
  or (_0115_, _0110_, _1302_);
  or (_0116_, _0108_, \oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbit_holder [0]);
  and (_0117_, _0116_, _1330_);
  and (_0120_, _0117_, _0115_);
  not (_0118_, \xm8051_golden_model_1.aes_bytes_processed [10]);
  and (_0119_, _0055_, _0118_);
  nor (_0121_, _0055_, _0118_);
  or (_0122_, _0121_, _0119_);
  nand (_0123_, _0122_, _0050_);
  or (_0124_, _0050_, _0118_);
  nand (_0125_, _0124_, _0123_);
  or (_0126_, _0125_, _1616_);
  nor (_0127_, _0067_, _0118_);
  and (_0128_, _0127_, _0071_);
  or (_0129_, _0128_, _1596_);
  and (_0130_, _0127_, _0076_);
  or (_0131_, _0130_, _0075_);
  or (_0132_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [10]);
  and (_0133_, _0132_, _0082_);
  and (_0134_, _0127_, _0081_);
  or (_0135_, _0134_, _0086_);
  or (_0136_, _0135_, _0133_);
  and (_0137_, _0136_, _0079_);
  or (_0138_, _0137_, _0131_);
  and (_0139_, _0138_, _0074_);
  or (_0140_, _0139_, _0129_);
  and (_0141_, _0140_, _0126_);
  or (_0142_, _0141_, _1757_);
  or (_0143_, _0127_, _0096_);
  and (_0144_, _0143_, _1330_);
  and (_1892_[10], _0144_, _0142_);
  nor (_0145_, _1513_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [13]);
  and (_0146_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [12], _1529_);
  or (_0147_, _0146_, _0145_);
  and (_0148_, _1513_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [13]);
  and (_0149_, _1514_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [12]);
  or (_0150_, _0149_, _0148_);
  and (_0151_, _1538_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [14]);
  and (_0152_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [14], _1547_);
  and (_0153_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [15], _1537_);
  nor (_0154_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [15], _1537_);
  or (_0155_, _0154_, _0153_);
  or (_0156_, _0155_, _0152_);
  or (_0157_, _0156_, _0151_);
  or (_0158_, _0157_, _0150_);
  or (_0159_, _0158_, _0147_);
  and (_0160_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [11], _1492_);
  and (_0161_, _1493_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [10]);
  nor (_0162_, _0161_, _0160_);
  and (_0163_, _1491_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [11]);
  and (_0164_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [10], _1504_);
  nor (_0165_, _0164_, _0163_);
  nand (_0166_, _0165_, _0162_);
  and (_0167_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [9], _1468_);
  nor (_0168_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [8], _1483_);
  nor (_0169_, _0168_, _0167_);
  and (_0170_, _1467_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [9]);
  and (_0171_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [8], _1483_);
  nor (_0172_, _0171_, _0170_);
  nand (_0173_, _0172_, _0169_);
  or (_0174_, _0173_, _0166_);
  nor (_0175_, _0174_, _0159_);
  not (_0176_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [7]);
  or (_0177_, _0176_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [7]);
  or (_0178_, _1457_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [6]);
  and (_0179_, _0178_, _0177_);
  and (_0180_, _0176_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [7]);
  and (_0181_, _1457_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [6]);
  nor (_0183_, _0181_, _0180_);
  nand (_0184_, _0183_, _0179_);
  and (_0185_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [5], _1436_);
  and (_0186_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [4], _1427_);
  nor (_0187_, _0186_, _0185_);
  and (_0188_, _1435_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [5]);
  and (_0189_, _1426_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [4]);
  nor (_0190_, _0189_, _0188_);
  nand (_0191_, _0190_, _0187_);
  nor (_0192_, _0191_, _0184_);
  or (_0193_, _1407_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [3]);
  or (_0194_, _1417_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [2]);
  and (_0195_, _0194_, _0193_);
  and (_0196_, _1407_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [3]);
  and (_0197_, _1417_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [2]);
  nor (_0198_, _0197_, _0196_);
  and (_0199_, _0198_, _0195_);
  or (_0200_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [1], _1398_);
  and (_0201_, _1389_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [0]);
  and (_0202_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [1], _1398_);
  or (_0203_, _0202_, _0201_);
  nand (_0204_, _0203_, _0200_);
  nand (_0205_, _0204_, _0199_);
  or (_0206_, _0196_, _0195_);
  nand (_0207_, _0206_, _0205_);
  nand (_0208_, _0207_, _0192_);
  or (_0209_, _0180_, _0179_);
  or (_0210_, _0188_, _0187_);
  or (_0211_, _0210_, _0184_);
  and (_0212_, _0211_, _0209_);
  nand (_0213_, _0212_, _0208_);
  nand (_0214_, _0213_, _0175_);
  or (_0215_, _0170_, _0169_);
  or (_0216_, _0215_, _0166_);
  or (_0217_, _0163_, _0162_);
  and (_0218_, _0217_, _0216_);
  or (_0219_, _0159_, _0218_);
  not (_0220_, _0151_);
  nor (_0221_, _0220_, _0153_);
  nor (_0222_, _0221_, _0154_);
  not (_0223_, _0149_);
  nor (_0224_, _0223_, _0145_);
  nor (_0225_, _0224_, _0148_);
  or (_0226_, _0225_, _0157_);
  and (_0227_, _0226_, _0222_);
  and (_0228_, _0227_, _0219_);
  and (_0229_, _0228_, _0214_);
  or (_0230_, _1389_, \oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [0]);
  nand (_0231_, _0230_, _0200_);
  nor (_0232_, _0231_, _0203_);
  and (_0233_, _0232_, _0199_);
  and (_0234_, _0233_, _0192_);
  nand (_0235_, _0234_, _0175_);
  nand (_0236_, _0235_, ABINPUT000[161]);
  or (_0237_, _0236_, _0229_);
  and (_0238_, _0237_, _1373_);
  or (_0239_, _0238_, _1571_);
  and (_0240_, _1560_, _1390_);
  or (_0241_, _0240_, _0239_);
  and (_0182_, _0241_, _1330_);
  nand (_0242_, _0058_, _0050_);
  and (_0243_, _0242_, \xm8051_golden_model_1.aes_bytes_processed [13]);
  nor (_0244_, _0242_, \xm8051_golden_model_1.aes_bytes_processed [13]);
  or (_0245_, _0244_, _0243_);
  or (_0246_, _0245_, _1616_);
  and (_0247_, _0068_, \xm8051_golden_model_1.aes_bytes_processed [13]);
  and (_0248_, _0247_, _0071_);
  or (_0249_, _0248_, _1596_);
  and (_0250_, _0247_, _0076_);
  or (_0251_, _0250_, _0075_);
  or (_0252_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [13]);
  and (_0253_, _0252_, _0082_);
  and (_0254_, _0247_, _0081_);
  or (_0255_, _0254_, _0086_);
  or (_0256_, _0255_, _0253_);
  and (_0257_, _0256_, _0079_);
  or (_0258_, _0257_, _0251_);
  and (_0259_, _0258_, _0074_);
  or (_0260_, _0259_, _0249_);
  and (_0261_, _0260_, _0246_);
  or (_0262_, _0261_, _1757_);
  or (_0263_, _0247_, _0096_);
  and (_0264_, _0263_, _1330_);
  and (_1892_[13], _0264_, _0262_);
  and (_0279_, _1786_, _1330_);
  and (_0265_, _0057_, _0050_);
  or (_0266_, _0265_, \xm8051_golden_model_1.aes_bytes_processed [12]);
  and (_0267_, _0266_, _0242_);
  or (_0268_, _0267_, _1597_);
  and (_0269_, _0068_, \xm8051_golden_model_1.aes_bytes_processed [12]);
  or (_0270_, _0269_, _0079_);
  or (_0271_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [12]);
  and (_0272_, _0271_, _0082_);
  or (_0273_, _0272_, _0086_);
  and (_0274_, _0273_, _0270_);
  or (_0275_, _0274_, _0075_);
  and (_0276_, _0275_, _0267_);
  not (_0277_, _0086_);
  and (_0278_, _0269_, _0081_);
  not (_0280_, _0083_);
  and (_0281_, _0272_, _0280_);
  or (_0282_, _0281_, _0278_);
  and (_0283_, _0282_, _0277_);
  or (_0284_, _0283_, _0076_);
  not (_0285_, _0075_);
  and (_0286_, _0270_, _0285_);
  and (_0287_, _0286_, _0284_);
  or (_0288_, _0287_, _0276_);
  and (_0289_, _0288_, _0074_);
  and (_0290_, _0269_, _0071_);
  or (_0291_, _0290_, _1596_);
  or (_0292_, _0291_, _0289_);
  and (_0293_, _0292_, _0268_);
  or (_0294_, _0293_, _1757_);
  or (_0295_, _0269_, _0096_);
  and (_0296_, _0295_, _1330_);
  and (_1892_[12], _0296_, _0294_);
  and (_0318_, _1833_, _1330_);
  and (_0297_, _1343_, proc_addr[1]);
  and (_0298_, _0297_, _1309_);
  and (_0299_, _0298_, _1377_);
  and (_0300_, _0299_, _1332_);
  nor (_0301_, _0300_, _1389_);
  and (_0302_, _0300_, proc_data_in[0]);
  or (_0303_, _0302_, _0301_);
  and (_0331_, _0303_, _1330_);
  nor (_0304_, _0300_, _1398_);
  and (_0305_, _0300_, proc_data_in[1]);
  or (_0306_, _0305_, _0304_);
  and (_0343_, _0306_, _1330_);
  and (_0307_, _1349_, proc_data_in[1]);
  not (_0308_, \xm8051_golden_model_1.aes_len [1]);
  nor (_0309_, _1349_, _0308_);
  or (_0310_, _0309_, _0307_);
  and (_1893_[1], _0310_, _1330_);
  and (_0375_, _1402_, _1330_);
  not (_0311_, \xm8051_golden_model_1.aes_state [1]);
  and (_0312_, _0311_, \xm8051_golden_model_1.aes_state [0]);
  and (_0313_, _0070_, _0312_);
  and (_0314_, _0050_, _0313_);
  and (_0315_, _0312_, _1370_);
  and (_0316_, _0050_, _0315_);
  and (_0317_, _0080_, _0312_);
  nand (_0319_, _0317_, _0050_);
  or (_0320_, _0083_, _0311_);
  nand (_0321_, _0320_, _0319_);
  and (_0322_, _0321_, _0277_);
  or (_0323_, _0322_, _0316_);
  and (_0324_, _0323_, _0285_);
  or (_0325_, _0324_, _0314_);
  and (_0326_, _0325_, _1597_);
  and (_0327_, _1318_, _0311_);
  and (_0328_, _0327_, \xm8051_golden_model_1.aes_state [0]);
  and (_0329_, _0050_, _0328_);
  nand (_0330_, _0049_, _1759_);
  and (_0332_, _0330_, _1595_);
  or (_0333_, _0332_, _0329_);
  or (_0334_, _0333_, _0326_);
  and (_1894_[1], _0334_, _1330_);
  and (_0335_, _1575_, \xm8051_golden_model_1.sha_bytes_processed [6]);
  or (_0336_, _0335_, \xm8051_golden_model_1.sha_bytes_processed [7]);
  and (_0337_, _0336_, _1577_);
  and (_0338_, _0337_, _1370_);
  and (_0339_, _1318_, \xm8051_golden_model_1.sha_bytes_processed [7]);
  and (_0340_, _0339_, _1329_);
  and (_0341_, \xm8051_golden_model_1.sha_state [0], \xm8051_golden_model_1.sha_bytes_processed [7]);
  or (_0342_, _0341_, _0340_);
  or (_0344_, _0342_, _0338_);
  and (_1895_[7], _0344_, _1330_);
  nand (_0345_, \oc8051_xiommu_impl_1.oc8051_xram_i.cnt [0], _1330_);
  or (_0409_, _0345_, _1696_);
  nor (_0346_, _0300_, _1407_);
  and (_0347_, _0300_, proc_data_in[3]);
  or (_0348_, _0347_, _0346_);
  and (_0442_, _0348_, _1330_);
  and (_0349_, _1363_, proc_data_in[5]);
  not (_0350_, \xm8051_golden_model_1.aes_len [13]);
  nor (_0351_, _1363_, _0350_);
  or (_0352_, _0351_, _0349_);
  and (_1893_[13], _0352_, _1330_);
  nor (_0353_, _1639_, _1869_);
  and (_0354_, _1639_, proc_data_in[5]);
  or (_0355_, _0354_, _0353_);
  and (_0506_, _0355_, _1330_);
  and (_0542_, _0048_, _1330_);
  and (_0356_, _1386_, _1383_);
  and (_0357_, _0356_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [4]);
  or (_0358_, _0356_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [4]);
  and (_0359_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0], _1330_);
  nand (_0360_, _0359_, _0358_);
  nor (_0553_, _0360_, _0357_);
  nor (_0361_, _0300_, _1426_);
  and (_0362_, _0300_, proc_data_in[4]);
  or (_0363_, _0362_, _0361_);
  and (_0564_, _0363_, _1330_);
  and (_0573_, _1543_, _1330_);
  and (_0364_, _1363_, proc_data_in[6]);
  not (_0365_, \xm8051_golden_model_1.aes_len [14]);
  nor (_0366_, _1363_, _0365_);
  or (_0367_, _0366_, _0364_);
  and (_1893_[14], _0367_, _1330_);
  not (_0368_, \xm8051_golden_model_1.aes_bytes_processed [9]);
  and (_0369_, _0054_, _0368_);
  nor (_0370_, _0054_, _0368_);
  nor (_0371_, _0370_, _0369_);
  nor (_0372_, _0371_, _0330_);
  and (_0373_, _0330_, \xm8051_golden_model_1.aes_bytes_processed [9]);
  nor (_0374_, _0373_, _0372_);
  nand (_0376_, _0374_, _1595_);
  nor (_0377_, _0067_, _0368_);
  and (_0378_, _0377_, _0076_);
  or (_0379_, _0378_, _0075_);
  or (_0380_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [9]);
  and (_0381_, _0380_, _0082_);
  and (_0382_, _0377_, _0081_);
  or (_0383_, _0382_, _0086_);
  or (_0384_, _0383_, _0381_);
  and (_0385_, _0384_, _0079_);
  or (_0386_, _0385_, _0379_);
  and (_0387_, _0386_, _0074_);
  and (_0388_, _0377_, _0071_);
  or (_0389_, _0388_, _1596_);
  or (_0390_, _0389_, _0387_);
  and (_0391_, _0390_, _0376_);
  or (_0392_, _0391_, _1757_);
  or (_0393_, _0377_, _0096_);
  and (_0394_, _0393_, _1330_);
  and (_1892_[9], _0394_, _0392_);
  not (_0395_, \xm8051_golden_model_1.sha_len [15]);
  and (_0396_, _0298_, _1314_);
  and (_0397_, _0396_, proc_addr[0]);
  nor (_0398_, _0397_, _0395_);
  and (_0399_, _0397_, proc_data_in[7]);
  or (_0400_, _0399_, _1319_);
  or (_0401_, _0400_, _0398_);
  or (_0402_, _1318_, \xm8051_golden_model_1.sha_len [15]);
  and (_0403_, _0402_, _1330_);
  and (_1896_[15], _0403_, _0401_);
  nor (_0404_, _1639_, _1891_);
  and (_0405_, _1639_, proc_data_in[0]);
  or (_0406_, _0405_, _0404_);
  and (_0618_, _0406_, _1330_);
  and (_0407_, _0061_, \xm8051_golden_model_1.aes_bytes_processed [15]);
  nor (_0408_, _0061_, \xm8051_golden_model_1.aes_bytes_processed [15]);
  or (_0410_, _0408_, _0407_);
  nor (_0411_, _0083_, _0086_);
  and (_0412_, _0411_, _0285_);
  or (_0413_, _0412_, _0410_);
  or (_0414_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [15]);
  and (_0415_, _0414_, _0082_);
  and (_0416_, _0068_, \xm8051_golden_model_1.aes_bytes_processed [15]);
  and (_0417_, _0416_, _0081_);
  or (_0418_, _0417_, _0086_);
  or (_0419_, _0418_, _0415_);
  and (_0420_, _0419_, _0079_);
  and (_0421_, _0416_, _0076_);
  or (_0422_, _0421_, _0075_);
  or (_0423_, _0422_, _0420_);
  and (_0424_, _0423_, _0413_);
  or (_0425_, _0424_, _0071_);
  or (_0426_, _0416_, _0074_);
  and (_0427_, _0426_, _1597_);
  and (_0428_, _0427_, _0425_);
  and (_0429_, _0410_, _1596_);
  or (_0430_, _0429_, _1757_);
  or (_0431_, _0430_, _0428_);
  or (_0432_, _0416_, _0096_);
  and (_0433_, _0432_, _1330_);
  and (_1892_[15], _0433_, _0431_);
  nor (_0434_, _1578_, \xm8051_golden_model_1.sha_bytes_processed [9]);
  nor (_0435_, _0434_, _1605_);
  and (_0436_, _0435_, _1370_);
  not (_0437_, \xm8051_golden_model_1.sha_state [1]);
  and (_0438_, _1329_, _0437_);
  or (_0439_, _0438_, \xm8051_golden_model_1.sha_state [0]);
  and (_0440_, _0439_, \xm8051_golden_model_1.sha_bytes_processed [9]);
  or (_0441_, _0440_, _0436_);
  and (_1895_[9], _0441_, _1330_);
  nand (_0443_, _1607_, _1602_);
  and (_0444_, _0443_, _1608_);
  and (_0445_, _0444_, _1370_);
  and (_0446_, _1318_, \xm8051_golden_model_1.sha_bytes_processed [12]);
  and (_0447_, _0446_, _1329_);
  and (_0448_, \xm8051_golden_model_1.sha_state [0], \xm8051_golden_model_1.sha_bytes_processed [12]);
  or (_0449_, _0448_, _0447_);
  or (_0450_, _0449_, _0445_);
  and (_1895_[12], _0450_, _1330_);
  and (_0652_, _1775_, _1666_);
  and (_0451_, \xm8051_golden_model_1.sha_bytes_processed [3], _1330_);
  and (_1895_[3], _0451_, _1329_);
  not (_0452_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [10]);
  nor (_0453_, _1359_, _0452_);
  and (_0454_, _1359_, proc_data_in[2]);
  or (_0455_, _0454_, _0453_);
  and (_0680_, _0455_, _1330_);
  and (_0456_, _0065_, _0365_);
  nor (_0457_, _0065_, _0365_);
  nor (_0458_, _0457_, _0456_);
  not (_0459_, \xm8051_golden_model_1.aes_len [15]);
  nand (_0460_, _0410_, _0459_);
  or (_0461_, _0410_, _0459_);
  and (_0462_, _0461_, _0460_);
  and (_0463_, _0462_, _0458_);
  nor (_0464_, _0245_, _0350_);
  nor (_0465_, _0267_, _1365_);
  or (_0466_, _0465_, _0464_);
  nand (_0467_, _0267_, _1365_);
  nand (_0468_, _0245_, _0350_);
  nand (_0469_, _0468_, _0467_);
  nor (_0470_, _0469_, _0466_);
  and (_0471_, _0470_, _0463_);
  not (_0472_, \xm8051_golden_model_1.aes_len [11]);
  nand (_0473_, _0056_, _0050_);
  and (_0474_, _0473_, \xm8051_golden_model_1.aes_bytes_processed [11]);
  nor (_0475_, _0473_, \xm8051_golden_model_1.aes_bytes_processed [11]);
  or (_0476_, _0475_, _0474_);
  or (_0477_, _0476_, _0472_);
  nand (_0478_, _0476_, _0472_);
  and (_0479_, _0478_, _0477_);
  and (_0480_, _0125_, _0100_);
  nor (_0481_, _0125_, _0100_);
  nor (_0482_, _0481_, _0480_);
  and (_0483_, _0482_, _0479_);
  not (_0484_, \xm8051_golden_model_1.aes_len [8]);
  nand (_0485_, _0054_, _0050_);
  not (_0486_, \xm8051_golden_model_1.aes_bytes_processed [8]);
  nand (_0487_, _0053_, _0050_);
  nand (_0488_, _0487_, _0486_);
  and (_0489_, _0488_, _0485_);
  nor (_0490_, _0489_, _0484_);
  and (_0491_, _0489_, _0484_);
  nor (_0492_, _0491_, _0490_);
  or (_0493_, _0374_, \xm8051_golden_model_1.aes_len [9]);
  nand (_0494_, _0374_, \xm8051_golden_model_1.aes_len [9]);
  and (_0495_, _0494_, _0493_);
  and (_0496_, _0495_, _0492_);
  and (_0497_, _0496_, _0483_);
  nand (_0498_, _0497_, _0471_);
  not (_0499_, \xm8051_golden_model_1.aes_len [7]);
  and (_0500_, _0052_, _0050_);
  or (_0501_, _0500_, \xm8051_golden_model_1.aes_bytes_processed [7]);
  and (_0502_, _0501_, _0487_);
  nor (_0503_, _0502_, _0499_);
  not (_0504_, \xm8051_golden_model_1.aes_len [6]);
  nand (_0505_, _0051_, _0050_);
  nand (_0507_, _0505_, \xm8051_golden_model_1.aes_bytes_processed [6]);
  or (_0509_, _0505_, \xm8051_golden_model_1.aes_bytes_processed [6]);
  nand (_0510_, _0509_, _0507_);
  and (_0511_, _0510_, _0504_);
  nor (_0512_, _0511_, _0503_);
  nand (_0513_, _0502_, _0499_);
  or (_0514_, _0510_, _0504_);
  and (_0515_, _0514_, _0513_);
  and (_0516_, _0515_, _0512_);
  not (_0517_, \xm8051_golden_model_1.aes_len [5]);
  nor (_0518_, \xm8051_golden_model_1.aes_bytes_processed [4], \xm8051_golden_model_1.aes_bytes_processed [5]);
  nor (_0519_, _0518_, _0051_);
  or (_0520_, _0519_, _0330_);
  or (_0521_, _0050_, \xm8051_golden_model_1.aes_bytes_processed [5]);
  and (_0522_, _0521_, _0520_);
  and (_0523_, _0522_, _0517_);
  nand (_0524_, _0521_, _0520_);
  and (_0525_, _0524_, \xm8051_golden_model_1.aes_len [5]);
  or (_0526_, _0050_, \xm8051_golden_model_1.aes_bytes_processed [4]);
  not (_0527_, \xm8051_golden_model_1.aes_bytes_processed [4]);
  or (_0528_, _0330_, _0527_);
  and (_0529_, _0528_, _0526_);
  or (_0530_, _0529_, _1351_);
  nand (_0531_, _0529_, _1351_);
  nand (_0532_, _0531_, _0530_);
  or (_0533_, _0532_, _0525_);
  nor (_0534_, _0533_, _0523_);
  nand (_0535_, _0534_, _0516_);
  not (_0536_, \xm8051_golden_model_1.aes_bytes_processed [3]);
  and (_0537_, _0536_, \xm8051_golden_model_1.aes_len [3]);
  and (_0538_, \xm8051_golden_model_1.aes_len [2], _0113_);
  nor (_0539_, _0538_, _0537_);
  nor (_0540_, _0536_, \xm8051_golden_model_1.aes_len [3]);
  nor (_0541_, \xm8051_golden_model_1.aes_len [2], _0113_);
  nor (_0543_, _0541_, _0540_);
  and (_0544_, _0543_, _0539_);
  not (_0545_, \xm8051_golden_model_1.aes_bytes_processed [1]);
  and (_0546_, \xm8051_golden_model_1.aes_len [1], _0545_);
  not (_0547_, \xm8051_golden_model_1.aes_bytes_processed [0]);
  or (_0548_, \xm8051_golden_model_1.aes_len [0], _0547_);
  and (_0549_, _0308_, \xm8051_golden_model_1.aes_bytes_processed [1]);
  nor (_0550_, _0549_, _0546_);
  and (_0551_, _0550_, _0548_);
  or (_0552_, _0551_, _0546_);
  and (_0554_, _0552_, _0544_);
  not (_0555_, _0540_);
  and (_0556_, _0555_, _0538_);
  or (_0557_, _0556_, _0537_);
  nor (_0558_, _0557_, _0554_);
  nor (_0559_, _0558_, _0535_);
  nor (_0560_, _0523_, _0530_);
  or (_0561_, _0560_, _0525_);
  and (_0562_, _0561_, _0516_);
  nor (_0563_, _0510_, _0504_);
  and (_0565_, _0563_, _0513_);
  or (_0566_, _0565_, _0503_);
  or (_0567_, _0566_, _0562_);
  nor (_0568_, _0567_, _0559_);
  nor (_0569_, _0568_, _0498_);
  nand (_0570_, _0493_, _0490_);
  nand (_0571_, _0570_, _0494_);
  and (_0572_, _0571_, _0483_);
  nand (_0574_, _0481_, _0478_);
  nand (_0575_, _0574_, _0477_);
  or (_0576_, _0575_, _0572_);
  and (_0577_, _0576_, _0471_);
  and (_0578_, _0468_, _0466_);
  and (_0579_, _0578_, _0463_);
  nand (_0580_, _0457_, _0460_);
  nand (_0581_, _0580_, _0461_);
  or (_0582_, _0581_, _0579_);
  or (_0583_, _0582_, _0577_);
  or (_0584_, _0583_, _0569_);
  nand (_0585_, \xm8051_golden_model_1.aes_len [0], _0547_);
  and (_0586_, _0551_, _0585_);
  nand (_0587_, _0586_, _0544_);
  or (_0588_, _0587_, _0535_);
  or (_0589_, _0588_, _0498_);
  and (_0590_, _0589_, _0584_);
  or (_0591_, _0590_, _0330_);
  and (_0592_, _0591_, _1595_);
  and (_0593_, _0071_, _0067_);
  and (_0594_, _0067_, _0076_);
  not (_0595_, \xm8051_golden_model_1.aes_state [0]);
  and (_0596_, \xm8051_golden_model_1.aes_state [1], _0595_);
  and (_0597_, _0596_, _1370_);
  and (_0598_, _0050_, _0597_);
  or (_0599_, _0598_, _0315_);
  and (_0600_, _0081_, _0067_);
  and (_0601_, _0080_, _0596_);
  and (_0602_, _0601_, _0050_);
  nor (_0603_, _0083_, _0595_);
  or (_0604_, _0603_, _0602_);
  and (_0605_, _0604_, _0319_);
  or (_0606_, _0605_, _0600_);
  and (_0607_, _0606_, _0277_);
  nor (_0608_, _0607_, _0599_);
  nor (_0609_, _0608_, _0316_);
  or (_0610_, _0609_, _0594_);
  and (_0611_, _0610_, _0285_);
  and (_0612_, _0596_, _0070_);
  and (_0613_, _0612_, _0050_);
  or (_0614_, _0613_, _0313_);
  nor (_0615_, _0614_, _0611_);
  nor (_0616_, _0615_, _0314_);
  or (_0617_, _0616_, _0593_);
  and (_0619_, _0617_, _1597_);
  and (_0620_, _0596_, _1318_);
  and (_0621_, _0050_, _0620_);
  or (_0622_, _0621_, _0328_);
  or (_0623_, _0622_, _0619_);
  nor (_0624_, _0623_, _0592_);
  nor (_0625_, _0624_, _0329_);
  and (_0626_, _0067_, _1757_);
  or (_0627_, _0626_, _0625_);
  and (_1894_[0], _0627_, _1330_);
  and (_0701_, _1666_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [3]);
  nor (_0628_, _1639_, _1860_);
  and (_0629_, _1639_, proc_data_in[4]);
  or (_0630_, _0629_, _0628_);
  and (_0711_, _0630_, _1330_);
  not (_0631_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [14]);
  nor (_0632_, _1359_, _0631_);
  and (_0633_, _1359_, proc_data_in[6]);
  or (_0634_, _0633_, _0632_);
  and (_0723_, _0634_, _1330_);
  and (_0635_, _1349_, proc_data_in[5]);
  nor (_0636_, _1349_, _0517_);
  or (_0637_, _0636_, _0635_);
  and (_1893_[5], _0637_, _1330_);
  not (_0638_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [6]);
  nor (_0639_, _1639_, _0638_);
  and (_0640_, _1639_, proc_data_in[6]);
  or (_0641_, _0640_, _0639_);
  and (_0798_, _0641_, _1330_);
  nor (_0642_, _1605_, \xm8051_golden_model_1.sha_bytes_processed [10]);
  nor (_0643_, _0642_, _1606_);
  or (_0644_, _0643_, _1600_);
  or (_0645_, _1319_, \xm8051_golden_model_1.sha_bytes_processed [10]);
  or (_0646_, _1369_, \xm8051_golden_model_1.sha_bytes_processed [10]);
  and (_0647_, _0646_, _1330_);
  and (_0648_, _0647_, _0645_);
  and (_0649_, _0648_, _1329_);
  and (_1895_[10], _0649_, _0644_);
  and (_0650_, \xm8051_golden_model_1.sha_bytes_processed [2], _1330_);
  and (_1895_[2], _0650_, _1329_);
  not (_0651_, \xm8051_golden_model_1.sha_len [14]);
  nor (_0653_, _0397_, _0651_);
  and (_0654_, _0397_, proc_data_in[6]);
  or (_0655_, _0654_, _1319_);
  or (_0656_, _0655_, _0653_);
  or (_0657_, _1318_, \xm8051_golden_model_1.sha_len [14]);
  and (_0658_, _0657_, _1330_);
  and (_1896_[14], _0658_, _0656_);
  and (_0821_, _1825_, _1666_);
  and (_0835_, _1666_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [2]);
  not (_0659_, \xm8051_golden_model_1.sha_len [13]);
  nor (_0660_, _0397_, _0659_);
  and (_0661_, _0397_, proc_data_in[5]);
  or (_0662_, _0661_, _1319_);
  or (_0663_, _0662_, _0660_);
  or (_0664_, _1318_, \xm8051_golden_model_1.sha_len [13]);
  and (_0665_, _0664_, _1330_);
  and (_1896_[13], _0665_, _0663_);
  and (_0880_, _1666_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [1]);
  not (_0666_, \xm8051_golden_model_1.sha_len [12]);
  nor (_0667_, _0397_, _0666_);
  and (_0668_, _0397_, proc_data_in[4]);
  or (_0669_, _0668_, _1319_);
  or (_0670_, _0669_, _0667_);
  or (_0671_, _1318_, \xm8051_golden_model_1.sha_len [12]);
  and (_0672_, _0671_, _1330_);
  and (_1896_[12], _0672_, _0670_);
  and (_0673_, _0299_, proc_addr[0]);
  nor (_0674_, _0673_, _1483_);
  and (_0675_, _0673_, proc_data_in[0]);
  or (_0676_, _0675_, _0674_);
  and (_0908_, _0676_, _1330_);
  or (_0677_, _0502_, _0412_);
  or (_0678_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [7]);
  and (_0679_, _0678_, _0082_);
  and (_0681_, _0068_, \xm8051_golden_model_1.aes_bytes_processed [7]);
  and (_0682_, _0681_, _0081_);
  or (_0683_, _0682_, _0086_);
  or (_0684_, _0683_, _0679_);
  and (_0685_, _0684_, _0079_);
  and (_0686_, _0681_, _0076_);
  or (_0687_, _0686_, _0075_);
  or (_0688_, _0687_, _0685_);
  and (_0689_, _0688_, _0677_);
  or (_0690_, _0689_, _0071_);
  or (_0691_, _0681_, _0074_);
  and (_0692_, _0691_, _1597_);
  and (_0693_, _0692_, _0690_);
  and (_0694_, _0502_, _1596_);
  or (_0695_, _0694_, _1757_);
  or (_0696_, _0695_, _0693_);
  or (_0697_, _0681_, _0096_);
  and (_0698_, _0697_, _1330_);
  and (_1892_[7], _0698_, _0696_);
  and (_0699_, _1349_, proc_data_in[2]);
  not (_0700_, _1349_);
  and (_0702_, _0700_, \xm8051_golden_model_1.aes_len [2]);
  or (_0703_, _0702_, _0699_);
  and (_1893_[2], _0703_, _1330_);
  nor (_0704_, _0673_, _1547_);
  and (_0705_, _0673_, proc_data_in[6]);
  or (_0706_, _0705_, _0704_);
  and (_0920_, _0706_, _1330_);
  and (_0707_, _1349_, proc_data_in[6]);
  nor (_0708_, _1349_, _0504_);
  or (_0709_, _0708_, _0707_);
  and (_1893_[6], _0709_, _1330_);
  and (_0710_, _1363_, proc_data_in[7]);
  nor (_0712_, _1363_, _0459_);
  or (_0713_, _0712_, _0710_);
  and (_1893_[15], _0713_, _1330_);
  not (_0714_, \xm8051_golden_model_1.sha_len [11]);
  nor (_0715_, _0397_, _0714_);
  and (_0716_, _0397_, proc_data_in[3]);
  or (_0717_, _0716_, _1319_);
  or (_0718_, _0717_, _0715_);
  or (_0719_, _1318_, \xm8051_golden_model_1.sha_len [11]);
  and (_0720_, _0719_, _1330_);
  and (_1896_[11], _0720_, _0718_);
  not (_0721_, \xm8051_golden_model_1.sha_len [10]);
  nor (_0722_, _0397_, _0721_);
  and (_0724_, _0397_, proc_data_in[2]);
  or (_0725_, _0724_, _1319_);
  or (_0726_, _0725_, _0722_);
  or (_0727_, _1318_, \xm8051_golden_model_1.sha_len [10]);
  and (_0728_, _0727_, _1330_);
  and (_1896_[10], _0728_, _0726_);
  or (_0729_, _1606_, \xm8051_golden_model_1.sha_bytes_processed [11]);
  and (_0730_, _0729_, _1607_);
  or (_0731_, _0730_, _1600_);
  or (_0732_, _1319_, \xm8051_golden_model_1.sha_bytes_processed [11]);
  or (_0733_, _1369_, \xm8051_golden_model_1.sha_bytes_processed [11]);
  and (_0734_, _0733_, _1330_);
  and (_0735_, _0734_, _0732_);
  and (_0736_, _0735_, _1329_);
  and (_1895_[11], _0736_, _0731_);
  not (_0737_, \xm8051_golden_model_1.sha_len [9]);
  nor (_0738_, _0397_, _0737_);
  and (_0739_, _0397_, proc_data_in[1]);
  or (_0740_, _0739_, _1319_);
  or (_0741_, _0740_, _0738_);
  or (_0742_, _1318_, \xm8051_golden_model_1.sha_len [9]);
  and (_0743_, _0742_, _1330_);
  and (_1896_[9], _0743_, _0741_);
  or (_0744_, _0510_, _1616_);
  and (_0745_, _0068_, \xm8051_golden_model_1.aes_bytes_processed [6]);
  and (_0746_, _0745_, _0076_);
  or (_0747_, _0746_, _0075_);
  or (_0748_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [6]);
  and (_0749_, _0748_, _0082_);
  and (_0750_, _0745_, _0081_);
  or (_0751_, _0750_, _0086_);
  or (_0752_, _0751_, _0749_);
  and (_0753_, _0752_, _0079_);
  or (_0754_, _0753_, _0747_);
  and (_0755_, _0754_, _0074_);
  and (_0756_, _0745_, _0071_);
  or (_0757_, _0756_, _1596_);
  or (_0758_, _0757_, _0755_);
  and (_0759_, _0758_, _0744_);
  or (_0760_, _0759_, _1757_);
  or (_0761_, _0745_, _0096_);
  and (_0762_, _0761_, _1330_);
  and (_1892_[6], _0762_, _0760_);
  nor (_0763_, _1359_, _1790_);
  and (_0764_, _1359_, proc_data_in[4]);
  or (_0765_, _0764_, _0763_);
  and (_0979_, _0765_, _1330_);
  not (_0766_, \xm8051_golden_model_1.sha_len [8]);
  nor (_0767_, _0397_, _0766_);
  and (_0768_, _0397_, proc_data_in[0]);
  or (_0769_, _0768_, _1319_);
  or (_0770_, _0769_, _0767_);
  or (_0771_, _1318_, \xm8051_golden_model_1.sha_len [8]);
  and (_0772_, _0771_, _1330_);
  and (_1896_[8], _0772_, _0770_);
  and (_0773_, _0068_, \xm8051_golden_model_1.aes_bytes_processed [5]);
  or (_0774_, _0773_, _0079_);
  and (_0775_, _0774_, _0285_);
  or (_0776_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [5]);
  and (_0777_, _0776_, _0082_);
  or (_0778_, _0777_, _0086_);
  and (_0779_, _0778_, _0775_);
  or (_0780_, _0779_, _0075_);
  and (_0781_, _0780_, _0074_);
  or (_0782_, _0781_, _1596_);
  and (_0783_, _0782_, _0522_);
  and (_0784_, _0773_, _0071_);
  and (_0785_, _0773_, _0081_);
  and (_0786_, _0777_, _0280_);
  or (_0787_, _0786_, _0785_);
  and (_0788_, _0787_, _0277_);
  or (_0789_, _0788_, _0076_);
  and (_0790_, _0775_, _0074_);
  and (_0791_, _0790_, _0789_);
  or (_0792_, _0791_, _0784_);
  and (_0793_, _0792_, _1597_);
  or (_0794_, _0793_, _1757_);
  or (_0795_, _0794_, _0783_);
  or (_0796_, _0773_, _0096_);
  and (_0797_, _0796_, _1330_);
  and (_1892_[5], _0797_, _0795_);
  or (_0799_, _0529_, _1616_);
  nor (_0800_, _0067_, _0527_);
  and (_0801_, _0800_, _0076_);
  or (_0802_, _0801_, _0075_);
  or (_0803_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [4]);
  and (_0804_, _0803_, _0082_);
  and (_0805_, _0800_, _0081_);
  or (_0806_, _0805_, _0086_);
  or (_0807_, _0806_, _0804_);
  and (_0808_, _0807_, _0079_);
  or (_0809_, _0808_, _0802_);
  and (_0810_, _0809_, _0074_);
  and (_0811_, _0800_, _0071_);
  or (_0812_, _0811_, _1596_);
  or (_0813_, _0812_, _0810_);
  and (_0814_, _0813_, _0799_);
  or (_0815_, _0814_, _1757_);
  or (_0816_, _0800_, _0096_);
  and (_0817_, _0816_, _1330_);
  and (_1892_[4], _0817_, _0815_);
  or (_0818_, _0536_, rst);
  nor (_1892_[3], _0818_, _0067_);
  and (_1001_, _1795_, _1666_);
  nor (_0819_, _1359_, _1828_);
  and (_0820_, _1359_, proc_data_in[1]);
  or (_0822_, _0820_, _0819_);
  and (_1004_, _0822_, _1330_);
  and (_0823_, \oc8051_xiommu_impl_1.oc8051_xram_i.cnt [0], \oc8051_xiommu_impl_1.oc8051_xram_i.cnt [1]);
  or (_0824_, _0823_, _1635_);
  nor (_0825_, _1636_, rst);
  nand (_0826_, _0825_, _0824_);
  nor (_1006_, _0826_, _1696_);
  and (_0827_, _1363_, proc_data_in[3]);
  nor (_0828_, _1363_, _0472_);
  or (_0829_, _0828_, _0827_);
  and (_1893_[11], _0829_, _1330_);
  nor (_0830_, _0673_, _1537_);
  and (_0831_, _0673_, proc_data_in[7]);
  or (_0832_, _0831_, _0830_);
  and (_1010_, _0832_, _1330_);
  nor (_0833_, _0673_, _1467_);
  and (_0834_, _0673_, proc_data_in[1]);
  or (_0836_, _0834_, _0833_);
  and (_1014_, _0836_, _1330_);
  not (_0837_, \xm8051_golden_model_1.sha_len [7]);
  and (_0838_, _0396_, _1332_);
  nor (_0839_, _0838_, _0837_);
  and (_0840_, _0838_, proc_data_in[7]);
  or (_0841_, _0840_, _1319_);
  or (_0842_, _0841_, _0839_);
  or (_0843_, _1318_, \xm8051_golden_model_1.sha_len [7]);
  and (_0844_, _0843_, _1330_);
  and (_1896_[7], _0844_, _0842_);
  nor (_0845_, _0673_, _1529_);
  and (_0846_, _0673_, proc_data_in[4]);
  or (_0847_, _0846_, _0845_);
  and (_1023_, _0847_, _1330_);
  not (_0848_, \xm8051_golden_model_1.sha_len [6]);
  nor (_0849_, _0838_, _0848_);
  and (_0850_, _0838_, proc_data_in[6]);
  or (_0851_, _0850_, _1319_);
  or (_0852_, _0851_, _0849_);
  or (_0853_, _1318_, \xm8051_golden_model_1.sha_len [6]);
  and (_0854_, _0853_, _1330_);
  and (_1896_[6], _0854_, _0852_);
  and (_0855_, _1363_, proc_data_in[1]);
  not (_0856_, \xm8051_golden_model_1.aes_len [9]);
  nor (_0857_, _1363_, _0856_);
  or (_0858_, _0857_, _0855_);
  and (_1893_[9], _0858_, _1330_);
  or (_0859_, _0545_, rst);
  nor (_1892_[1], _0859_, _0067_);
  and (_0860_, _1363_, proc_data_in[0]);
  nor (_0861_, _1363_, _0484_);
  or (_0862_, _0861_, _0860_);
  and (_1893_[8], _0862_, _1330_);
  and (_0863_, _1598_, \xm8051_golden_model_1.sha_bytes_processed [6]);
  and (_0864_, _1575_, _1370_);
  nor (_0865_, _0864_, _0863_);
  nor (_0866_, _1336_, _1319_);
  and (_0867_, _0866_, _1616_);
  and (_0868_, _0335_, _1370_);
  or (_0869_, _0868_, _0867_);
  nor (_0870_, _0869_, _0865_);
  and (_0871_, _1329_, \xm8051_golden_model_1.sha_bytes_processed [6]);
  and (_0872_, _0871_, _0867_);
  or (_0873_, _0872_, _1757_);
  or (_0874_, _0873_, _0870_);
  or (_0875_, _0871_, _0096_);
  and (_0876_, _0875_, _1330_);
  and (_1895_[6], _0876_, _0874_);
  nor (_0877_, _0673_, _1491_);
  and (_0878_, _0673_, proc_data_in[3]);
  or (_0879_, _0878_, _0877_);
  and (_1072_, _0879_, _1330_);
  nor (_0881_, _0673_, _1504_);
  and (_0882_, _0673_, proc_data_in[2]);
  or (_0883_, _0882_, _0881_);
  and (_1077_, _0883_, _1330_);
  or (_0884_, _0547_, rst);
  nor (_1892_[0], _0884_, _0067_);
  not (_0885_, \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [13]);
  nor (_0886_, _0673_, _0885_);
  and (_0887_, _0673_, proc_data_in[5]);
  or (_0888_, _0887_, _0886_);
  and (_1092_, _0888_, _1330_);
  not (_0889_, \xm8051_golden_model_1.sha_len [5]);
  nor (_0890_, _0838_, _0889_);
  and (_0891_, _0838_, proc_data_in[5]);
  or (_0892_, _0891_, _1319_);
  or (_0893_, _0892_, _0890_);
  or (_0894_, _1318_, \xm8051_golden_model_1.sha_len [5]);
  and (_0895_, _0894_, _1330_);
  and (_1896_[5], _0895_, _0893_);
  not (_0896_, \xm8051_golden_model_1.sha_len [4]);
  nor (_0897_, _0838_, _0896_);
  and (_0898_, _0838_, proc_data_in[4]);
  or (_0899_, _0898_, _1319_);
  or (_0900_, _0899_, _0897_);
  or (_0901_, _1318_, \xm8051_golden_model_1.sha_len [4]);
  and (_0902_, _0901_, _1330_);
  and (_1896_[4], _0902_, _0900_);
  not (_0903_, \xm8051_golden_model_1.sha_len [3]);
  nor (_0904_, _0838_, _0903_);
  and (_0905_, _0838_, proc_data_in[3]);
  or (_0906_, _0905_, _1319_);
  or (_0907_, _0906_, _0904_);
  or (_0909_, _1318_, \xm8051_golden_model_1.sha_len [3]);
  and (_0910_, _0909_, _1330_);
  and (_1896_[3], _0910_, _0907_);
  or (_0911_, _0476_, _0412_);
  or (_0912_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [11]);
  and (_0913_, _0912_, _0082_);
  and (_0914_, _0068_, \xm8051_golden_model_1.aes_bytes_processed [11]);
  and (_0915_, _0914_, _0081_);
  or (_0916_, _0915_, _0086_);
  or (_0917_, _0916_, _0913_);
  and (_0918_, _0917_, _0079_);
  and (_0919_, _0914_, _0076_);
  or (_0921_, _0919_, _0075_);
  or (_0922_, _0921_, _0918_);
  and (_0923_, _0922_, _0911_);
  or (_0924_, _0923_, _0071_);
  or (_0925_, _0914_, _0074_);
  and (_0926_, _0925_, _1597_);
  and (_0927_, _0926_, _0924_);
  and (_0928_, _0476_, _1596_);
  or (_0929_, _0928_, _1757_);
  or (_0930_, _0929_, _0927_);
  or (_0931_, _0914_, _0096_);
  and (_0932_, _0931_, _1330_);
  and (_1892_[11], _0932_, _0930_);
  not (_0933_, \xm8051_golden_model_1.sha_len [2]);
  nor (_0934_, _0838_, _0933_);
  and (_0935_, _0838_, proc_data_in[2]);
  or (_0936_, _0935_, _1319_);
  or (_0937_, _0936_, _0934_);
  or (_0938_, _1318_, \xm8051_golden_model_1.sha_len [2]);
  and (_0939_, _0938_, _1330_);
  and (_1896_[2], _0939_, _0937_);
  not (_0940_, \xm8051_golden_model_1.sha_len [1]);
  nor (_0941_, _0838_, _0940_);
  and (_0942_, _0838_, proc_data_in[1]);
  or (_0943_, _0942_, _1319_);
  or (_0944_, _0943_, _0941_);
  or (_0945_, _1318_, \xm8051_golden_model_1.sha_len [1]);
  and (_0946_, _0945_, _1330_);
  and (_1896_[1], _0946_, _0944_);
  not (_0947_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [8]);
  nor (_0948_, _1359_, _0947_);
  and (_0949_, _1359_, proc_data_in[0]);
  or (_0950_, _0949_, _0948_);
  and (_1118_, _0950_, _1330_);
  not (_0951_, \xm8051_golden_model_1.sha_len [0]);
  nor (_0952_, _0838_, _0951_);
  and (_0953_, _0838_, proc_data_in[0]);
  or (_0954_, _0953_, _1319_);
  or (_0955_, _0954_, _0952_);
  or (_0956_, _1318_, \xm8051_golden_model_1.sha_len [0]);
  and (_0957_, _0956_, _1330_);
  and (_1896_[0], _0957_, _0955_);
  and (_1134_, _1854_, _1666_);
  and (_1137_, _1864_, _1330_);
  nor (_0958_, _0300_, _1457_);
  and (_0959_, _0300_, proc_data_in[6]);
  or (_0960_, _0959_, _0958_);
  and (_1139_, _0960_, _1330_);
  or (_0961_, _1329_, _0311_);
  nand (_0962_, _0961_, \xm8051_golden_model_1.sha_bytes_processed [15]);
  nand (_0963_, _0962_, _1614_);
  not (_0964_, \xm8051_golden_model_1.sha_bytes_processed [15]);
  nor (_0965_, _1614_, _0964_);
  nor (_0966_, _0965_, _0327_);
  and (_0967_, _0966_, _0963_);
  and (_0968_, _0327_, \xm8051_golden_model_1.sha_bytes_processed [15]);
  and (_0969_, _0968_, _1329_);
  or (_0970_, _0969_, _0967_);
  and (_1895_[15], _0970_, _1330_);
  nor (_0971_, _1359_, _1806_);
  and (_0972_, _1359_, proc_data_in[3]);
  or (_0973_, _0972_, _0971_);
  and (_1149_, _0973_, _1330_);
  or (_0974_, _1699_, \oc8051_xiommu_impl_1.aes_top_i.byte_counter [3]);
  and (_0975_, _0974_, _1649_);
  and (_1161_, _0975_, _1666_);
  and (_0976_, _1349_, proc_data_in[7]);
  nor (_0977_, _1349_, _0499_);
  or (_0978_, _0977_, _0976_);
  and (_1893_[7], _0978_, _1330_);
  nand (_0980_, _0357_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [5]);
  or (_0981_, _0357_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [5]);
  and (_0982_, _0981_, _0980_);
  and (_1198_, _0982_, _0359_);
  and (_0983_, _1564_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [2]);
  or (_0984_, _0983_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [3]);
  nand (_0985_, _0984_, _0359_);
  nor (_1201_, _0985_, _0356_);
  nor (_0986_, _1564_, _1563_);
  or (_0987_, _0986_, _1565_);
  and (_1203_, _0987_, _0359_);
  and (_0988_, _1383_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [0]);
  or (_0989_, _0988_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [1]);
  nand (_0990_, _0989_, _0359_);
  nor (_1205_, _0990_, _1564_);
  nor (_0991_, _1383_, \oc8051_xiommu_impl_1.sha_top_i.byte_counter [0]);
  nor (_0992_, _0991_, _0988_);
  and (_1210_, _0992_, _0359_);
  and (_1212_, _1573_, _1330_);
  and (_1215_, _1550_, _1330_);
  nor (_0993_, _0300_, _0176_);
  and (_0994_, _0300_, proc_data_in[7]);
  or (_0995_, _0994_, _0993_);
  and (_1219_, _0995_, _1330_);
  nor (_0996_, _0300_, _1435_);
  and (_0997_, _0300_, proc_data_in[5]);
  or (_0998_, _0997_, _0996_);
  and (_1222_, _0998_, _1330_);
  and (_0999_, _1649_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [1]);
  not (_1000_, _1355_);
  nand (_1002_, _1623_, _1000_);
  nor (_1003_, _1002_, _1649_);
  or (_1005_, _1003_, _0999_);
  and (_1225_, _1005_, _1330_);
  and (_1007_, _1700_, \oc8051_xiommu_impl_1.aes_top_i.byte_counter [0]);
  or (_1008_, _1007_, \oc8051_xiommu_impl_1.aes_top_i.byte_counter [1]);
  nand (_1009_, _1008_, _1666_);
  nor (_1231_, _1009_, _1701_);
  and (_1249_, _1525_, _1330_);
  and (_1253_, _1532_, _1330_);
  or (_1011_, _1634_, rst);
  or (_1012_, _1011_, _1635_);
  nor (_1254_, _1012_, _1696_);
  and (_1255_, _1499_, _1330_);
  and (_1256_, _1666_, \oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [0]);
  nor (_1013_, _0300_, _1417_);
  and (_1015_, _0300_, proc_data_in[2]);
  or (_1016_, _1015_, _1013_);
  and (_1257_, _1016_, _1330_);
  and (_1017_, _1705_, \xm8051_golden_model_1.sha_state [1]);
  or (_1018_, _1017_, _1370_);
  and (_1019_, \xm8051_golden_model_1.sha_bytes_processed [12], \xm8051_golden_model_1.sha_bytes_processed [13]);
  and (_1020_, _1708_, _1019_);
  and (_1021_, _1020_, _1612_);
  nor (_1022_, _1020_, _1612_);
  nor (_1024_, _1022_, _1021_);
  or (_1025_, _1024_, _1705_);
  or (_1026_, _1575_, _1612_);
  and (_1027_, _1026_, _1025_);
  or (_1028_, _1027_, \xm8051_golden_model_1.sha_len [14]);
  nand (_1029_, _1027_, \xm8051_golden_model_1.sha_len [14]);
  and (_1030_, _1029_, _1028_);
  and (_1031_, _1020_, \xm8051_golden_model_1.sha_bytes_processed [14]);
  and (_1032_, _1031_, _0964_);
  nor (_1033_, _1031_, _0964_);
  nor (_1034_, _1033_, _1032_);
  or (_1035_, _1034_, _1705_);
  or (_1036_, _1575_, _0964_);
  and (_1037_, _1036_, _1035_);
  or (_1038_, _1037_, \xm8051_golden_model_1.sha_len [15]);
  nand (_1039_, _1037_, \xm8051_golden_model_1.sha_len [15]);
  and (_1040_, _1039_, _1038_);
  nand (_1041_, _1040_, _1030_);
  or (_1042_, _1716_, _0659_);
  or (_1043_, _0444_, _0666_);
  and (_1044_, _1716_, _0659_);
  or (_1045_, _1044_, _1043_);
  and (_1046_, _1045_, _1042_);
  or (_1047_, _1046_, _1041_);
  nand (_1048_, _1039_, _1029_);
  nand (_1049_, _1048_, _1038_);
  and (_1050_, _1049_, _1047_);
  nand (_1051_, _0444_, _0666_);
  and (_1052_, _1051_, _1043_);
  and (_1053_, _1052_, _1042_);
  nor (_1054_, _1044_, _1041_);
  and (_1055_, _1054_, _1053_);
  and (_1056_, _0730_, _0714_);
  or (_1057_, _0730_, _0714_);
  or (_1058_, _0643_, _0721_);
  and (_1059_, _1058_, _1057_);
  or (_1060_, _1059_, _1056_);
  and (_1061_, _0643_, _0721_);
  nor (_1062_, _1061_, _1056_);
  and (_1063_, _1062_, _1059_);
  and (_1064_, _0435_, _0737_);
  or (_1065_, _0435_, _0737_);
  or (_1066_, _1580_, _0766_);
  and (_1067_, _1066_, _1065_);
  nor (_1068_, _1067_, _1064_);
  nand (_1069_, _1068_, _1063_);
  nand (_1070_, _1069_, _1060_);
  nand (_1071_, _1070_, _1055_);
  and (_1073_, _1071_, _1050_);
  nor (_1074_, _1575_, \xm8051_golden_model_1.sha_bytes_processed [6]);
  nor (_1075_, _1074_, _0335_);
  or (_1076_, _1075_, _0848_);
  nand (_1078_, _1075_, _0848_);
  nand (_1079_, _1078_, _1076_);
  and (_1080_, _0337_, _0837_);
  nor (_1081_, _0337_, _0837_);
  or (_1082_, _1081_, _1080_);
  or (_1083_, _1082_, _1079_);
  nor (_1084_, _0889_, \xm8051_golden_model_1.sha_bytes_processed [5]);
  nor (_1085_, _0896_, \xm8051_golden_model_1.sha_bytes_processed [4]);
  nor (_1086_, _1085_, _1084_);
  and (_1087_, _0896_, \xm8051_golden_model_1.sha_bytes_processed [4]);
  and (_1088_, _0889_, \xm8051_golden_model_1.sha_bytes_processed [5]);
  nor (_1089_, _1088_, _1087_);
  nand (_1090_, _1089_, _1086_);
  nor (_1091_, _1090_, _1083_);
  or (_1093_, _0903_, \xm8051_golden_model_1.sha_bytes_processed [3]);
  or (_1094_, _0933_, \xm8051_golden_model_1.sha_bytes_processed [2]);
  and (_1095_, _1094_, _1093_);
  and (_1096_, _0903_, \xm8051_golden_model_1.sha_bytes_processed [3]);
  and (_1097_, _0933_, \xm8051_golden_model_1.sha_bytes_processed [2]);
  nor (_1098_, _1097_, _1096_);
  and (_1099_, _1098_, _1095_);
  nor (_1100_, _0940_, \xm8051_golden_model_1.sha_bytes_processed [1]);
  and (_1101_, _0951_, \xm8051_golden_model_1.sha_bytes_processed [0]);
  and (_1102_, _0940_, \xm8051_golden_model_1.sha_bytes_processed [1]);
  or (_1103_, _1102_, _1100_);
  nor (_1104_, _1103_, _1101_);
  or (_1105_, _1104_, _1100_);
  nand (_1106_, _1105_, _1099_);
  or (_1107_, _1096_, _1094_);
  and (_1108_, _1107_, _1093_);
  nand (_1109_, _1108_, _1106_);
  nand (_1110_, _1109_, _1091_);
  or (_1111_, _1088_, _1086_);
  or (_1112_, _1111_, _1083_);
  nor (_1113_, _1076_, _1080_);
  nor (_1114_, _1113_, _1081_);
  and (_1115_, _1114_, _1112_);
  nand (_1116_, _1115_, _1110_);
  and (_1117_, _1580_, _0766_);
  nor (_1119_, _1117_, _1064_);
  and (_1120_, _1119_, _1067_);
  and (_1121_, _1120_, _1063_);
  and (_1122_, _1121_, _1055_);
  nand (_1123_, _1122_, _1116_);
  and (_1124_, _1123_, _1073_);
  not (_1125_, _0864_);
  or (_1126_, _0951_, \xm8051_golden_model_1.sha_bytes_processed [0]);
  and (_1127_, _1126_, _1099_);
  and (_1128_, _1127_, _1104_);
  and (_1129_, _1128_, _1091_);
  and (_1130_, _1129_, _1122_);
  or (_1131_, _1130_, _1125_);
  or (_1132_, _1131_, _1124_);
  and (_1133_, _1132_, _1018_);
  and (_1135_, _0070_, _1575_);
  or (_1136_, _1135_, _1133_);
  and (_1897_[1], _1136_, _1330_);
  and (_1258_, _1507_, _1330_);
  and (_1259_, _1479_, _1330_);
  and (_1260_, _1486_, _1330_);
  and (_1261_, _1453_, _1330_);
  and (_1262_, _1460_, _1330_);
  and (_1263_, _1443_, _1330_);
  and (_1264_, _1431_, _1330_);
  and (_1265_, _1413_, _1330_);
  and (_1266_, _1420_, _1330_);
  and (_1138_, _1349_, proc_data_in[3]);
  and (_1140_, _0700_, \xm8051_golden_model_1.aes_len [3]);
  or (_1141_, _1140_, _1138_);
  and (_1893_[3], _1141_, _1330_);
  and (_1142_, \xm8051_golden_model_1.sha_bytes_processed [4], _1330_);
  and (_1895_[4], _1142_, _1329_);
  or (_1143_, _1700_, \oc8051_xiommu_impl_1.aes_top_i.byte_counter [0]);
  nand (_1144_, _1143_, _1666_);
  nor (_1267_, _1144_, _1007_);
  and (_1145_, _1705_, \xm8051_golden_model_1.sha_state [0]);
  nand (_1146_, _1125_, _1329_);
  or (_1147_, _1146_, _1145_);
  and (_1897_[0], _1147_, _1330_);
  nor (_1148_, _1639_, _1844_);
  and (_1150_, _1639_, proc_data_in[7]);
  or (_1151_, _1150_, _1148_);
  and (_1268_, _1151_, _1330_);
  and (_1269_, _1813_, _1666_);
  or (_1152_, _0489_, _1616_);
  nor (_1153_, _0067_, _0486_);
  and (_1154_, _1153_, _0076_);
  or (_1155_, _1154_, _0075_);
  or (_1156_, _0083_, \xm8051_golden_model_1.aes_bytes_processed [8]);
  and (_1157_, _1156_, _0082_);
  and (_1158_, _1153_, _0081_);
  or (_1159_, _1158_, _0086_);
  or (_1160_, _1159_, _1157_);
  and (_1162_, _1160_, _0079_);
  or (_1163_, _1162_, _1155_);
  and (_1164_, _1163_, _0074_);
  and (_1165_, _1153_, _0071_);
  or (_1166_, _1165_, _1596_);
  or (_1167_, _1166_, _1164_);
  and (_1168_, _1167_, _1152_);
  or (_1169_, _1168_, _1757_);
  or (_1170_, _1153_, _0096_);
  and (_1171_, _1170_, _1330_);
  and (_1892_[8], _1171_, _1169_);
  nand (_1172_, proc_stb_r, _1270_);
  or (_1173_, _1172_, _1306_);
  and (_1174_, _1173_, proc_stb_valid);
  or (_1175_, \xm8051_golden_model_1.aes_len [1], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [1]);
  nand (_1176_, \xm8051_golden_model_1.aes_len [1], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [1]);
  and (_1177_, _1176_, _1175_);
  or (_1178_, \xm8051_golden_model_1.aes_len [0], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [0]);
  nand (_1179_, \xm8051_golden_model_1.aes_len [0], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [0]);
  and (_1180_, _1179_, _1178_);
  or (_1181_, _1180_, _1177_);
  nand (_1182_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [2], \xm8051_golden_model_1.aes_len [2]);
  or (_1183_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [2], \xm8051_golden_model_1.aes_len [2]);
  and (_1184_, _1183_, _1182_);
  or (_1185_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [3], \xm8051_golden_model_1.aes_len [3]);
  nand (_1186_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [3], \xm8051_golden_model_1.aes_len [3]);
  and (_1187_, _1186_, _1185_);
  or (_1188_, _1187_, _1184_);
  or (_1189_, _1188_, _1181_);
  nand (_1190_, \xm8051_golden_model_1.aes_len [6], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [6]);
  or (_1191_, \xm8051_golden_model_1.aes_len [6], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [6]);
  and (_1192_, _1191_, _1190_);
  or (_1193_, \xm8051_golden_model_1.aes_len [7], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [7]);
  nand (_1194_, \xm8051_golden_model_1.aes_len [7], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [7]);
  and (_1195_, _1194_, _1193_);
  or (_1196_, _1195_, _1192_);
  and (_1197_, _1351_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [4]);
  and (_1199_, \xm8051_golden_model_1.aes_len [4], _1860_);
  or (_1200_, _1199_, _1197_);
  and (_1202_, _0517_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [5]);
  and (_1204_, \xm8051_golden_model_1.aes_len [5], _1869_);
  or (_1206_, _1204_, _1202_);
  or (_1207_, _1206_, _1200_);
  or (_1208_, _1207_, _1196_);
  or (_1209_, _1208_, _1189_);
  and (_1211_, _1828_, \xm8051_golden_model_1.aes_len [9]);
  and (_1213_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [9], _0856_);
  or (_1214_, _1213_, _1211_);
  and (_1216_, _0484_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [8]);
  and (_1217_, \xm8051_golden_model_1.aes_len [8], _0947_);
  or (_1218_, _1217_, _1216_);
  or (_1220_, _1218_, _1214_);
  and (_1221_, _0100_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [10]);
  and (_1223_, \xm8051_golden_model_1.aes_len [10], _0452_);
  or (_1224_, _1223_, _1221_);
  nand (_1226_, \xm8051_golden_model_1.aes_len [11], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [11]);
  or (_1227_, \xm8051_golden_model_1.aes_len [11], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [11]);
  and (_1228_, _1227_, _1226_);
  or (_1229_, _1228_, _1224_);
  or (_1230_, _1229_, _1220_);
  and (_1232_, _0350_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [13]);
  and (_1233_, \xm8051_golden_model_1.aes_len [13], _1354_);
  or (_1234_, _1233_, _1232_);
  and (_1235_, _1790_, \xm8051_golden_model_1.aes_len [12]);
  and (_1236_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [12], _1365_);
  or (_1237_, _1236_, _1235_);
  or (_1238_, _1237_, _1234_);
  nand (_1239_, \xm8051_golden_model_1.aes_len [15], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [15]);
  or (_1240_, \xm8051_golden_model_1.aes_len [15], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [15]);
  and (_1241_, _1240_, _1239_);
  and (_1242_, \xm8051_golden_model_1.aes_len [14], _0631_);
  and (_1243_, _0365_, \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [14]);
  or (_1244_, _1243_, _1242_);
  or (_1245_, _1244_, _1241_);
  or (_1246_, _1245_, _1238_);
  or (_1247_, _1246_, _1230_);
  or (_1248_, _1247_, _1209_);
  and (property_invalid_aes_len, _1248_, _1174_);
  and (_0000_, proc_stb, _1330_);
  or (_0001_, _1174_, rst);
  and (_1250_, _1349_, proc_data_in[0]);
  and (_1251_, _0700_, \xm8051_golden_model_1.aes_len [0]);
  or (_1252_, _1251_, _1250_);
  and (_1893_[0], _1252_, _1330_);
  dff (proc_stb_valid, _0001_);
  dff (proc_stb_r, _0000_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [0], _0542_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [1], _1225_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [0], _1256_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [1], _0880_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [2], _0835_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [3], _0701_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [4], _1137_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [5], _1834_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [6], _1134_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [7], _1837_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [8], _0821_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [9], _0318_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [10], _1551_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [11], _1269_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [12], _1001_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [13], _0279_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [14], _1554_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.operated_bytes_count [15], _0652_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.byte_counter [0], _1267_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.byte_counter [1], _1231_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.byte_counter [2], _1709_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.byte_counter [3], _1161_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [0], _0618_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [1], _1500_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [2], _1588_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [3], _1656_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [4], _0711_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [5], _0506_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [6], _0798_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [7], _1268_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [8], _1118_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [9], _1004_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [10], _0680_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [11], _1149_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [12], _0979_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [13], _0508_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [14], _0723_);
  dff (\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [15], _1667_);
  dff (\oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbit_holder [0], _0120_);
  dff (\oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbit_holder [1], _0064_);
  dff (\oc8051_xiommu_impl_1.oc8051_memarbiter_i.arbiter_state , _0062_);
  dff (\oc8051_xiommu_impl_1.oc8051_xram_i.cnt [0], _0409_);
  dff (\oc8051_xiommu_impl_1.oc8051_xram_i.cnt [1], _1006_);
  dff (\oc8051_xiommu_impl_1.oc8051_xram_i.cnt [2], _1254_);
  dff (\oc8051_xiommu_impl_1.oc8051_xram_i.ackr , _1703_);
  dff (\oc8051_xiommu_impl_1.oc8051_xram_i.ackw , _1497_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [0], _1684_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [1], _0375_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [2], _1266_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [3], _1265_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [4], _1264_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [5], _1263_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [6], _1262_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [7], _1261_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [8], _1260_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [9], _1259_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [10], _1258_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [11], _1255_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [12], _1253_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [13], _1249_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [14], _1215_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.reg_bytes_read [15], _0573_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0], _1212_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [1], _0182_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.byte_counter [0], _1210_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.byte_counter [1], _1205_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.byte_counter [2], _1203_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.byte_counter [3], _1201_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.byte_counter [4], _0553_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.byte_counter [5], _1198_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [0], _0331_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [1], _0343_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [2], _1257_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [3], _0442_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [4], _0564_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [5], _1222_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [6], _1139_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [7], _1219_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [8], _0908_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [9], _1014_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [10], _1077_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [11], _1072_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [12], _1023_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [13], _1092_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [14], _0920_);
  dff (\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [15], _1010_);
  dff (\xm8051_golden_model_1.sha_bytes_processed [0], _1895_[0]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [1], _1895_[1]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [2], _1895_[2]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [3], _1895_[3]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [4], _1895_[4]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [5], _1895_[5]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [6], _1895_[6]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [7], _1895_[7]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [8], _1895_[8]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [9], _1895_[9]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [10], _1895_[10]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [11], _1895_[11]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [12], _1895_[12]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [13], _1895_[13]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [14], _1895_[14]);
  dff (\xm8051_golden_model_1.sha_bytes_processed [15], _1895_[15]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [0], _1892_[0]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [1], _1892_[1]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [2], _1892_[2]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [3], _1892_[3]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [4], _1892_[4]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [5], _1892_[5]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [6], _1892_[6]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [7], _1892_[7]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [8], _1892_[8]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [9], _1892_[9]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [10], _1892_[10]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [11], _1892_[11]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [12], _1892_[12]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [13], _1892_[13]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [14], _1892_[14]);
  dff (\xm8051_golden_model_1.aes_bytes_processed [15], _1892_[15]);
  dff (\xm8051_golden_model_1.sha_len [0], _1896_[0]);
  dff (\xm8051_golden_model_1.sha_len [1], _1896_[1]);
  dff (\xm8051_golden_model_1.sha_len [2], _1896_[2]);
  dff (\xm8051_golden_model_1.sha_len [3], _1896_[3]);
  dff (\xm8051_golden_model_1.sha_len [4], _1896_[4]);
  dff (\xm8051_golden_model_1.sha_len [5], _1896_[5]);
  dff (\xm8051_golden_model_1.sha_len [6], _1896_[6]);
  dff (\xm8051_golden_model_1.sha_len [7], _1896_[7]);
  dff (\xm8051_golden_model_1.sha_len [8], _1896_[8]);
  dff (\xm8051_golden_model_1.sha_len [9], _1896_[9]);
  dff (\xm8051_golden_model_1.sha_len [10], _1896_[10]);
  dff (\xm8051_golden_model_1.sha_len [11], _1896_[11]);
  dff (\xm8051_golden_model_1.sha_len [12], _1896_[12]);
  dff (\xm8051_golden_model_1.sha_len [13], _1896_[13]);
  dff (\xm8051_golden_model_1.sha_len [14], _1896_[14]);
  dff (\xm8051_golden_model_1.sha_len [15], _1896_[15]);
  dff (\xm8051_golden_model_1.aes_len [0], _1893_[0]);
  dff (\xm8051_golden_model_1.aes_len [1], _1893_[1]);
  dff (\xm8051_golden_model_1.aes_len [2], _1893_[2]);
  dff (\xm8051_golden_model_1.aes_len [3], _1893_[3]);
  dff (\xm8051_golden_model_1.aes_len [4], _1893_[4]);
  dff (\xm8051_golden_model_1.aes_len [5], _1893_[5]);
  dff (\xm8051_golden_model_1.aes_len [6], _1893_[6]);
  dff (\xm8051_golden_model_1.aes_len [7], _1893_[7]);
  dff (\xm8051_golden_model_1.aes_len [8], _1893_[8]);
  dff (\xm8051_golden_model_1.aes_len [9], _1893_[9]);
  dff (\xm8051_golden_model_1.aes_len [10], _1893_[10]);
  dff (\xm8051_golden_model_1.aes_len [11], _1893_[11]);
  dff (\xm8051_golden_model_1.aes_len [12], _1893_[12]);
  dff (\xm8051_golden_model_1.aes_len [13], _1893_[13]);
  dff (\xm8051_golden_model_1.aes_len [14], _1893_[14]);
  dff (\xm8051_golden_model_1.aes_len [15], _1893_[15]);
  dff (\xm8051_golden_model_1.sha_state [0], _1897_[0]);
  dff (\xm8051_golden_model_1.sha_state [1], _1897_[1]);
  dff (\xm8051_golden_model_1.sha_state [2], 1'b0);
  dff (\xm8051_golden_model_1.sha_state [3], 1'b0);
  dff (\xm8051_golden_model_1.sha_state [4], 1'b0);
  dff (\xm8051_golden_model_1.sha_state [5], 1'b0);
  dff (\xm8051_golden_model_1.sha_state [6], 1'b0);
  dff (\xm8051_golden_model_1.sha_state [7], 1'b0);
  dff (\xm8051_golden_model_1.aes_state [0], _1894_[0]);
  dff (\xm8051_golden_model_1.aes_state [1], _1894_[1]);
  dff (\xm8051_golden_model_1.aes_state [2], 1'b0);
  dff (\xm8051_golden_model_1.aes_state [3], 1'b0);
  dff (\xm8051_golden_model_1.aes_state [4], 1'b0);
  dff (\xm8051_golden_model_1.aes_state [5], 1'b0);
  dff (\xm8051_golden_model_1.aes_state [6], 1'b0);
  dff (\xm8051_golden_model_1.aes_state [7], 1'b0);
  buf(\xm8051_golden_model_1.n0881 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0881 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0881 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0881 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0881 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0881 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0881 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0881 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0881 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0881 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0881 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0881 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0881 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0881 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0881 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0881 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0881 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0881 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0881 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0881 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0881 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0881 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0881 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0881 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0881 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0881 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0881 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0881 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0881 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0881 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0881 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0881 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0881 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0881 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0881 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0881 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0881 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0881 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0881 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0881 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0881 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0881 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0881 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0881 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0881 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0881 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0881 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0881 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0881 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0881 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0881 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0881 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0881 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0881 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0881 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0881 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0881 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0881 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0881 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0881 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0881 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0881 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0881 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0881 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0881 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0881 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0881 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0881 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0881 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0881 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0881 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0881 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0881 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0881 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0881 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0881 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0881 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0881 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0881 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0881 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0881 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0881 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0881 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0881 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0881 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0881 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0881 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0881 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0881 [88], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0881 [89], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0881 [90], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0881 [91], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0881 [92], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0881 [93], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0881 [94], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0881 [95], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0881 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0881 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0881 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0881 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0881 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0881 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0881 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0881 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0881 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0881 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0881 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0881 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0881 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0881 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0881 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0881 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0881 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0881 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0881 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0881 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0881 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0881 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0881 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0881 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0881 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0881 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0881 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0881 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0881 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0881 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0881 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0881 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0880 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0880 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0880 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0880 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0880 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0880 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0880 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0880 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0880 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0880 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0880 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0880 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0880 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0880 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0880 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0880 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0880 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0880 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0880 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0880 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0880 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0880 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0880 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0880 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0880 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0880 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0880 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0880 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0880 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0880 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0880 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0880 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0880 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0880 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0880 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0880 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0880 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0880 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0880 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0880 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0880 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0880 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0880 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0880 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0880 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0880 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0880 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0880 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0880 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0880 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0880 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0880 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0880 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0880 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0880 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0880 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0880 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0880 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0880 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0880 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0880 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0880 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0880 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0880 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0880 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0880 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0880 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0880 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0880 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0880 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0880 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0880 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0880 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0880 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0880 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0880 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0880 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0880 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0880 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0880 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0880 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0880 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0880 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0880 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0880 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0880 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0880 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0880 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0453 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0453 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0453 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n0879 [0], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0879 [1], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0879 [2], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0879 [3], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0879 [4], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0879 [5], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0879 [6], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0879 [7], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0879 [8], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0879 [9], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0879 [10], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0879 [11], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0879 [12], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0879 [13], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0879 [14], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0879 [15], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0879 [16], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0879 [17], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0879 [18], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0879 [19], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0879 [20], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0879 [21], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0879 [22], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0879 [23], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0879 [24], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0879 [25], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0879 [26], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0879 [27], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0879 [28], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0879 [29], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0879 [30], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0879 [31], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0878 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0878 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0878 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0878 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0878 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0878 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0878 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0878 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0878 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0878 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0878 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0878 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0878 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0878 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0878 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0878 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0878 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0878 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0878 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0878 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0878 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0878 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0878 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0878 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0878 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0878 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0878 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0878 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0878 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0878 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0878 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0878 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0878 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0878 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0878 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0878 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0878 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0878 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0878 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0878 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0878 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0878 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0878 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0878 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0878 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0878 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0878 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0878 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0878 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0878 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0878 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0878 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0878 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0878 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0878 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0878 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0878 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0878 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0878 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0878 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0878 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0878 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0878 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0878 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0878 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0878 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0878 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0878 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0878 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0878 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0878 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0878 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0878 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0878 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0878 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0878 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0878 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0878 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0878 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0878 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0878 [80], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0878 [81], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0878 [82], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0878 [83], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0878 [84], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0878 [85], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0878 [86], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0878 [87], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0878 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0878 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0878 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0878 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0878 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0878 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0878 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0878 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0878 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0878 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0878 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0878 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0878 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0878 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0878 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0878 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0878 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0878 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0878 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0878 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0878 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0878 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0878 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0878 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0878 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0878 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0878 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0878 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0878 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0878 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0878 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0878 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0878 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0878 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0878 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0878 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0878 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0878 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0878 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0878 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0877 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0877 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0877 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0877 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0877 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0877 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0877 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0877 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0877 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0877 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0877 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0877 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0877 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0877 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0877 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0877 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0877 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0877 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0877 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0877 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0877 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0877 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0877 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0877 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0877 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0877 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0877 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0877 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0877 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0877 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0877 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0877 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0877 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0877 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0877 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0877 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0877 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0877 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0877 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0877 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0877 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0877 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0877 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0877 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0877 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0877 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0877 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0877 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0877 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0877 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0877 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0877 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0877 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0877 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0877 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0877 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0877 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0877 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0877 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0877 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0877 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0877 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0877 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0877 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0877 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0877 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0877 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0877 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0877 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0877 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0877 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0877 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0877 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0877 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0877 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0877 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0877 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0877 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0877 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0877 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0876 [0], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0876 [1], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0876 [2], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0876 [3], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0876 [4], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0876 [5], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0876 [6], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0876 [7], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0876 [8], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0876 [9], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0876 [10], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0876 [11], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0876 [12], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0876 [13], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0876 [14], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0876 [15], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0876 [16], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0876 [17], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0876 [18], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0876 [19], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0876 [20], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0876 [21], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0876 [22], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0876 [23], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0876 [24], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0876 [25], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0876 [26], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0876 [27], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0876 [28], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0876 [29], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0876 [30], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0876 [31], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0876 [32], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0876 [33], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0876 [34], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0876 [35], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0876 [36], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0876 [37], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0876 [38], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0876 [39], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0875 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0875 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0875 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0875 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0875 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0875 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0875 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0875 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0875 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0875 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0875 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0875 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0875 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0875 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0875 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0875 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0875 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0875 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0875 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0875 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0875 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0875 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0875 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0875 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0875 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0875 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0875 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0875 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0875 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0875 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0875 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0875 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0875 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0875 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0875 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0875 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0875 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0875 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0875 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0875 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0875 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0875 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0875 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0875 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0875 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0875 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0875 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0875 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0875 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0875 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0875 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0875 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0875 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0875 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0875 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0875 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0875 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0875 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0875 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0875 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0875 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0875 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0875 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0875 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0875 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0875 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0875 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0875 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0875 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0875 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0875 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0875 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0875 [72], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0875 [73], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0875 [74], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0875 [75], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0875 [76], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0875 [77], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0875 [78], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0875 [79], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0875 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0875 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0875 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0875 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0875 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0875 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0875 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0875 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0875 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0875 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0875 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0875 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0875 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0875 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0875 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0875 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0875 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0875 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0875 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0875 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0875 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0875 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0875 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0875 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0875 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0875 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0875 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0875 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0875 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0875 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0875 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0875 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0875 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0875 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0875 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0875 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0875 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0875 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0875 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0875 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0875 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0875 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0875 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0875 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0875 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0875 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0875 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0875 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0874 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0874 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0874 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0874 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0874 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0874 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0874 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0874 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0874 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0874 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0874 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0874 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0874 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0874 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0874 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0874 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0874 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0874 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0874 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0874 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0874 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0874 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0874 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0874 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0874 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0874 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0874 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0874 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0874 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0874 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0874 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0874 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0874 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0874 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0874 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0874 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0874 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0874 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0874 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0874 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0874 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0874 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0874 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0874 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0874 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0874 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0874 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0874 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0874 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0874 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0874 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0874 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0874 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0874 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0874 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0874 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0874 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0874 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0874 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0874 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0874 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0874 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0874 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0874 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0874 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0874 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0874 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0874 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0874 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0874 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0874 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0874 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0873 [0], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0873 [1], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0873 [2], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0873 [3], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0873 [4], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0873 [5], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0873 [6], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0873 [7], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0873 [8], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0873 [9], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0873 [10], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0873 [11], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0873 [12], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0873 [13], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0873 [14], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0873 [15], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0873 [16], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0873 [17], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0873 [18], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0873 [19], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0873 [20], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0873 [21], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0873 [22], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0873 [23], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0873 [24], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0873 [25], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0873 [26], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0873 [27], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0873 [28], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0873 [29], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0873 [30], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0873 [31], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0873 [32], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0873 [33], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0873 [34], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0873 [35], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0873 [36], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0873 [37], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0873 [38], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0873 [39], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0873 [40], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0873 [41], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0873 [42], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0873 [43], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0873 [44], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0873 [45], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0873 [46], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0873 [47], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0872 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0872 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0872 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0872 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0872 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0872 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0872 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0872 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0872 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0872 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0872 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0872 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0872 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0872 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0872 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0872 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0872 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0872 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0872 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0872 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0872 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0872 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0872 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0872 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0872 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0872 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0872 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0872 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0872 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0872 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0872 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0872 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0872 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0872 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0872 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0872 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0872 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0872 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0872 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0872 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0872 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0872 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0872 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0872 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0872 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0872 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0872 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0872 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0872 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0872 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0872 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0872 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0872 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0872 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0872 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0872 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0872 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0872 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0872 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0872 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0872 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0872 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0872 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0872 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0872 [64], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0872 [65], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0872 [66], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0872 [67], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0872 [68], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0872 [69], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0872 [70], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0872 [71], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0872 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0872 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0872 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0872 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0872 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0872 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0872 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0872 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0872 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0872 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0872 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0872 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0872 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0872 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0872 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0872 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0872 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0872 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0872 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0872 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0872 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0872 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0872 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0872 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0872 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0872 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0872 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0872 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0872 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0872 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0872 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0872 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0872 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0872 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0872 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0872 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0872 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0872 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0872 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0872 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0872 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0872 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0872 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0872 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0872 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0872 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0872 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0872 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0872 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0872 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0872 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0872 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0872 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0872 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0872 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0872 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0871 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0871 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0871 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0871 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0871 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0871 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0871 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0871 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0871 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0871 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0871 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0871 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0871 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0871 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0871 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0871 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0871 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0871 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0871 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0871 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0871 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0871 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0871 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0871 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0871 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0871 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0871 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0871 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0871 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0871 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0871 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0871 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0871 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0871 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0871 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0871 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0871 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0871 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0871 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0871 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0871 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0871 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0871 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0871 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0871 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0871 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0871 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0871 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0871 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0871 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0871 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0871 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0871 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0871 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0871 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0871 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0871 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0871 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0871 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0871 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0871 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0871 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0871 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0871 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0e [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.n0443 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0443 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0443 [2], \xm8051_golden_model_1.n0483 [2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0c [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.n0870 [0], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0870 [1], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0870 [2], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0870 [3], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0870 [4], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0870 [5], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0870 [6], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0870 [7], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0870 [8], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0870 [9], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0870 [10], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0870 [11], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0870 [12], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0870 [13], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0870 [14], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0870 [15], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0870 [16], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0870 [17], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0870 [18], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0870 [19], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0870 [20], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0870 [21], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0870 [22], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0870 [23], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0870 [24], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0870 [25], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0870 [26], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0870 [27], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0870 [28], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0870 [29], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0870 [30], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0870 [31], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0870 [32], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0870 [33], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0870 [34], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0870 [35], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0870 [36], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0870 [37], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0870 [38], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0870 [39], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0870 [40], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0870 [41], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0870 [42], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0870 [43], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0870 [44], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0870 [45], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0870 [46], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0870 [47], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0870 [48], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0870 [49], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0870 [50], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0870 [51], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0870 [52], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0870 [53], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0870 [54], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0870 [55], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_0a [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_09 [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_08 [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.n0869 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0869 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0869 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0869 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0869 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0869 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0869 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0869 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0869 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0869 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0869 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0869 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0869 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0869 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0869 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0869 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0869 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0869 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0869 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0869 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0869 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0869 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0869 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0869 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0869 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0869 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0869 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0869 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0869 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0869 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0869 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0869 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0869 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0869 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0869 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0869 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0869 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0869 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0869 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0869 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0869 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0869 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0869 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0869 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0869 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0869 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0869 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0869 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0869 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0869 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0869 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0869 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0869 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0869 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0869 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0869 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0869 [56], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0869 [57], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0869 [58], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0869 [59], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0869 [60], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0869 [61], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0869 [62], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0869 [63], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0869 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0869 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0869 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0869 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0869 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0869 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0869 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0869 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0869 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0869 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0869 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0869 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0869 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0869 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0869 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0869 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0869 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0869 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0869 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0869 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0869 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0869 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0869 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0869 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0869 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0869 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0869 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0869 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0869 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0869 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0869 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0869 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0869 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0869 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0869 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0869 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0869 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0869 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0869 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0869 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0869 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0869 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0869 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0869 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0869 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0869 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0869 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0869 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0869 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0869 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0869 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0869 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0869 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0869 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0869 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0869 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0869 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0869 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0869 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0869 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0869 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0869 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0869 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0869 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_06 [15], proc_addr[15]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.data_in_A [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.data_in_A [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.data_in_A [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.data_in_A [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.data_in_A [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.data_in_A [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.data_in_A [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.data_in_A [7], proc_data_in[7]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [0], proc_addr[0]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [1], proc_addr[1]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [2], proc_addr[2]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [3], proc_addr[3]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [4], proc_addr[4]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [5], proc_addr[5]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [6], proc_addr[6]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [7], proc_addr[7]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [8], proc_addr[8]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [9], proc_addr[9]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [10], proc_addr[10]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [11], proc_addr[11]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [12], proc_addr[12]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [13], proc_addr[13]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [14], proc_addr[14]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.addr_A [15], proc_addr[15]);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.rst , rst);
  buf(\oc8051_xiommu_impl_1.oc8051_memarbiter_i.clk , clk);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [0], ABINPUT[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [1], ABINPUT[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [2], ABINPUT[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [3], ABINPUT[3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [4], ABINPUT[4]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [5], ABINPUT[5]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [6], ABINPUT[6]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [7], ABINPUT[7]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [8], ABINPUT[8]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [9], ABINPUT[9]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [10], ABINPUT[10]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [11], ABINPUT[11]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [12], ABINPUT[12]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [13], ABINPUT[13]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [14], ABINPUT[14]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [15], ABINPUT[15]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [16], ABINPUT[16]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [17], ABINPUT[17]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [18], ABINPUT[18]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [19], ABINPUT[19]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [20], ABINPUT[20]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [21], ABINPUT[21]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [22], ABINPUT[22]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [23], ABINPUT[23]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [24], ABINPUT[24]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [25], ABINPUT[25]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [26], ABINPUT[26]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [27], ABINPUT[27]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [28], ABINPUT[28]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [29], ABINPUT[29]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [30], ABINPUT[30]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [31], ABINPUT[31]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [32], ABINPUT[32]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [33], ABINPUT[33]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [34], ABINPUT[34]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [35], ABINPUT[35]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [36], ABINPUT[36]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [37], ABINPUT[37]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [38], ABINPUT[38]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [39], ABINPUT[39]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [40], ABINPUT[40]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [41], ABINPUT[41]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [42], ABINPUT[42]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [43], ABINPUT[43]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [44], ABINPUT[44]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [45], ABINPUT[45]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [46], ABINPUT[46]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [47], ABINPUT[47]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [48], ABINPUT[48]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [49], ABINPUT[49]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [50], ABINPUT[50]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [51], ABINPUT[51]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [52], ABINPUT[52]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [53], ABINPUT[53]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [54], ABINPUT[54]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [55], ABINPUT[55]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [56], ABINPUT[56]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [57], ABINPUT[57]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [58], ABINPUT[58]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [59], ABINPUT[59]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [60], ABINPUT[60]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [61], ABINPUT[61]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [62], ABINPUT[62]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [63], ABINPUT[63]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [64], ABINPUT[64]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [65], ABINPUT[65]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [66], ABINPUT[66]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [67], ABINPUT[67]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [68], ABINPUT[68]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [69], ABINPUT[69]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [70], ABINPUT[70]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [71], ABINPUT[71]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [72], ABINPUT[72]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [73], ABINPUT[73]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [74], ABINPUT[74]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [75], ABINPUT[75]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [76], ABINPUT[76]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [77], ABINPUT[77]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [78], ABINPUT[78]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [79], ABINPUT[79]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [80], ABINPUT[80]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [81], ABINPUT[81]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [82], ABINPUT[82]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [83], ABINPUT[83]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [84], ABINPUT[84]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [85], ABINPUT[85]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [86], ABINPUT[86]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [87], ABINPUT[87]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [88], ABINPUT[88]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [89], ABINPUT[89]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [90], ABINPUT[90]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [91], ABINPUT[91]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [92], ABINPUT[92]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [93], ABINPUT[93]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [94], ABINPUT[94]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [95], ABINPUT[95]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [96], ABINPUT[96]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [97], ABINPUT[97]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [98], ABINPUT[98]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [99], ABINPUT[99]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [100], ABINPUT[100]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [101], ABINPUT[101]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [102], ABINPUT[102]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [103], ABINPUT[103]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [104], ABINPUT[104]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [105], ABINPUT[105]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [106], ABINPUT[106]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [107], ABINPUT[107]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [108], ABINPUT[108]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [109], ABINPUT[109]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [110], ABINPUT[110]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [111], ABINPUT[111]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [112], ABINPUT[112]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [113], ABINPUT[113]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [114], ABINPUT[114]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [115], ABINPUT[115]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [116], ABINPUT[116]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [117], ABINPUT[117]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [118], ABINPUT[118]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [119], ABINPUT[119]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [120], ABINPUT[120]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [121], ABINPUT[121]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [122], ABINPUT[122]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [123], ABINPUT[123]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [124], ABINPUT[124]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [125], ABINPUT[125]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [126], ABINPUT[126]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_out [127], ABINPUT[127]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_05 [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_04 [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.n0868 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0868 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0868 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0868 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0868 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0868 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0868 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0868 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0868 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0868 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0868 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0868 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0868 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0868 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0868 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0868 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0868 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0868 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0868 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0868 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0868 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0868 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0868 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0868 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0868 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0868 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0868 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0868 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0868 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0868 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0868 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0868 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0868 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0868 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0868 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0868 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0868 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0868 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0868 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0868 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0868 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0868 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0868 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0868 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0868 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0868 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0868 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0868 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0868 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0868 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0868 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0868 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0868 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0868 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0868 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0868 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_02 [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_01 [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.WR_XRAM_ADDR_00 [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_119 , nondet_memwrite_choice_119);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_118 , nondet_memwrite_choice_118);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_117 , nondet_memwrite_choice_117);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_116 , nondet_memwrite_choice_116);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [0], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [1], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [2], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [3], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [4], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [4]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [5], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [5]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [6], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [6]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [7], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [7]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [8], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [8]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [9], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [9]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [10], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [10]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [11], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [11]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [12], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [12]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [13], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [13]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [14], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [14]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_len [15], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [15]);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_115 , nondet_memwrite_choice_115);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_114 , nondet_memwrite_choice_114);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_113 , nondet_memwrite_choice_113);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_112 , nondet_memwrite_choice_112);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_111 , nondet_memwrite_choice_111);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_110 , nondet_memwrite_choice_110);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_state [0], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_state [1], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [1]);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_109 , nondet_memwrite_choice_109);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_108 , nondet_memwrite_choice_108);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_107 , nondet_memwrite_choice_107);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_106 , nondet_memwrite_choice_106);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_105 , nondet_memwrite_choice_105);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_104 , nondet_memwrite_choice_104);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_103 , nondet_memwrite_choice_103);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_102 , nondet_memwrite_choice_102);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_101 , nondet_memwrite_choice_101);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_100 , nondet_memwrite_choice_100);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_99 , nondet_memwrite_choice_99);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_98 , nondet_memwrite_choice_98);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_97 , nondet_memwrite_choice_97);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_96 , nondet_memwrite_choice_96);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_95 , nondet_memwrite_choice_95);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_94 , nondet_memwrite_choice_94);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [0], proc_addr[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [1], proc_addr[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [2], proc_addr[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [3], proc_addr[3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [4], proc_addr[4]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [5], proc_addr[5]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [6], proc_addr[6]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [7], proc_addr[7]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [8], proc_addr[8]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [9], proc_addr[9]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [10], proc_addr[10]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [11], proc_addr[11]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [12], proc_addr[12]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [13], proc_addr[13]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [14], proc_addr[14]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.addr [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_93 , nondet_memwrite_choice_93);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_92 , nondet_memwrite_choice_92);
  buf(\oc8051_xiommu_impl_1.aes_top_i.data_in [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.data_in [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.data_in [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.data_in [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.data_in [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.data_in [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.data_in [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.data_in [7], proc_data_in[7]);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_91 , nondet_memwrite_choice_91);
  buf(\oc8051_xiommu_impl_1.aes_top_i.rst , rst);
  buf(\oc8051_xiommu_impl_1.aes_top_i.clk , clk);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_90 , nondet_memwrite_choice_90);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [9], ABINPUT[9]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [10], ABINPUT[10]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [11], ABINPUT[11]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [12], ABINPUT[12]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [13], ABINPUT[13]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [14], ABINPUT[14]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [15], ABINPUT[15]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [16], ABINPUT[16]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [17], ABINPUT[17]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [18], ABINPUT[18]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [19], ABINPUT[19]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [20], ABINPUT[20]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [21], ABINPUT[21]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [22], ABINPUT[22]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [23], ABINPUT[23]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [24], ABINPUT[24]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [25], ABINPUT[25]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [26], ABINPUT[26]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [27], ABINPUT[27]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [28], ABINPUT[28]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [29], ABINPUT[29]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [30], ABINPUT[30]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [31], ABINPUT[31]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [32], ABINPUT[32]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [33], ABINPUT[33]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [34], ABINPUT[34]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [35], ABINPUT[35]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [36], ABINPUT[36]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [37], ABINPUT[37]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [38], ABINPUT[38]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [39], ABINPUT[39]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [40], ABINPUT[40]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [41], ABINPUT[41]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [42], ABINPUT[42]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [43], ABINPUT[43]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [44], ABINPUT[44]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [45], ABINPUT[45]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [46], ABINPUT[46]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [47], ABINPUT[47]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [48], ABINPUT[48]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [49], ABINPUT[49]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [50], ABINPUT[50]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [51], ABINPUT[51]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [52], ABINPUT[52]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [53], ABINPUT[53]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [54], ABINPUT[54]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [55], ABINPUT[55]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [56], ABINPUT[56]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [57], ABINPUT[57]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [58], ABINPUT[58]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [59], ABINPUT[59]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [60], ABINPUT[60]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [61], ABINPUT[61]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [62], ABINPUT[62]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [63], ABINPUT[63]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [64], ABINPUT[64]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [65], ABINPUT[65]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [66], ABINPUT[66]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [67], ABINPUT[67]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [68], ABINPUT[68]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [69], ABINPUT[69]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [70], ABINPUT[70]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [71], ABINPUT[71]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [72], ABINPUT[72]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [73], ABINPUT[73]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [74], ABINPUT[74]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [75], ABINPUT[75]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [76], ABINPUT[76]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [77], ABINPUT[77]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [78], ABINPUT[78]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [79], ABINPUT[79]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [80], ABINPUT[80]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [81], ABINPUT[81]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [82], ABINPUT[82]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [83], ABINPUT[83]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [84], ABINPUT[84]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [85], ABINPUT[85]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [86], ABINPUT[86]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [87], ABINPUT[87]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [88], ABINPUT[88]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [89], ABINPUT[89]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [90], ABINPUT[90]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [91], ABINPUT[91]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [92], ABINPUT[92]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [93], ABINPUT[93]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [94], ABINPUT[94]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [95], ABINPUT[95]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [96], ABINPUT[96]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [97], ABINPUT[97]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [98], ABINPUT[98]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [99], ABINPUT[99]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [100], ABINPUT[100]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [101], ABINPUT[101]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [102], ABINPUT[102]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [103], ABINPUT[103]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [104], ABINPUT[104]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [105], ABINPUT[105]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [106], ABINPUT[106]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [107], ABINPUT[107]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [108], ABINPUT[108]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [109], ABINPUT[109]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [110], ABINPUT[110]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [111], ABINPUT[111]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [112], ABINPUT[112]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [113], ABINPUT[113]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [114], ABINPUT[114]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [115], ABINPUT[115]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [116], ABINPUT[116]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [117], ABINPUT[117]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [118], ABINPUT[118]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [119], ABINPUT[119]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [120], ABINPUT[120]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [121], ABINPUT[121]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [122], ABINPUT[122]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [123], ABINPUT[123]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [124], ABINPUT[124]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [125], ABINPUT[125]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [126], ABINPUT[126]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.ABINPUT [127], ABINPUT[127]);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_89 , nondet_memwrite_choice_89);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_88 , nondet_memwrite_choice_88);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_87 , nondet_memwrite_choice_87);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_86 , nondet_memwrite_choice_86);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_85 , nondet_memwrite_choice_85);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_84 , nondet_memwrite_choice_84);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_83 , nondet_memwrite_choice_83);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_82 , nondet_memwrite_choice_82);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_81 , nondet_memwrite_choice_81);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_80 , nondet_memwrite_choice_80);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_79 , nondet_memwrite_choice_79);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_78 , nondet_memwrite_choice_78);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_77 , nondet_memwrite_choice_77);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_76 , nondet_memwrite_choice_76);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_75 , nondet_memwrite_choice_75);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_74 , nondet_memwrite_choice_74);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_73 , nondet_memwrite_choice_73);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_72 , nondet_memwrite_choice_72);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_71 , nondet_memwrite_choice_71);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_70 , nondet_memwrite_choice_70);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_69 , nondet_memwrite_choice_69);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_68 , nondet_memwrite_choice_68);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_67 , nondet_memwrite_choice_67);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_66 , nondet_memwrite_choice_66);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_65 , nondet_memwrite_choice_65);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_64 , nondet_memwrite_choice_64);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_63 , nondet_memwrite_choice_63);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_62 , nondet_memwrite_choice_62);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_61 , nondet_memwrite_choice_61);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_60 , nondet_memwrite_choice_60);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_59 , nondet_memwrite_choice_59);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [0], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [1], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [2], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [3], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [4], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [4]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [5], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [5]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [6], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [6]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [7], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [7]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [8], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [8]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [9], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [9]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [10], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [10]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [11], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [11]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [12], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [12]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [13], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [13]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [14], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [14]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen [15], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [15]);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_58 , nondet_memwrite_choice_58);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_57 , nondet_memwrite_choice_57);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_56 , nondet_memwrite_choice_56);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_55 , nondet_memwrite_choice_55);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_54 , nondet_memwrite_choice_54);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_53 , nondet_memwrite_choice_53);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_52 , nondet_memwrite_choice_52);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_51 , nondet_memwrite_choice_51);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_50 , nondet_memwrite_choice_50);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_49 , nondet_memwrite_choice_49);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_48 , nondet_memwrite_choice_48);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_47 , nondet_memwrite_choice_47);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_46 , nondet_memwrite_choice_46);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_45 , nondet_memwrite_choice_45);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_44 , nondet_memwrite_choice_44);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_43 , nondet_memwrite_choice_43);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_42 , nondet_memwrite_choice_42);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_41 , nondet_memwrite_choice_41);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_40 , nondet_memwrite_choice_40);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_39 , nondet_memwrite_choice_39);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_38 , nondet_memwrite_choice_38);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_37 , nondet_memwrite_choice_37);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_36 , nondet_memwrite_choice_36);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_35 , nondet_memwrite_choice_35);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_34 , nondet_memwrite_choice_34);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_33 , nondet_memwrite_choice_33);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_32 , nondet_memwrite_choice_32);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_31 , nondet_memwrite_choice_31);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_30 , nondet_memwrite_choice_30);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_29 , nondet_memwrite_choice_29);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_28 , nondet_memwrite_choice_28);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_27 , nondet_memwrite_choice_27);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_26 , nondet_memwrite_choice_26);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_25 , nondet_memwrite_choice_25);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_24 , nondet_memwrite_choice_24);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_23 , nondet_memwrite_choice_23);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_22 , nondet_memwrite_choice_22);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_21 , nondet_memwrite_choice_21);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_20 , nondet_memwrite_choice_20);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_19 , nondet_memwrite_choice_19);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_18 , nondet_memwrite_choice_18);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_17 , nondet_memwrite_choice_17);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_16 , nondet_memwrite_choice_16);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_15 , nondet_memwrite_choice_15);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_14 , nondet_memwrite_choice_14);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_13 , nondet_memwrite_choice_13);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_12 , nondet_memwrite_choice_12);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_11 , nondet_memwrite_choice_11);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_10 , nondet_memwrite_choice_10);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_9 , nondet_memwrite_choice_9);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_8 , nondet_memwrite_choice_8);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_7 , nondet_memwrite_choice_7);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_6 , nondet_memwrite_choice_6);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_5 , nondet_memwrite_choice_5);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_4 , nondet_memwrite_choice_4);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_3 , nondet_memwrite_choice_3);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_2 , nondet_memwrite_choice_2);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_1 , nondet_memwrite_choice_1);
  buf(\xm8051_golden_model_1.nondet_memwrite_choice_0 , nondet_memwrite_choice_0);
  buf(\xm8051_golden_model_1.RD_xram_80 [0], RD_xram_80[0]);
  buf(\xm8051_golden_model_1.RD_xram_80 [1], RD_xram_80[1]);
  buf(\xm8051_golden_model_1.RD_xram_80 [2], RD_xram_80[2]);
  buf(\xm8051_golden_model_1.RD_xram_80 [3], RD_xram_80[3]);
  buf(\xm8051_golden_model_1.RD_xram_80 [4], RD_xram_80[4]);
  buf(\xm8051_golden_model_1.RD_xram_80 [5], RD_xram_80[5]);
  buf(\xm8051_golden_model_1.RD_xram_80 [6], RD_xram_80[6]);
  buf(\xm8051_golden_model_1.RD_xram_80 [7], RD_xram_80[7]);
  buf(\xm8051_golden_model_1.RD_xram_79 [0], RD_xram_79[0]);
  buf(\xm8051_golden_model_1.RD_xram_79 [1], RD_xram_79[1]);
  buf(\xm8051_golden_model_1.RD_xram_79 [2], RD_xram_79[2]);
  buf(\xm8051_golden_model_1.RD_xram_79 [3], RD_xram_79[3]);
  buf(\xm8051_golden_model_1.RD_xram_79 [4], RD_xram_79[4]);
  buf(\xm8051_golden_model_1.RD_xram_79 [5], RD_xram_79[5]);
  buf(\xm8051_golden_model_1.RD_xram_79 [6], RD_xram_79[6]);
  buf(\xm8051_golden_model_1.RD_xram_79 [7], RD_xram_79[7]);
  buf(\xm8051_golden_model_1.RD_xram_78 [0], RD_xram_78[0]);
  buf(\xm8051_golden_model_1.RD_xram_78 [1], RD_xram_78[1]);
  buf(\xm8051_golden_model_1.RD_xram_78 [2], RD_xram_78[2]);
  buf(\xm8051_golden_model_1.RD_xram_78 [3], RD_xram_78[3]);
  buf(\xm8051_golden_model_1.RD_xram_78 [4], RD_xram_78[4]);
  buf(\xm8051_golden_model_1.RD_xram_78 [5], RD_xram_78[5]);
  buf(\xm8051_golden_model_1.RD_xram_78 [6], RD_xram_78[6]);
  buf(\xm8051_golden_model_1.RD_xram_78 [7], RD_xram_78[7]);
  buf(\xm8051_golden_model_1.RD_xram_77 [0], RD_xram_77[0]);
  buf(\xm8051_golden_model_1.RD_xram_77 [1], RD_xram_77[1]);
  buf(\xm8051_golden_model_1.RD_xram_77 [2], RD_xram_77[2]);
  buf(\xm8051_golden_model_1.RD_xram_77 [3], RD_xram_77[3]);
  buf(\xm8051_golden_model_1.RD_xram_77 [4], RD_xram_77[4]);
  buf(\xm8051_golden_model_1.RD_xram_77 [5], RD_xram_77[5]);
  buf(\xm8051_golden_model_1.RD_xram_77 [6], RD_xram_77[6]);
  buf(\xm8051_golden_model_1.RD_xram_77 [7], RD_xram_77[7]);
  buf(\xm8051_golden_model_1.RD_xram_76 [0], RD_xram_76[0]);
  buf(\xm8051_golden_model_1.RD_xram_76 [1], RD_xram_76[1]);
  buf(\xm8051_golden_model_1.RD_xram_76 [2], RD_xram_76[2]);
  buf(\xm8051_golden_model_1.RD_xram_76 [3], RD_xram_76[3]);
  buf(\xm8051_golden_model_1.RD_xram_76 [4], RD_xram_76[4]);
  buf(\xm8051_golden_model_1.RD_xram_76 [5], RD_xram_76[5]);
  buf(\xm8051_golden_model_1.RD_xram_76 [6], RD_xram_76[6]);
  buf(\xm8051_golden_model_1.RD_xram_76 [7], RD_xram_76[7]);
  buf(\xm8051_golden_model_1.RD_xram_75 [0], RD_xram_75[0]);
  buf(\xm8051_golden_model_1.RD_xram_75 [1], RD_xram_75[1]);
  buf(\xm8051_golden_model_1.RD_xram_75 [2], RD_xram_75[2]);
  buf(\xm8051_golden_model_1.RD_xram_75 [3], RD_xram_75[3]);
  buf(\xm8051_golden_model_1.RD_xram_75 [4], RD_xram_75[4]);
  buf(\xm8051_golden_model_1.RD_xram_75 [5], RD_xram_75[5]);
  buf(\xm8051_golden_model_1.RD_xram_75 [6], RD_xram_75[6]);
  buf(\xm8051_golden_model_1.RD_xram_75 [7], RD_xram_75[7]);
  buf(\xm8051_golden_model_1.RD_xram_74 [0], RD_xram_74[0]);
  buf(\xm8051_golden_model_1.RD_xram_74 [1], RD_xram_74[1]);
  buf(\xm8051_golden_model_1.RD_xram_74 [2], RD_xram_74[2]);
  buf(\xm8051_golden_model_1.RD_xram_74 [3], RD_xram_74[3]);
  buf(\xm8051_golden_model_1.RD_xram_74 [4], RD_xram_74[4]);
  buf(\xm8051_golden_model_1.RD_xram_74 [5], RD_xram_74[5]);
  buf(\xm8051_golden_model_1.RD_xram_74 [6], RD_xram_74[6]);
  buf(\xm8051_golden_model_1.RD_xram_74 [7], RD_xram_74[7]);
  buf(\xm8051_golden_model_1.RD_xram_73 [0], RD_xram_73[0]);
  buf(\xm8051_golden_model_1.RD_xram_73 [1], RD_xram_73[1]);
  buf(\xm8051_golden_model_1.RD_xram_73 [2], RD_xram_73[2]);
  buf(\xm8051_golden_model_1.RD_xram_73 [3], RD_xram_73[3]);
  buf(\xm8051_golden_model_1.RD_xram_73 [4], RD_xram_73[4]);
  buf(\xm8051_golden_model_1.RD_xram_73 [5], RD_xram_73[5]);
  buf(\xm8051_golden_model_1.RD_xram_73 [6], RD_xram_73[6]);
  buf(\xm8051_golden_model_1.RD_xram_73 [7], RD_xram_73[7]);
  buf(\xm8051_golden_model_1.RD_xram_72 [0], RD_xram_72[0]);
  buf(\xm8051_golden_model_1.RD_xram_72 [1], RD_xram_72[1]);
  buf(\xm8051_golden_model_1.RD_xram_72 [2], RD_xram_72[2]);
  buf(\xm8051_golden_model_1.RD_xram_72 [3], RD_xram_72[3]);
  buf(\xm8051_golden_model_1.RD_xram_72 [4], RD_xram_72[4]);
  buf(\xm8051_golden_model_1.RD_xram_72 [5], RD_xram_72[5]);
  buf(\xm8051_golden_model_1.RD_xram_72 [6], RD_xram_72[6]);
  buf(\xm8051_golden_model_1.RD_xram_72 [7], RD_xram_72[7]);
  buf(\xm8051_golden_model_1.RD_xram_71 [0], RD_xram_71[0]);
  buf(\xm8051_golden_model_1.RD_xram_71 [1], RD_xram_71[1]);
  buf(\xm8051_golden_model_1.RD_xram_71 [2], RD_xram_71[2]);
  buf(\xm8051_golden_model_1.RD_xram_71 [3], RD_xram_71[3]);
  buf(\xm8051_golden_model_1.RD_xram_71 [4], RD_xram_71[4]);
  buf(\xm8051_golden_model_1.RD_xram_71 [5], RD_xram_71[5]);
  buf(\xm8051_golden_model_1.RD_xram_71 [6], RD_xram_71[6]);
  buf(\xm8051_golden_model_1.RD_xram_71 [7], RD_xram_71[7]);
  buf(\xm8051_golden_model_1.RD_xram_70 [0], RD_xram_70[0]);
  buf(\xm8051_golden_model_1.RD_xram_70 [1], RD_xram_70[1]);
  buf(\xm8051_golden_model_1.RD_xram_70 [2], RD_xram_70[2]);
  buf(\xm8051_golden_model_1.RD_xram_70 [3], RD_xram_70[3]);
  buf(\xm8051_golden_model_1.RD_xram_70 [4], RD_xram_70[4]);
  buf(\xm8051_golden_model_1.RD_xram_70 [5], RD_xram_70[5]);
  buf(\xm8051_golden_model_1.RD_xram_70 [6], RD_xram_70[6]);
  buf(\xm8051_golden_model_1.RD_xram_70 [7], RD_xram_70[7]);
  buf(\xm8051_golden_model_1.RD_xram_69 [0], RD_xram_69[0]);
  buf(\xm8051_golden_model_1.RD_xram_69 [1], RD_xram_69[1]);
  buf(\xm8051_golden_model_1.RD_xram_69 [2], RD_xram_69[2]);
  buf(\xm8051_golden_model_1.RD_xram_69 [3], RD_xram_69[3]);
  buf(\xm8051_golden_model_1.RD_xram_69 [4], RD_xram_69[4]);
  buf(\xm8051_golden_model_1.RD_xram_69 [5], RD_xram_69[5]);
  buf(\xm8051_golden_model_1.RD_xram_69 [6], RD_xram_69[6]);
  buf(\xm8051_golden_model_1.RD_xram_69 [7], RD_xram_69[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.data_in [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.data_in [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.data_in [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.data_in [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.data_in [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.data_in [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.data_in [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.data_in [7], proc_data_in[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.addr , proc_addr[0]);
  buf(\xm8051_golden_model_1.RD_xram_68 [0], RD_xram_68[0]);
  buf(\xm8051_golden_model_1.RD_xram_68 [1], RD_xram_68[1]);
  buf(\xm8051_golden_model_1.RD_xram_68 [2], RD_xram_68[2]);
  buf(\xm8051_golden_model_1.RD_xram_68 [3], RD_xram_68[3]);
  buf(\xm8051_golden_model_1.RD_xram_68 [4], RD_xram_68[4]);
  buf(\xm8051_golden_model_1.RD_xram_68 [5], RD_xram_68[5]);
  buf(\xm8051_golden_model_1.RD_xram_68 [6], RD_xram_68[6]);
  buf(\xm8051_golden_model_1.RD_xram_68 [7], RD_xram_68[7]);
  buf(\xm8051_golden_model_1.RD_xram_67 [0], RD_xram_67[0]);
  buf(\xm8051_golden_model_1.RD_xram_67 [1], RD_xram_67[1]);
  buf(\xm8051_golden_model_1.RD_xram_67 [2], RD_xram_67[2]);
  buf(\xm8051_golden_model_1.RD_xram_67 [3], RD_xram_67[3]);
  buf(\xm8051_golden_model_1.RD_xram_67 [4], RD_xram_67[4]);
  buf(\xm8051_golden_model_1.RD_xram_67 [5], RD_xram_67[5]);
  buf(\xm8051_golden_model_1.RD_xram_67 [6], RD_xram_67[6]);
  buf(\xm8051_golden_model_1.RD_xram_67 [7], RD_xram_67[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.rst , rst);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_rd_addr_i.clk , clk);
  buf(\xm8051_golden_model_1.RD_xram_66 [0], RD_xram_66[0]);
  buf(\xm8051_golden_model_1.RD_xram_66 [1], RD_xram_66[1]);
  buf(\xm8051_golden_model_1.RD_xram_66 [2], RD_xram_66[2]);
  buf(\xm8051_golden_model_1.RD_xram_66 [3], RD_xram_66[3]);
  buf(\xm8051_golden_model_1.RD_xram_66 [4], RD_xram_66[4]);
  buf(\xm8051_golden_model_1.RD_xram_66 [5], RD_xram_66[5]);
  buf(\xm8051_golden_model_1.RD_xram_66 [6], RD_xram_66[6]);
  buf(\xm8051_golden_model_1.RD_xram_66 [7], RD_xram_66[7]);
  buf(\xm8051_golden_model_1.RD_xram_65 [0], RD_xram_65[0]);
  buf(\xm8051_golden_model_1.RD_xram_65 [1], RD_xram_65[1]);
  buf(\xm8051_golden_model_1.RD_xram_65 [2], RD_xram_65[2]);
  buf(\xm8051_golden_model_1.RD_xram_65 [3], RD_xram_65[3]);
  buf(\xm8051_golden_model_1.RD_xram_65 [4], RD_xram_65[4]);
  buf(\xm8051_golden_model_1.RD_xram_65 [5], RD_xram_65[5]);
  buf(\xm8051_golden_model_1.RD_xram_65 [6], RD_xram_65[6]);
  buf(\xm8051_golden_model_1.RD_xram_65 [7], RD_xram_65[7]);
  buf(\xm8051_golden_model_1.RD_xram_64 [0], RD_xram_64[0]);
  buf(\xm8051_golden_model_1.RD_xram_64 [1], RD_xram_64[1]);
  buf(\xm8051_golden_model_1.RD_xram_64 [2], RD_xram_64[2]);
  buf(\xm8051_golden_model_1.RD_xram_64 [3], RD_xram_64[3]);
  buf(\xm8051_golden_model_1.RD_xram_64 [4], RD_xram_64[4]);
  buf(\xm8051_golden_model_1.RD_xram_64 [5], RD_xram_64[5]);
  buf(\xm8051_golden_model_1.RD_xram_64 [6], RD_xram_64[6]);
  buf(\xm8051_golden_model_1.RD_xram_64 [7], RD_xram_64[7]);
  buf(\xm8051_golden_model_1.RD_xram_63 [0], RD_xram_63[0]);
  buf(\xm8051_golden_model_1.RD_xram_63 [1], RD_xram_63[1]);
  buf(\xm8051_golden_model_1.RD_xram_63 [2], RD_xram_63[2]);
  buf(\xm8051_golden_model_1.RD_xram_63 [3], RD_xram_63[3]);
  buf(\xm8051_golden_model_1.RD_xram_63 [4], RD_xram_63[4]);
  buf(\xm8051_golden_model_1.RD_xram_63 [5], RD_xram_63[5]);
  buf(\xm8051_golden_model_1.RD_xram_63 [6], RD_xram_63[6]);
  buf(\xm8051_golden_model_1.RD_xram_63 [7], RD_xram_63[7]);
  buf(\xm8051_golden_model_1.RD_xram_62 [0], RD_xram_62[0]);
  buf(\xm8051_golden_model_1.RD_xram_62 [1], RD_xram_62[1]);
  buf(\xm8051_golden_model_1.RD_xram_62 [2], RD_xram_62[2]);
  buf(\xm8051_golden_model_1.RD_xram_62 [3], RD_xram_62[3]);
  buf(\xm8051_golden_model_1.RD_xram_62 [4], RD_xram_62[4]);
  buf(\xm8051_golden_model_1.RD_xram_62 [5], RD_xram_62[5]);
  buf(\xm8051_golden_model_1.RD_xram_62 [6], RD_xram_62[6]);
  buf(\xm8051_golden_model_1.RD_xram_62 [7], RD_xram_62[7]);
  buf(\xm8051_golden_model_1.RD_xram_61 [0], RD_xram_61[0]);
  buf(\xm8051_golden_model_1.RD_xram_61 [1], RD_xram_61[1]);
  buf(\xm8051_golden_model_1.RD_xram_61 [2], RD_xram_61[2]);
  buf(\xm8051_golden_model_1.RD_xram_61 [3], RD_xram_61[3]);
  buf(\xm8051_golden_model_1.RD_xram_61 [4], RD_xram_61[4]);
  buf(\xm8051_golden_model_1.RD_xram_61 [5], RD_xram_61[5]);
  buf(\xm8051_golden_model_1.RD_xram_61 [6], RD_xram_61[6]);
  buf(\xm8051_golden_model_1.RD_xram_61 [7], RD_xram_61[7]);
  buf(\xm8051_golden_model_1.RD_xram_60 [0], RD_xram_60[0]);
  buf(\xm8051_golden_model_1.RD_xram_60 [1], RD_xram_60[1]);
  buf(\xm8051_golden_model_1.RD_xram_60 [2], RD_xram_60[2]);
  buf(\xm8051_golden_model_1.RD_xram_60 [3], RD_xram_60[3]);
  buf(\xm8051_golden_model_1.RD_xram_60 [4], RD_xram_60[4]);
  buf(\xm8051_golden_model_1.RD_xram_60 [5], RD_xram_60[5]);
  buf(\xm8051_golden_model_1.RD_xram_60 [6], RD_xram_60[6]);
  buf(\xm8051_golden_model_1.RD_xram_60 [7], RD_xram_60[7]);
  buf(\xm8051_golden_model_1.RD_xram_59 [0], RD_xram_59[0]);
  buf(\xm8051_golden_model_1.RD_xram_59 [1], RD_xram_59[1]);
  buf(\xm8051_golden_model_1.RD_xram_59 [2], RD_xram_59[2]);
  buf(\xm8051_golden_model_1.RD_xram_59 [3], RD_xram_59[3]);
  buf(\xm8051_golden_model_1.RD_xram_59 [4], RD_xram_59[4]);
  buf(\xm8051_golden_model_1.RD_xram_59 [5], RD_xram_59[5]);
  buf(\xm8051_golden_model_1.RD_xram_59 [6], RD_xram_59[6]);
  buf(\xm8051_golden_model_1.RD_xram_59 [7], RD_xram_59[7]);
  buf(\xm8051_golden_model_1.RD_xram_58 [0], RD_xram_58[0]);
  buf(\xm8051_golden_model_1.RD_xram_58 [1], RD_xram_58[1]);
  buf(\xm8051_golden_model_1.RD_xram_58 [2], RD_xram_58[2]);
  buf(\xm8051_golden_model_1.RD_xram_58 [3], RD_xram_58[3]);
  buf(\xm8051_golden_model_1.RD_xram_58 [4], RD_xram_58[4]);
  buf(\xm8051_golden_model_1.RD_xram_58 [5], RD_xram_58[5]);
  buf(\xm8051_golden_model_1.RD_xram_58 [6], RD_xram_58[6]);
  buf(\xm8051_golden_model_1.RD_xram_58 [7], RD_xram_58[7]);
  buf(\xm8051_golden_model_1.RD_xram_57 [0], RD_xram_57[0]);
  buf(\xm8051_golden_model_1.RD_xram_57 [1], RD_xram_57[1]);
  buf(\xm8051_golden_model_1.RD_xram_57 [2], RD_xram_57[2]);
  buf(\xm8051_golden_model_1.RD_xram_57 [3], RD_xram_57[3]);
  buf(\xm8051_golden_model_1.RD_xram_57 [4], RD_xram_57[4]);
  buf(\xm8051_golden_model_1.RD_xram_57 [5], RD_xram_57[5]);
  buf(\xm8051_golden_model_1.RD_xram_57 [6], RD_xram_57[6]);
  buf(\xm8051_golden_model_1.RD_xram_57 [7], RD_xram_57[7]);
  buf(\xm8051_golden_model_1.RD_xram_56 [0], RD_xram_56[0]);
  buf(\xm8051_golden_model_1.RD_xram_56 [1], RD_xram_56[1]);
  buf(\xm8051_golden_model_1.RD_xram_56 [2], RD_xram_56[2]);
  buf(\xm8051_golden_model_1.RD_xram_56 [3], RD_xram_56[3]);
  buf(\xm8051_golden_model_1.RD_xram_56 [4], RD_xram_56[4]);
  buf(\xm8051_golden_model_1.RD_xram_56 [5], RD_xram_56[5]);
  buf(\xm8051_golden_model_1.RD_xram_56 [6], RD_xram_56[6]);
  buf(\xm8051_golden_model_1.RD_xram_56 [7], RD_xram_56[7]);
  buf(\xm8051_golden_model_1.RD_xram_55 [0], RD_xram_55[0]);
  buf(\xm8051_golden_model_1.RD_xram_55 [1], RD_xram_55[1]);
  buf(\xm8051_golden_model_1.RD_xram_55 [2], RD_xram_55[2]);
  buf(\xm8051_golden_model_1.RD_xram_55 [3], RD_xram_55[3]);
  buf(\xm8051_golden_model_1.RD_xram_55 [4], RD_xram_55[4]);
  buf(\xm8051_golden_model_1.RD_xram_55 [5], RD_xram_55[5]);
  buf(\xm8051_golden_model_1.RD_xram_55 [6], RD_xram_55[6]);
  buf(\xm8051_golden_model_1.RD_xram_55 [7], RD_xram_55[7]);
  buf(\xm8051_golden_model_1.RD_xram_54 [0], RD_xram_54[0]);
  buf(\xm8051_golden_model_1.RD_xram_54 [1], RD_xram_54[1]);
  buf(\xm8051_golden_model_1.RD_xram_54 [2], RD_xram_54[2]);
  buf(\xm8051_golden_model_1.RD_xram_54 [3], RD_xram_54[3]);
  buf(\xm8051_golden_model_1.RD_xram_54 [4], RD_xram_54[4]);
  buf(\xm8051_golden_model_1.RD_xram_54 [5], RD_xram_54[5]);
  buf(\xm8051_golden_model_1.RD_xram_54 [6], RD_xram_54[6]);
  buf(\xm8051_golden_model_1.RD_xram_54 [7], RD_xram_54[7]);
  buf(\xm8051_golden_model_1.RD_xram_53 [0], RD_xram_53[0]);
  buf(\xm8051_golden_model_1.RD_xram_53 [1], RD_xram_53[1]);
  buf(\xm8051_golden_model_1.RD_xram_53 [2], RD_xram_53[2]);
  buf(\xm8051_golden_model_1.RD_xram_53 [3], RD_xram_53[3]);
  buf(\xm8051_golden_model_1.RD_xram_53 [4], RD_xram_53[4]);
  buf(\xm8051_golden_model_1.RD_xram_53 [5], RD_xram_53[5]);
  buf(\xm8051_golden_model_1.RD_xram_53 [6], RD_xram_53[6]);
  buf(\xm8051_golden_model_1.RD_xram_53 [7], RD_xram_53[7]);
  buf(\xm8051_golden_model_1.RD_xram_52 [0], RD_xram_52[0]);
  buf(\xm8051_golden_model_1.RD_xram_52 [1], RD_xram_52[1]);
  buf(\xm8051_golden_model_1.RD_xram_52 [2], RD_xram_52[2]);
  buf(\xm8051_golden_model_1.RD_xram_52 [3], RD_xram_52[3]);
  buf(\xm8051_golden_model_1.RD_xram_52 [4], RD_xram_52[4]);
  buf(\xm8051_golden_model_1.RD_xram_52 [5], RD_xram_52[5]);
  buf(\xm8051_golden_model_1.RD_xram_52 [6], RD_xram_52[6]);
  buf(\xm8051_golden_model_1.RD_xram_52 [7], RD_xram_52[7]);
  buf(\xm8051_golden_model_1.RD_xram_51 [0], RD_xram_51[0]);
  buf(\xm8051_golden_model_1.RD_xram_51 [1], RD_xram_51[1]);
  buf(\xm8051_golden_model_1.RD_xram_51 [2], RD_xram_51[2]);
  buf(\xm8051_golden_model_1.RD_xram_51 [3], RD_xram_51[3]);
  buf(\xm8051_golden_model_1.RD_xram_51 [4], RD_xram_51[4]);
  buf(\xm8051_golden_model_1.RD_xram_51 [5], RD_xram_51[5]);
  buf(\xm8051_golden_model_1.RD_xram_51 [6], RD_xram_51[6]);
  buf(\xm8051_golden_model_1.RD_xram_51 [7], RD_xram_51[7]);
  buf(\xm8051_golden_model_1.RD_xram_50 [0], RD_xram_50[0]);
  buf(\xm8051_golden_model_1.RD_xram_50 [1], RD_xram_50[1]);
  buf(\xm8051_golden_model_1.RD_xram_50 [2], RD_xram_50[2]);
  buf(\xm8051_golden_model_1.RD_xram_50 [3], RD_xram_50[3]);
  buf(\xm8051_golden_model_1.RD_xram_50 [4], RD_xram_50[4]);
  buf(\xm8051_golden_model_1.RD_xram_50 [5], RD_xram_50[5]);
  buf(\xm8051_golden_model_1.RD_xram_50 [6], RD_xram_50[6]);
  buf(\xm8051_golden_model_1.RD_xram_50 [7], RD_xram_50[7]);
  buf(\xm8051_golden_model_1.RD_xram_49 [0], RD_xram_49[0]);
  buf(\xm8051_golden_model_1.RD_xram_49 [1], RD_xram_49[1]);
  buf(\xm8051_golden_model_1.RD_xram_49 [2], RD_xram_49[2]);
  buf(\xm8051_golden_model_1.RD_xram_49 [3], RD_xram_49[3]);
  buf(\xm8051_golden_model_1.RD_xram_49 [4], RD_xram_49[4]);
  buf(\xm8051_golden_model_1.RD_xram_49 [5], RD_xram_49[5]);
  buf(\xm8051_golden_model_1.RD_xram_49 [6], RD_xram_49[6]);
  buf(\xm8051_golden_model_1.RD_xram_49 [7], RD_xram_49[7]);
  buf(\xm8051_golden_model_1.RD_xram_48 [0], RD_xram_48[0]);
  buf(\xm8051_golden_model_1.RD_xram_48 [1], RD_xram_48[1]);
  buf(\xm8051_golden_model_1.RD_xram_48 [2], RD_xram_48[2]);
  buf(\xm8051_golden_model_1.RD_xram_48 [3], RD_xram_48[3]);
  buf(\xm8051_golden_model_1.RD_xram_48 [4], RD_xram_48[4]);
  buf(\xm8051_golden_model_1.RD_xram_48 [5], RD_xram_48[5]);
  buf(\xm8051_golden_model_1.RD_xram_48 [6], RD_xram_48[6]);
  buf(\xm8051_golden_model_1.RD_xram_48 [7], RD_xram_48[7]);
  buf(\xm8051_golden_model_1.RD_xram_47 [0], RD_xram_47[0]);
  buf(\xm8051_golden_model_1.RD_xram_47 [1], RD_xram_47[1]);
  buf(\xm8051_golden_model_1.RD_xram_47 [2], RD_xram_47[2]);
  buf(\xm8051_golden_model_1.RD_xram_47 [3], RD_xram_47[3]);
  buf(\xm8051_golden_model_1.RD_xram_47 [4], RD_xram_47[4]);
  buf(\xm8051_golden_model_1.RD_xram_47 [5], RD_xram_47[5]);
  buf(\xm8051_golden_model_1.RD_xram_47 [6], RD_xram_47[6]);
  buf(\xm8051_golden_model_1.RD_xram_47 [7], RD_xram_47[7]);
  buf(\xm8051_golden_model_1.RD_xram_46 [0], RD_xram_46[0]);
  buf(\xm8051_golden_model_1.RD_xram_46 [1], RD_xram_46[1]);
  buf(\xm8051_golden_model_1.RD_xram_46 [2], RD_xram_46[2]);
  buf(\xm8051_golden_model_1.RD_xram_46 [3], RD_xram_46[3]);
  buf(\xm8051_golden_model_1.RD_xram_46 [4], RD_xram_46[4]);
  buf(\xm8051_golden_model_1.RD_xram_46 [5], RD_xram_46[5]);
  buf(\xm8051_golden_model_1.RD_xram_46 [6], RD_xram_46[6]);
  buf(\xm8051_golden_model_1.RD_xram_46 [7], RD_xram_46[7]);
  buf(\xm8051_golden_model_1.RD_xram_45 [0], RD_xram_45[0]);
  buf(\xm8051_golden_model_1.RD_xram_45 [1], RD_xram_45[1]);
  buf(\xm8051_golden_model_1.RD_xram_45 [2], RD_xram_45[2]);
  buf(\xm8051_golden_model_1.RD_xram_45 [3], RD_xram_45[3]);
  buf(\xm8051_golden_model_1.RD_xram_45 [4], RD_xram_45[4]);
  buf(\xm8051_golden_model_1.RD_xram_45 [5], RD_xram_45[5]);
  buf(\xm8051_golden_model_1.RD_xram_45 [6], RD_xram_45[6]);
  buf(\xm8051_golden_model_1.RD_xram_45 [7], RD_xram_45[7]);
  buf(\xm8051_golden_model_1.RD_xram_44 [0], RD_xram_44[0]);
  buf(\xm8051_golden_model_1.RD_xram_44 [1], RD_xram_44[1]);
  buf(\xm8051_golden_model_1.RD_xram_44 [2], RD_xram_44[2]);
  buf(\xm8051_golden_model_1.RD_xram_44 [3], RD_xram_44[3]);
  buf(\xm8051_golden_model_1.RD_xram_44 [4], RD_xram_44[4]);
  buf(\xm8051_golden_model_1.RD_xram_44 [5], RD_xram_44[5]);
  buf(\xm8051_golden_model_1.RD_xram_44 [6], RD_xram_44[6]);
  buf(\xm8051_golden_model_1.RD_xram_44 [7], RD_xram_44[7]);
  buf(\xm8051_golden_model_1.RD_xram_43 [0], RD_xram_43[0]);
  buf(\xm8051_golden_model_1.RD_xram_43 [1], RD_xram_43[1]);
  buf(\xm8051_golden_model_1.RD_xram_43 [2], RD_xram_43[2]);
  buf(\xm8051_golden_model_1.RD_xram_43 [3], RD_xram_43[3]);
  buf(\xm8051_golden_model_1.RD_xram_43 [4], RD_xram_43[4]);
  buf(\xm8051_golden_model_1.RD_xram_43 [5], RD_xram_43[5]);
  buf(\xm8051_golden_model_1.RD_xram_43 [6], RD_xram_43[6]);
  buf(\xm8051_golden_model_1.RD_xram_43 [7], RD_xram_43[7]);
  buf(\xm8051_golden_model_1.RD_xram_42 [0], RD_xram_42[0]);
  buf(\xm8051_golden_model_1.RD_xram_42 [1], RD_xram_42[1]);
  buf(\xm8051_golden_model_1.RD_xram_42 [2], RD_xram_42[2]);
  buf(\xm8051_golden_model_1.RD_xram_42 [3], RD_xram_42[3]);
  buf(\xm8051_golden_model_1.RD_xram_42 [4], RD_xram_42[4]);
  buf(\xm8051_golden_model_1.RD_xram_42 [5], RD_xram_42[5]);
  buf(\xm8051_golden_model_1.RD_xram_42 [6], RD_xram_42[6]);
  buf(\xm8051_golden_model_1.RD_xram_42 [7], RD_xram_42[7]);
  buf(\xm8051_golden_model_1.RD_xram_41 [0], RD_xram_41[0]);
  buf(\xm8051_golden_model_1.RD_xram_41 [1], RD_xram_41[1]);
  buf(\xm8051_golden_model_1.RD_xram_41 [2], RD_xram_41[2]);
  buf(\xm8051_golden_model_1.RD_xram_41 [3], RD_xram_41[3]);
  buf(\xm8051_golden_model_1.RD_xram_41 [4], RD_xram_41[4]);
  buf(\xm8051_golden_model_1.RD_xram_41 [5], RD_xram_41[5]);
  buf(\xm8051_golden_model_1.RD_xram_41 [6], RD_xram_41[6]);
  buf(\xm8051_golden_model_1.RD_xram_41 [7], RD_xram_41[7]);
  buf(\xm8051_golden_model_1.RD_xram_40 [0], RD_xram_40[0]);
  buf(\xm8051_golden_model_1.RD_xram_40 [1], RD_xram_40[1]);
  buf(\xm8051_golden_model_1.RD_xram_40 [2], RD_xram_40[2]);
  buf(\xm8051_golden_model_1.RD_xram_40 [3], RD_xram_40[3]);
  buf(\xm8051_golden_model_1.RD_xram_40 [4], RD_xram_40[4]);
  buf(\xm8051_golden_model_1.RD_xram_40 [5], RD_xram_40[5]);
  buf(\xm8051_golden_model_1.RD_xram_40 [6], RD_xram_40[6]);
  buf(\xm8051_golden_model_1.RD_xram_40 [7], RD_xram_40[7]);
  buf(\xm8051_golden_model_1.RD_xram_39 [0], RD_xram_39[0]);
  buf(\xm8051_golden_model_1.RD_xram_39 [1], RD_xram_39[1]);
  buf(\xm8051_golden_model_1.RD_xram_39 [2], RD_xram_39[2]);
  buf(\xm8051_golden_model_1.RD_xram_39 [3], RD_xram_39[3]);
  buf(\xm8051_golden_model_1.RD_xram_39 [4], RD_xram_39[4]);
  buf(\xm8051_golden_model_1.RD_xram_39 [5], RD_xram_39[5]);
  buf(\xm8051_golden_model_1.RD_xram_39 [6], RD_xram_39[6]);
  buf(\xm8051_golden_model_1.RD_xram_39 [7], RD_xram_39[7]);
  buf(\xm8051_golden_model_1.RD_xram_38 [0], RD_xram_38[0]);
  buf(\xm8051_golden_model_1.RD_xram_38 [1], RD_xram_38[1]);
  buf(\xm8051_golden_model_1.RD_xram_38 [2], RD_xram_38[2]);
  buf(\xm8051_golden_model_1.RD_xram_38 [3], RD_xram_38[3]);
  buf(\xm8051_golden_model_1.RD_xram_38 [4], RD_xram_38[4]);
  buf(\xm8051_golden_model_1.RD_xram_38 [5], RD_xram_38[5]);
  buf(\xm8051_golden_model_1.RD_xram_38 [6], RD_xram_38[6]);
  buf(\xm8051_golden_model_1.RD_xram_38 [7], RD_xram_38[7]);
  buf(\xm8051_golden_model_1.RD_xram_37 [0], RD_xram_37[0]);
  buf(\xm8051_golden_model_1.RD_xram_37 [1], RD_xram_37[1]);
  buf(\xm8051_golden_model_1.RD_xram_37 [2], RD_xram_37[2]);
  buf(\xm8051_golden_model_1.RD_xram_37 [3], RD_xram_37[3]);
  buf(\xm8051_golden_model_1.RD_xram_37 [4], RD_xram_37[4]);
  buf(\xm8051_golden_model_1.RD_xram_37 [5], RD_xram_37[5]);
  buf(\xm8051_golden_model_1.RD_xram_37 [6], RD_xram_37[6]);
  buf(\xm8051_golden_model_1.RD_xram_37 [7], RD_xram_37[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.data_in [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.data_in [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.data_in [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.data_in [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.data_in [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.data_in [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.data_in [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.data_in [7], proc_data_in[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.addr , proc_addr[0]);
  buf(\xm8051_golden_model_1.RD_xram_36 [0], RD_xram_36[0]);
  buf(\xm8051_golden_model_1.RD_xram_36 [1], RD_xram_36[1]);
  buf(\xm8051_golden_model_1.RD_xram_36 [2], RD_xram_36[2]);
  buf(\xm8051_golden_model_1.RD_xram_36 [3], RD_xram_36[3]);
  buf(\xm8051_golden_model_1.RD_xram_36 [4], RD_xram_36[4]);
  buf(\xm8051_golden_model_1.RD_xram_36 [5], RD_xram_36[5]);
  buf(\xm8051_golden_model_1.RD_xram_36 [6], RD_xram_36[6]);
  buf(\xm8051_golden_model_1.RD_xram_36 [7], RD_xram_36[7]);
  buf(\xm8051_golden_model_1.RD_xram_35 [0], RD_xram_35[0]);
  buf(\xm8051_golden_model_1.RD_xram_35 [1], RD_xram_35[1]);
  buf(\xm8051_golden_model_1.RD_xram_35 [2], RD_xram_35[2]);
  buf(\xm8051_golden_model_1.RD_xram_35 [3], RD_xram_35[3]);
  buf(\xm8051_golden_model_1.RD_xram_35 [4], RD_xram_35[4]);
  buf(\xm8051_golden_model_1.RD_xram_35 [5], RD_xram_35[5]);
  buf(\xm8051_golden_model_1.RD_xram_35 [6], RD_xram_35[6]);
  buf(\xm8051_golden_model_1.RD_xram_35 [7], RD_xram_35[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.rst , rst);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_wr_addr_i.clk , clk);
  buf(\xm8051_golden_model_1.RD_xram_34 [0], RD_xram_34[0]);
  buf(\xm8051_golden_model_1.RD_xram_34 [1], RD_xram_34[1]);
  buf(\xm8051_golden_model_1.RD_xram_34 [2], RD_xram_34[2]);
  buf(\xm8051_golden_model_1.RD_xram_34 [3], RD_xram_34[3]);
  buf(\xm8051_golden_model_1.RD_xram_34 [4], RD_xram_34[4]);
  buf(\xm8051_golden_model_1.RD_xram_34 [5], RD_xram_34[5]);
  buf(\xm8051_golden_model_1.RD_xram_34 [6], RD_xram_34[6]);
  buf(\xm8051_golden_model_1.RD_xram_34 [7], RD_xram_34[7]);
  buf(\xm8051_golden_model_1.RD_xram_33 [0], RD_xram_33[0]);
  buf(\xm8051_golden_model_1.RD_xram_33 [1], RD_xram_33[1]);
  buf(\xm8051_golden_model_1.RD_xram_33 [2], RD_xram_33[2]);
  buf(\xm8051_golden_model_1.RD_xram_33 [3], RD_xram_33[3]);
  buf(\xm8051_golden_model_1.RD_xram_33 [4], RD_xram_33[4]);
  buf(\xm8051_golden_model_1.RD_xram_33 [5], RD_xram_33[5]);
  buf(\xm8051_golden_model_1.RD_xram_33 [6], RD_xram_33[6]);
  buf(\xm8051_golden_model_1.RD_xram_33 [7], RD_xram_33[7]);
  buf(\xm8051_golden_model_1.RD_xram_32 [0], RD_xram_32[0]);
  buf(\xm8051_golden_model_1.RD_xram_32 [1], RD_xram_32[1]);
  buf(\xm8051_golden_model_1.RD_xram_32 [2], RD_xram_32[2]);
  buf(\xm8051_golden_model_1.RD_xram_32 [3], RD_xram_32[3]);
  buf(\xm8051_golden_model_1.RD_xram_32 [4], RD_xram_32[4]);
  buf(\xm8051_golden_model_1.RD_xram_32 [5], RD_xram_32[5]);
  buf(\xm8051_golden_model_1.RD_xram_32 [6], RD_xram_32[6]);
  buf(\xm8051_golden_model_1.RD_xram_32 [7], RD_xram_32[7]);
  buf(\xm8051_golden_model_1.RD_xram_31 [0], RD_xram_31[0]);
  buf(\xm8051_golden_model_1.RD_xram_31 [1], RD_xram_31[1]);
  buf(\xm8051_golden_model_1.RD_xram_31 [2], RD_xram_31[2]);
  buf(\xm8051_golden_model_1.RD_xram_31 [3], RD_xram_31[3]);
  buf(\xm8051_golden_model_1.RD_xram_31 [4], RD_xram_31[4]);
  buf(\xm8051_golden_model_1.RD_xram_31 [5], RD_xram_31[5]);
  buf(\xm8051_golden_model_1.RD_xram_31 [6], RD_xram_31[6]);
  buf(\xm8051_golden_model_1.RD_xram_31 [7], RD_xram_31[7]);
  buf(\xm8051_golden_model_1.RD_xram_30 [0], RD_xram_30[0]);
  buf(\xm8051_golden_model_1.RD_xram_30 [1], RD_xram_30[1]);
  buf(\xm8051_golden_model_1.RD_xram_30 [2], RD_xram_30[2]);
  buf(\xm8051_golden_model_1.RD_xram_30 [3], RD_xram_30[3]);
  buf(\xm8051_golden_model_1.RD_xram_30 [4], RD_xram_30[4]);
  buf(\xm8051_golden_model_1.RD_xram_30 [5], RD_xram_30[5]);
  buf(\xm8051_golden_model_1.RD_xram_30 [6], RD_xram_30[6]);
  buf(\xm8051_golden_model_1.RD_xram_30 [7], RD_xram_30[7]);
  buf(\xm8051_golden_model_1.RD_xram_29 [0], RD_xram_29[0]);
  buf(\xm8051_golden_model_1.RD_xram_29 [1], RD_xram_29[1]);
  buf(\xm8051_golden_model_1.RD_xram_29 [2], RD_xram_29[2]);
  buf(\xm8051_golden_model_1.RD_xram_29 [3], RD_xram_29[3]);
  buf(\xm8051_golden_model_1.RD_xram_29 [4], RD_xram_29[4]);
  buf(\xm8051_golden_model_1.RD_xram_29 [5], RD_xram_29[5]);
  buf(\xm8051_golden_model_1.RD_xram_29 [6], RD_xram_29[6]);
  buf(\xm8051_golden_model_1.RD_xram_29 [7], RD_xram_29[7]);
  buf(\xm8051_golden_model_1.RD_xram_28 [0], RD_xram_28[0]);
  buf(\xm8051_golden_model_1.RD_xram_28 [1], RD_xram_28[1]);
  buf(\xm8051_golden_model_1.RD_xram_28 [2], RD_xram_28[2]);
  buf(\xm8051_golden_model_1.RD_xram_28 [3], RD_xram_28[3]);
  buf(\xm8051_golden_model_1.RD_xram_28 [4], RD_xram_28[4]);
  buf(\xm8051_golden_model_1.RD_xram_28 [5], RD_xram_28[5]);
  buf(\xm8051_golden_model_1.RD_xram_28 [6], RD_xram_28[6]);
  buf(\xm8051_golden_model_1.RD_xram_28 [7], RD_xram_28[7]);
  buf(\xm8051_golden_model_1.RD_xram_27 [0], RD_xram_27[0]);
  buf(\xm8051_golden_model_1.RD_xram_27 [1], RD_xram_27[1]);
  buf(\xm8051_golden_model_1.RD_xram_27 [2], RD_xram_27[2]);
  buf(\xm8051_golden_model_1.RD_xram_27 [3], RD_xram_27[3]);
  buf(\xm8051_golden_model_1.RD_xram_27 [4], RD_xram_27[4]);
  buf(\xm8051_golden_model_1.RD_xram_27 [5], RD_xram_27[5]);
  buf(\xm8051_golden_model_1.RD_xram_27 [6], RD_xram_27[6]);
  buf(\xm8051_golden_model_1.RD_xram_27 [7], RD_xram_27[7]);
  buf(\xm8051_golden_model_1.RD_xram_26 [0], RD_xram_26[0]);
  buf(\xm8051_golden_model_1.RD_xram_26 [1], RD_xram_26[1]);
  buf(\xm8051_golden_model_1.RD_xram_26 [2], RD_xram_26[2]);
  buf(\xm8051_golden_model_1.RD_xram_26 [3], RD_xram_26[3]);
  buf(\xm8051_golden_model_1.RD_xram_26 [4], RD_xram_26[4]);
  buf(\xm8051_golden_model_1.RD_xram_26 [5], RD_xram_26[5]);
  buf(\xm8051_golden_model_1.RD_xram_26 [6], RD_xram_26[6]);
  buf(\xm8051_golden_model_1.RD_xram_26 [7], RD_xram_26[7]);
  buf(\xm8051_golden_model_1.RD_xram_25 [0], RD_xram_25[0]);
  buf(\xm8051_golden_model_1.RD_xram_25 [1], RD_xram_25[1]);
  buf(\xm8051_golden_model_1.RD_xram_25 [2], RD_xram_25[2]);
  buf(\xm8051_golden_model_1.RD_xram_25 [3], RD_xram_25[3]);
  buf(\xm8051_golden_model_1.RD_xram_25 [4], RD_xram_25[4]);
  buf(\xm8051_golden_model_1.RD_xram_25 [5], RD_xram_25[5]);
  buf(\xm8051_golden_model_1.RD_xram_25 [6], RD_xram_25[6]);
  buf(\xm8051_golden_model_1.RD_xram_25 [7], RD_xram_25[7]);
  buf(\xm8051_golden_model_1.RD_xram_24 [0], RD_xram_24[0]);
  buf(\xm8051_golden_model_1.RD_xram_24 [1], RD_xram_24[1]);
  buf(\xm8051_golden_model_1.RD_xram_24 [2], RD_xram_24[2]);
  buf(\xm8051_golden_model_1.RD_xram_24 [3], RD_xram_24[3]);
  buf(\xm8051_golden_model_1.RD_xram_24 [4], RD_xram_24[4]);
  buf(\xm8051_golden_model_1.RD_xram_24 [5], RD_xram_24[5]);
  buf(\xm8051_golden_model_1.RD_xram_24 [6], RD_xram_24[6]);
  buf(\xm8051_golden_model_1.RD_xram_24 [7], RD_xram_24[7]);
  buf(\xm8051_golden_model_1.RD_xram_23 [0], RD_xram_23[0]);
  buf(\xm8051_golden_model_1.RD_xram_23 [1], RD_xram_23[1]);
  buf(\xm8051_golden_model_1.RD_xram_23 [2], RD_xram_23[2]);
  buf(\xm8051_golden_model_1.RD_xram_23 [3], RD_xram_23[3]);
  buf(\xm8051_golden_model_1.RD_xram_23 [4], RD_xram_23[4]);
  buf(\xm8051_golden_model_1.RD_xram_23 [5], RD_xram_23[5]);
  buf(\xm8051_golden_model_1.RD_xram_23 [6], RD_xram_23[6]);
  buf(\xm8051_golden_model_1.RD_xram_23 [7], RD_xram_23[7]);
  buf(\xm8051_golden_model_1.RD_xram_22 [0], RD_xram_22[0]);
  buf(\xm8051_golden_model_1.RD_xram_22 [1], RD_xram_22[1]);
  buf(\xm8051_golden_model_1.RD_xram_22 [2], RD_xram_22[2]);
  buf(\xm8051_golden_model_1.RD_xram_22 [3], RD_xram_22[3]);
  buf(\xm8051_golden_model_1.RD_xram_22 [4], RD_xram_22[4]);
  buf(\xm8051_golden_model_1.RD_xram_22 [5], RD_xram_22[5]);
  buf(\xm8051_golden_model_1.RD_xram_22 [6], RD_xram_22[6]);
  buf(\xm8051_golden_model_1.RD_xram_22 [7], RD_xram_22[7]);
  buf(\xm8051_golden_model_1.RD_xram_21 [0], RD_xram_21[0]);
  buf(\xm8051_golden_model_1.RD_xram_21 [1], RD_xram_21[1]);
  buf(\xm8051_golden_model_1.RD_xram_21 [2], RD_xram_21[2]);
  buf(\xm8051_golden_model_1.RD_xram_21 [3], RD_xram_21[3]);
  buf(\xm8051_golden_model_1.RD_xram_21 [4], RD_xram_21[4]);
  buf(\xm8051_golden_model_1.RD_xram_21 [5], RD_xram_21[5]);
  buf(\xm8051_golden_model_1.RD_xram_21 [6], RD_xram_21[6]);
  buf(\xm8051_golden_model_1.RD_xram_21 [7], RD_xram_21[7]);
  buf(\xm8051_golden_model_1.RD_xram_20 [0], RD_xram_20[0]);
  buf(\xm8051_golden_model_1.RD_xram_20 [1], RD_xram_20[1]);
  buf(\xm8051_golden_model_1.RD_xram_20 [2], RD_xram_20[2]);
  buf(\xm8051_golden_model_1.RD_xram_20 [3], RD_xram_20[3]);
  buf(\xm8051_golden_model_1.RD_xram_20 [4], RD_xram_20[4]);
  buf(\xm8051_golden_model_1.RD_xram_20 [5], RD_xram_20[5]);
  buf(\xm8051_golden_model_1.RD_xram_20 [6], RD_xram_20[6]);
  buf(\xm8051_golden_model_1.RD_xram_20 [7], RD_xram_20[7]);
  buf(\xm8051_golden_model_1.RD_xram_19 [0], RD_xram_19[0]);
  buf(\xm8051_golden_model_1.RD_xram_19 [1], RD_xram_19[1]);
  buf(\xm8051_golden_model_1.RD_xram_19 [2], RD_xram_19[2]);
  buf(\xm8051_golden_model_1.RD_xram_19 [3], RD_xram_19[3]);
  buf(\xm8051_golden_model_1.RD_xram_19 [4], RD_xram_19[4]);
  buf(\xm8051_golden_model_1.RD_xram_19 [5], RD_xram_19[5]);
  buf(\xm8051_golden_model_1.RD_xram_19 [6], RD_xram_19[6]);
  buf(\xm8051_golden_model_1.RD_xram_19 [7], RD_xram_19[7]);
  buf(\xm8051_golden_model_1.RD_xram_18 [0], RD_xram_18[0]);
  buf(\xm8051_golden_model_1.RD_xram_18 [1], RD_xram_18[1]);
  buf(\xm8051_golden_model_1.RD_xram_18 [2], RD_xram_18[2]);
  buf(\xm8051_golden_model_1.RD_xram_18 [3], RD_xram_18[3]);
  buf(\xm8051_golden_model_1.RD_xram_18 [4], RD_xram_18[4]);
  buf(\xm8051_golden_model_1.RD_xram_18 [5], RD_xram_18[5]);
  buf(\xm8051_golden_model_1.RD_xram_18 [6], RD_xram_18[6]);
  buf(\xm8051_golden_model_1.RD_xram_18 [7], RD_xram_18[7]);
  buf(\xm8051_golden_model_1.RD_xram_17 [0], RD_xram_17[0]);
  buf(\xm8051_golden_model_1.RD_xram_17 [1], RD_xram_17[1]);
  buf(\xm8051_golden_model_1.RD_xram_17 [2], RD_xram_17[2]);
  buf(\xm8051_golden_model_1.RD_xram_17 [3], RD_xram_17[3]);
  buf(\xm8051_golden_model_1.RD_xram_17 [4], RD_xram_17[4]);
  buf(\xm8051_golden_model_1.RD_xram_17 [5], RD_xram_17[5]);
  buf(\xm8051_golden_model_1.RD_xram_17 [6], RD_xram_17[6]);
  buf(\xm8051_golden_model_1.RD_xram_17 [7], RD_xram_17[7]);
  buf(\xm8051_golden_model_1.RD_xram_16 [0], RD_xram_16[0]);
  buf(\xm8051_golden_model_1.RD_xram_16 [1], RD_xram_16[1]);
  buf(\xm8051_golden_model_1.RD_xram_16 [2], RD_xram_16[2]);
  buf(\xm8051_golden_model_1.RD_xram_16 [3], RD_xram_16[3]);
  buf(\xm8051_golden_model_1.RD_xram_16 [4], RD_xram_16[4]);
  buf(\xm8051_golden_model_1.RD_xram_16 [5], RD_xram_16[5]);
  buf(\xm8051_golden_model_1.RD_xram_16 [6], RD_xram_16[6]);
  buf(\xm8051_golden_model_1.RD_xram_16 [7], RD_xram_16[7]);
  buf(\xm8051_golden_model_1.RD_xram_15 [0], RD_xram_15[0]);
  buf(\xm8051_golden_model_1.RD_xram_15 [1], RD_xram_15[1]);
  buf(\xm8051_golden_model_1.RD_xram_15 [2], RD_xram_15[2]);
  buf(\xm8051_golden_model_1.RD_xram_15 [3], RD_xram_15[3]);
  buf(\xm8051_golden_model_1.RD_xram_15 [4], RD_xram_15[4]);
  buf(\xm8051_golden_model_1.RD_xram_15 [5], RD_xram_15[5]);
  buf(\xm8051_golden_model_1.RD_xram_15 [6], RD_xram_15[6]);
  buf(\xm8051_golden_model_1.RD_xram_15 [7], RD_xram_15[7]);
  buf(\xm8051_golden_model_1.RD_xram_14 [0], RD_xram_14[0]);
  buf(\xm8051_golden_model_1.RD_xram_14 [1], RD_xram_14[1]);
  buf(\xm8051_golden_model_1.RD_xram_14 [2], RD_xram_14[2]);
  buf(\xm8051_golden_model_1.RD_xram_14 [3], RD_xram_14[3]);
  buf(\xm8051_golden_model_1.RD_xram_14 [4], RD_xram_14[4]);
  buf(\xm8051_golden_model_1.RD_xram_14 [5], RD_xram_14[5]);
  buf(\xm8051_golden_model_1.RD_xram_14 [6], RD_xram_14[6]);
  buf(\xm8051_golden_model_1.RD_xram_14 [7], RD_xram_14[7]);
  buf(\xm8051_golden_model_1.RD_xram_13 [0], RD_xram_13[0]);
  buf(\xm8051_golden_model_1.RD_xram_13 [1], RD_xram_13[1]);
  buf(\xm8051_golden_model_1.RD_xram_13 [2], RD_xram_13[2]);
  buf(\xm8051_golden_model_1.RD_xram_13 [3], RD_xram_13[3]);
  buf(\xm8051_golden_model_1.RD_xram_13 [4], RD_xram_13[4]);
  buf(\xm8051_golden_model_1.RD_xram_13 [5], RD_xram_13[5]);
  buf(\xm8051_golden_model_1.RD_xram_13 [6], RD_xram_13[6]);
  buf(\xm8051_golden_model_1.RD_xram_13 [7], RD_xram_13[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.data_in [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.data_in [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.data_in [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.data_in [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.data_in [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.data_in [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.data_in [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.data_in [7], proc_data_in[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.addr , proc_addr[0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.rst , rst);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.clk , clk);
  buf(\xm8051_golden_model_1.RD_xram_12 [0], RD_xram_12[0]);
  buf(\xm8051_golden_model_1.RD_xram_12 [1], RD_xram_12[1]);
  buf(\xm8051_golden_model_1.RD_xram_12 [2], RD_xram_12[2]);
  buf(\xm8051_golden_model_1.RD_xram_12 [3], RD_xram_12[3]);
  buf(\xm8051_golden_model_1.RD_xram_12 [4], RD_xram_12[4]);
  buf(\xm8051_golden_model_1.RD_xram_12 [5], RD_xram_12[5]);
  buf(\xm8051_golden_model_1.RD_xram_12 [6], RD_xram_12[6]);
  buf(\xm8051_golden_model_1.RD_xram_12 [7], RD_xram_12[7]);
  buf(\xm8051_golden_model_1.RD_xram_11 [0], RD_xram_11[0]);
  buf(\xm8051_golden_model_1.RD_xram_11 [1], RD_xram_11[1]);
  buf(\xm8051_golden_model_1.RD_xram_11 [2], RD_xram_11[2]);
  buf(\xm8051_golden_model_1.RD_xram_11 [3], RD_xram_11[3]);
  buf(\xm8051_golden_model_1.RD_xram_11 [4], RD_xram_11[4]);
  buf(\xm8051_golden_model_1.RD_xram_11 [5], RD_xram_11[5]);
  buf(\xm8051_golden_model_1.RD_xram_11 [6], RD_xram_11[6]);
  buf(\xm8051_golden_model_1.RD_xram_11 [7], RD_xram_11[7]);
  buf(\xm8051_golden_model_1.RD_xram_10 [0], RD_xram_10[0]);
  buf(\xm8051_golden_model_1.RD_xram_10 [1], RD_xram_10[1]);
  buf(\xm8051_golden_model_1.RD_xram_10 [2], RD_xram_10[2]);
  buf(\xm8051_golden_model_1.RD_xram_10 [3], RD_xram_10[3]);
  buf(\xm8051_golden_model_1.RD_xram_10 [4], RD_xram_10[4]);
  buf(\xm8051_golden_model_1.RD_xram_10 [5], RD_xram_10[5]);
  buf(\xm8051_golden_model_1.RD_xram_10 [6], RD_xram_10[6]);
  buf(\xm8051_golden_model_1.RD_xram_10 [7], RD_xram_10[7]);
  buf(\xm8051_golden_model_1.RD_xram_9 [0], RD_xram_9[0]);
  buf(\xm8051_golden_model_1.RD_xram_9 [1], RD_xram_9[1]);
  buf(\xm8051_golden_model_1.RD_xram_9 [2], RD_xram_9[2]);
  buf(\xm8051_golden_model_1.RD_xram_9 [3], RD_xram_9[3]);
  buf(\xm8051_golden_model_1.RD_xram_9 [4], RD_xram_9[4]);
  buf(\xm8051_golden_model_1.RD_xram_9 [5], RD_xram_9[5]);
  buf(\xm8051_golden_model_1.RD_xram_9 [6], RD_xram_9[6]);
  buf(\xm8051_golden_model_1.RD_xram_9 [7], RD_xram_9[7]);
  buf(\xm8051_golden_model_1.RD_xram_8 [0], RD_xram_8[0]);
  buf(\xm8051_golden_model_1.RD_xram_8 [1], RD_xram_8[1]);
  buf(\xm8051_golden_model_1.RD_xram_8 [2], RD_xram_8[2]);
  buf(\xm8051_golden_model_1.RD_xram_8 [3], RD_xram_8[3]);
  buf(\xm8051_golden_model_1.RD_xram_8 [4], RD_xram_8[4]);
  buf(\xm8051_golden_model_1.RD_xram_8 [5], RD_xram_8[5]);
  buf(\xm8051_golden_model_1.RD_xram_8 [6], RD_xram_8[6]);
  buf(\xm8051_golden_model_1.RD_xram_8 [7], RD_xram_8[7]);
  buf(\xm8051_golden_model_1.RD_xram_7 [0], RD_xram_7[0]);
  buf(\xm8051_golden_model_1.RD_xram_7 [1], RD_xram_7[1]);
  buf(\xm8051_golden_model_1.RD_xram_7 [2], RD_xram_7[2]);
  buf(\xm8051_golden_model_1.RD_xram_7 [3], RD_xram_7[3]);
  buf(\xm8051_golden_model_1.RD_xram_7 [4], RD_xram_7[4]);
  buf(\xm8051_golden_model_1.RD_xram_7 [5], RD_xram_7[5]);
  buf(\xm8051_golden_model_1.RD_xram_7 [6], RD_xram_7[6]);
  buf(\xm8051_golden_model_1.RD_xram_7 [7], RD_xram_7[7]);
  buf(\xm8051_golden_model_1.RD_xram_6 [0], RD_xram_6[0]);
  buf(\xm8051_golden_model_1.RD_xram_6 [1], RD_xram_6[1]);
  buf(\xm8051_golden_model_1.RD_xram_6 [2], RD_xram_6[2]);
  buf(\xm8051_golden_model_1.RD_xram_6 [3], RD_xram_6[3]);
  buf(\xm8051_golden_model_1.RD_xram_6 [4], RD_xram_6[4]);
  buf(\xm8051_golden_model_1.RD_xram_6 [5], RD_xram_6[5]);
  buf(\xm8051_golden_model_1.RD_xram_6 [6], RD_xram_6[6]);
  buf(\xm8051_golden_model_1.RD_xram_6 [7], RD_xram_6[7]);
  buf(\xm8051_golden_model_1.RD_xram_5 [0], RD_xram_5[0]);
  buf(\xm8051_golden_model_1.RD_xram_5 [1], RD_xram_5[1]);
  buf(\xm8051_golden_model_1.RD_xram_5 [2], RD_xram_5[2]);
  buf(\xm8051_golden_model_1.RD_xram_5 [3], RD_xram_5[3]);
  buf(\xm8051_golden_model_1.RD_xram_5 [4], RD_xram_5[4]);
  buf(\xm8051_golden_model_1.RD_xram_5 [5], RD_xram_5[5]);
  buf(\xm8051_golden_model_1.RD_xram_5 [6], RD_xram_5[6]);
  buf(\xm8051_golden_model_1.RD_xram_5 [7], RD_xram_5[7]);
  buf(\xm8051_golden_model_1.RD_xram_4 [0], RD_xram_4[0]);
  buf(\xm8051_golden_model_1.RD_xram_4 [1], RD_xram_4[1]);
  buf(\xm8051_golden_model_1.RD_xram_4 [2], RD_xram_4[2]);
  buf(\xm8051_golden_model_1.RD_xram_4 [3], RD_xram_4[3]);
  buf(\xm8051_golden_model_1.RD_xram_4 [4], RD_xram_4[4]);
  buf(\xm8051_golden_model_1.RD_xram_4 [5], RD_xram_4[5]);
  buf(\xm8051_golden_model_1.RD_xram_4 [6], RD_xram_4[6]);
  buf(\xm8051_golden_model_1.RD_xram_4 [7], RD_xram_4[7]);
  buf(\xm8051_golden_model_1.RD_xram_3 [0], RD_xram_3[0]);
  buf(\xm8051_golden_model_1.RD_xram_3 [1], RD_xram_3[1]);
  buf(\xm8051_golden_model_1.RD_xram_3 [2], RD_xram_3[2]);
  buf(\xm8051_golden_model_1.RD_xram_3 [3], RD_xram_3[3]);
  buf(\xm8051_golden_model_1.RD_xram_3 [4], RD_xram_3[4]);
  buf(\xm8051_golden_model_1.RD_xram_3 [5], RD_xram_3[5]);
  buf(\xm8051_golden_model_1.RD_xram_3 [6], RD_xram_3[6]);
  buf(\xm8051_golden_model_1.RD_xram_3 [7], RD_xram_3[7]);
  buf(\xm8051_golden_model_1.RD_xram_2 [0], RD_xram_2[0]);
  buf(\xm8051_golden_model_1.RD_xram_2 [1], RD_xram_2[1]);
  buf(\xm8051_golden_model_1.RD_xram_2 [2], RD_xram_2[2]);
  buf(\xm8051_golden_model_1.RD_xram_2 [3], RD_xram_2[3]);
  buf(\xm8051_golden_model_1.RD_xram_2 [4], RD_xram_2[4]);
  buf(\xm8051_golden_model_1.RD_xram_2 [5], RD_xram_2[5]);
  buf(\xm8051_golden_model_1.RD_xram_2 [6], RD_xram_2[6]);
  buf(\xm8051_golden_model_1.RD_xram_2 [7], RD_xram_2[7]);
  buf(\xm8051_golden_model_1.RD_xram_1 [0], RD_xram_1[0]);
  buf(\xm8051_golden_model_1.RD_xram_1 [1], RD_xram_1[1]);
  buf(\xm8051_golden_model_1.RD_xram_1 [2], RD_xram_1[2]);
  buf(\xm8051_golden_model_1.RD_xram_1 [3], RD_xram_1[3]);
  buf(\xm8051_golden_model_1.RD_xram_1 [4], RD_xram_1[4]);
  buf(\xm8051_golden_model_1.RD_xram_1 [5], RD_xram_1[5]);
  buf(\xm8051_golden_model_1.RD_xram_1 [6], RD_xram_1[6]);
  buf(\xm8051_golden_model_1.RD_xram_1 [7], RD_xram_1[7]);
  buf(\xm8051_golden_model_1.RD_xram_0 [0], RD_xram_0[0]);
  buf(\xm8051_golden_model_1.RD_xram_0 [1], RD_xram_0[1]);
  buf(\xm8051_golden_model_1.RD_xram_0 [2], RD_xram_0[2]);
  buf(\xm8051_golden_model_1.RD_xram_0 [3], RD_xram_0[3]);
  buf(\xm8051_golden_model_1.RD_xram_0 [4], RD_xram_0[4]);
  buf(\xm8051_golden_model_1.RD_xram_0 [5], RD_xram_0[5]);
  buf(\xm8051_golden_model_1.RD_xram_0 [6], RD_xram_0[6]);
  buf(\xm8051_golden_model_1.RD_xram_0 [7], RD_xram_0[7]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [0], input_sha_func_55[0]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [1], input_sha_func_55[1]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [2], input_sha_func_55[2]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [3], input_sha_func_55[3]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [4], input_sha_func_55[4]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [5], input_sha_func_55[5]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [6], input_sha_func_55[6]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [7], input_sha_func_55[7]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [8], input_sha_func_55[8]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [9], input_sha_func_55[9]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [10], input_sha_func_55[10]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [11], input_sha_func_55[11]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [12], input_sha_func_55[12]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [13], input_sha_func_55[13]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [14], input_sha_func_55[14]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [15], input_sha_func_55[15]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [16], input_sha_func_55[16]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [17], input_sha_func_55[17]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [18], input_sha_func_55[18]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [19], input_sha_func_55[19]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [20], input_sha_func_55[20]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [21], input_sha_func_55[21]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [22], input_sha_func_55[22]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [23], input_sha_func_55[23]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [24], input_sha_func_55[24]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [25], input_sha_func_55[25]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [26], input_sha_func_55[26]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [27], input_sha_func_55[27]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [28], input_sha_func_55[28]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [29], input_sha_func_55[29]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [30], input_sha_func_55[30]);
  buf(\xm8051_golden_model_1.input_sha_func_55 [31], input_sha_func_55[31]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [0], input_sha_func_54[0]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [1], input_sha_func_54[1]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [2], input_sha_func_54[2]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [3], input_sha_func_54[3]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [4], input_sha_func_54[4]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [5], input_sha_func_54[5]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [6], input_sha_func_54[6]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [7], input_sha_func_54[7]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [8], input_sha_func_54[8]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [9], input_sha_func_54[9]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [10], input_sha_func_54[10]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [11], input_sha_func_54[11]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [12], input_sha_func_54[12]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [13], input_sha_func_54[13]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [14], input_sha_func_54[14]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [15], input_sha_func_54[15]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [16], input_sha_func_54[16]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [17], input_sha_func_54[17]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [18], input_sha_func_54[18]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [19], input_sha_func_54[19]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [20], input_sha_func_54[20]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [21], input_sha_func_54[21]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [22], input_sha_func_54[22]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [23], input_sha_func_54[23]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [24], input_sha_func_54[24]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [25], input_sha_func_54[25]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [26], input_sha_func_54[26]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [27], input_sha_func_54[27]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [28], input_sha_func_54[28]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [29], input_sha_func_54[29]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [30], input_sha_func_54[30]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [31], input_sha_func_54[31]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [32], input_sha_func_54[32]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [33], input_sha_func_54[33]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [34], input_sha_func_54[34]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [35], input_sha_func_54[35]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [36], input_sha_func_54[36]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [37], input_sha_func_54[37]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [38], input_sha_func_54[38]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [39], input_sha_func_54[39]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [40], input_sha_func_54[40]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [41], input_sha_func_54[41]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [42], input_sha_func_54[42]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [43], input_sha_func_54[43]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [44], input_sha_func_54[44]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [45], input_sha_func_54[45]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [46], input_sha_func_54[46]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [47], input_sha_func_54[47]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [48], input_sha_func_54[48]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [49], input_sha_func_54[49]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [50], input_sha_func_54[50]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [51], input_sha_func_54[51]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [52], input_sha_func_54[52]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [53], input_sha_func_54[53]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [54], input_sha_func_54[54]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [55], input_sha_func_54[55]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [56], input_sha_func_54[56]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [57], input_sha_func_54[57]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [58], input_sha_func_54[58]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [59], input_sha_func_54[59]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [60], input_sha_func_54[60]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [61], input_sha_func_54[61]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [62], input_sha_func_54[62]);
  buf(\xm8051_golden_model_1.input_sha_func_54 [63], input_sha_func_54[63]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [0], input_sha_func_53[0]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [1], input_sha_func_53[1]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [2], input_sha_func_53[2]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [3], input_sha_func_53[3]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [4], input_sha_func_53[4]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [5], input_sha_func_53[5]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [6], input_sha_func_53[6]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [7], input_sha_func_53[7]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [8], input_sha_func_53[8]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [9], input_sha_func_53[9]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [10], input_sha_func_53[10]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [11], input_sha_func_53[11]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [12], input_sha_func_53[12]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [13], input_sha_func_53[13]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [14], input_sha_func_53[14]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [15], input_sha_func_53[15]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [16], input_sha_func_53[16]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [17], input_sha_func_53[17]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [18], input_sha_func_53[18]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [19], input_sha_func_53[19]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [20], input_sha_func_53[20]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [21], input_sha_func_53[21]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [22], input_sha_func_53[22]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [23], input_sha_func_53[23]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [24], input_sha_func_53[24]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [25], input_sha_func_53[25]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [26], input_sha_func_53[26]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [27], input_sha_func_53[27]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [28], input_sha_func_53[28]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [29], input_sha_func_53[29]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [30], input_sha_func_53[30]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [31], input_sha_func_53[31]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [32], input_sha_func_53[32]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [33], input_sha_func_53[33]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [34], input_sha_func_53[34]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [35], input_sha_func_53[35]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [36], input_sha_func_53[36]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [37], input_sha_func_53[37]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [38], input_sha_func_53[38]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [39], input_sha_func_53[39]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [40], input_sha_func_53[40]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [41], input_sha_func_53[41]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [42], input_sha_func_53[42]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [43], input_sha_func_53[43]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [44], input_sha_func_53[44]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [45], input_sha_func_53[45]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [46], input_sha_func_53[46]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [47], input_sha_func_53[47]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [48], input_sha_func_53[48]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [49], input_sha_func_53[49]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [50], input_sha_func_53[50]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [51], input_sha_func_53[51]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [52], input_sha_func_53[52]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [53], input_sha_func_53[53]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [54], input_sha_func_53[54]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [55], input_sha_func_53[55]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [56], input_sha_func_53[56]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [57], input_sha_func_53[57]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [58], input_sha_func_53[58]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [59], input_sha_func_53[59]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [60], input_sha_func_53[60]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [61], input_sha_func_53[61]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [62], input_sha_func_53[62]);
  buf(\xm8051_golden_model_1.input_sha_func_53 [63], input_sha_func_53[63]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [0], input_aes_func_52[0]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [1], input_aes_func_52[1]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [2], input_aes_func_52[2]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [3], input_aes_func_52[3]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [4], input_aes_func_52[4]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [5], input_aes_func_52[5]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [6], input_aes_func_52[6]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [7], input_aes_func_52[7]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [8], input_aes_func_52[8]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [9], input_aes_func_52[9]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [10], input_aes_func_52[10]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [11], input_aes_func_52[11]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [12], input_aes_func_52[12]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [13], input_aes_func_52[13]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [14], input_aes_func_52[14]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [15], input_aes_func_52[15]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [16], input_aes_func_52[16]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [17], input_aes_func_52[17]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [18], input_aes_func_52[18]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [19], input_aes_func_52[19]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [20], input_aes_func_52[20]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [21], input_aes_func_52[21]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [22], input_aes_func_52[22]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [23], input_aes_func_52[23]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [24], input_aes_func_52[24]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [25], input_aes_func_52[25]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [26], input_aes_func_52[26]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [27], input_aes_func_52[27]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [28], input_aes_func_52[28]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [29], input_aes_func_52[29]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [30], input_aes_func_52[30]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [31], input_aes_func_52[31]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [32], input_aes_func_52[32]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [33], input_aes_func_52[33]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [34], input_aes_func_52[34]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [35], input_aes_func_52[35]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [36], input_aes_func_52[36]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [37], input_aes_func_52[37]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [38], input_aes_func_52[38]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [39], input_aes_func_52[39]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [40], input_aes_func_52[40]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [41], input_aes_func_52[41]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [42], input_aes_func_52[42]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [43], input_aes_func_52[43]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [44], input_aes_func_52[44]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [45], input_aes_func_52[45]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [46], input_aes_func_52[46]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [47], input_aes_func_52[47]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [48], input_aes_func_52[48]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [49], input_aes_func_52[49]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [50], input_aes_func_52[50]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [51], input_aes_func_52[51]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [52], input_aes_func_52[52]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [53], input_aes_func_52[53]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [54], input_aes_func_52[54]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [55], input_aes_func_52[55]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [56], input_aes_func_52[56]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [57], input_aes_func_52[57]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [58], input_aes_func_52[58]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [59], input_aes_func_52[59]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [60], input_aes_func_52[60]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [61], input_aes_func_52[61]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [62], input_aes_func_52[62]);
  buf(\xm8051_golden_model_1.input_aes_func_52 [63], input_aes_func_52[63]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [0], input_aes_func_51[0]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [1], input_aes_func_51[1]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [2], input_aes_func_51[2]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [3], input_aes_func_51[3]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [4], input_aes_func_51[4]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [5], input_aes_func_51[5]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [6], input_aes_func_51[6]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [7], input_aes_func_51[7]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [8], input_aes_func_51[8]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [9], input_aes_func_51[9]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [10], input_aes_func_51[10]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [11], input_aes_func_51[11]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [12], input_aes_func_51[12]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [13], input_aes_func_51[13]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [14], input_aes_func_51[14]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [15], input_aes_func_51[15]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [16], input_aes_func_51[16]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [17], input_aes_func_51[17]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [18], input_aes_func_51[18]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [19], input_aes_func_51[19]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [20], input_aes_func_51[20]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [21], input_aes_func_51[21]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [22], input_aes_func_51[22]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [23], input_aes_func_51[23]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [24], input_aes_func_51[24]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [25], input_aes_func_51[25]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [26], input_aes_func_51[26]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [27], input_aes_func_51[27]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [28], input_aes_func_51[28]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [29], input_aes_func_51[29]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [30], input_aes_func_51[30]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [31], input_aes_func_51[31]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [32], input_aes_func_51[32]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [33], input_aes_func_51[33]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [34], input_aes_func_51[34]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [35], input_aes_func_51[35]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [36], input_aes_func_51[36]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [37], input_aes_func_51[37]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [38], input_aes_func_51[38]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [39], input_aes_func_51[39]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [40], input_aes_func_51[40]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [41], input_aes_func_51[41]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [42], input_aes_func_51[42]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [43], input_aes_func_51[43]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [44], input_aes_func_51[44]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [45], input_aes_func_51[45]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [46], input_aes_func_51[46]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [47], input_aes_func_51[47]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [48], input_aes_func_51[48]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [49], input_aes_func_51[49]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [50], input_aes_func_51[50]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [51], input_aes_func_51[51]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [52], input_aes_func_51[52]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [53], input_aes_func_51[53]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [54], input_aes_func_51[54]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [55], input_aes_func_51[55]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [56], input_aes_func_51[56]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [57], input_aes_func_51[57]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [58], input_aes_func_51[58]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [59], input_aes_func_51[59]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [60], input_aes_func_51[60]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [61], input_aes_func_51[61]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [62], input_aes_func_51[62]);
  buf(\xm8051_golden_model_1.input_aes_func_51 [63], input_aes_func_51[63]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [0], input_sha_func_50[0]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [1], input_sha_func_50[1]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [2], input_sha_func_50[2]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [3], input_sha_func_50[3]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [4], input_sha_func_50[4]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [5], input_sha_func_50[5]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [6], input_sha_func_50[6]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [7], input_sha_func_50[7]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [8], input_sha_func_50[8]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [9], input_sha_func_50[9]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [10], input_sha_func_50[10]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [11], input_sha_func_50[11]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [12], input_sha_func_50[12]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [13], input_sha_func_50[13]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [14], input_sha_func_50[14]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [15], input_sha_func_50[15]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [16], input_sha_func_50[16]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [17], input_sha_func_50[17]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [18], input_sha_func_50[18]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [19], input_sha_func_50[19]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [20], input_sha_func_50[20]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [21], input_sha_func_50[21]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [22], input_sha_func_50[22]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [23], input_sha_func_50[23]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [24], input_sha_func_50[24]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [25], input_sha_func_50[25]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [26], input_sha_func_50[26]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [27], input_sha_func_50[27]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [28], input_sha_func_50[28]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [29], input_sha_func_50[29]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [30], input_sha_func_50[30]);
  buf(\xm8051_golden_model_1.input_sha_func_50 [31], input_sha_func_50[31]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [0], input_sha_func_49[0]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [1], input_sha_func_49[1]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [2], input_sha_func_49[2]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [3], input_sha_func_49[3]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [4], input_sha_func_49[4]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [5], input_sha_func_49[5]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [6], input_sha_func_49[6]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [7], input_sha_func_49[7]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [8], input_sha_func_49[8]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [9], input_sha_func_49[9]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [10], input_sha_func_49[10]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [11], input_sha_func_49[11]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [12], input_sha_func_49[12]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [13], input_sha_func_49[13]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [14], input_sha_func_49[14]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [15], input_sha_func_49[15]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [16], input_sha_func_49[16]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [17], input_sha_func_49[17]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [18], input_sha_func_49[18]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [19], input_sha_func_49[19]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [20], input_sha_func_49[20]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [21], input_sha_func_49[21]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [22], input_sha_func_49[22]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [23], input_sha_func_49[23]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [24], input_sha_func_49[24]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [25], input_sha_func_49[25]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [26], input_sha_func_49[26]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [27], input_sha_func_49[27]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [28], input_sha_func_49[28]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [29], input_sha_func_49[29]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [30], input_sha_func_49[30]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [31], input_sha_func_49[31]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [32], input_sha_func_49[32]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [33], input_sha_func_49[33]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [34], input_sha_func_49[34]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [35], input_sha_func_49[35]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [36], input_sha_func_49[36]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [37], input_sha_func_49[37]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [38], input_sha_func_49[38]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [39], input_sha_func_49[39]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [40], input_sha_func_49[40]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [41], input_sha_func_49[41]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [42], input_sha_func_49[42]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [43], input_sha_func_49[43]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [44], input_sha_func_49[44]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [45], input_sha_func_49[45]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [46], input_sha_func_49[46]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [47], input_sha_func_49[47]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [48], input_sha_func_49[48]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [49], input_sha_func_49[49]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [50], input_sha_func_49[50]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [51], input_sha_func_49[51]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [52], input_sha_func_49[52]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [53], input_sha_func_49[53]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [54], input_sha_func_49[54]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [55], input_sha_func_49[55]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [56], input_sha_func_49[56]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [57], input_sha_func_49[57]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [58], input_sha_func_49[58]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [59], input_sha_func_49[59]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [60], input_sha_func_49[60]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [61], input_sha_func_49[61]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [62], input_sha_func_49[62]);
  buf(\xm8051_golden_model_1.input_sha_func_49 [63], input_sha_func_49[63]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [0], input_sha_func_48[0]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [1], input_sha_func_48[1]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [2], input_sha_func_48[2]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [3], input_sha_func_48[3]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [4], input_sha_func_48[4]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [5], input_sha_func_48[5]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [6], input_sha_func_48[6]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [7], input_sha_func_48[7]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [8], input_sha_func_48[8]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [9], input_sha_func_48[9]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [10], input_sha_func_48[10]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [11], input_sha_func_48[11]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [12], input_sha_func_48[12]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [13], input_sha_func_48[13]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [14], input_sha_func_48[14]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [15], input_sha_func_48[15]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [16], input_sha_func_48[16]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [17], input_sha_func_48[17]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [18], input_sha_func_48[18]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [19], input_sha_func_48[19]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [20], input_sha_func_48[20]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [21], input_sha_func_48[21]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [22], input_sha_func_48[22]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [23], input_sha_func_48[23]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [24], input_sha_func_48[24]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [25], input_sha_func_48[25]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [26], input_sha_func_48[26]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [27], input_sha_func_48[27]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [28], input_sha_func_48[28]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [29], input_sha_func_48[29]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [30], input_sha_func_48[30]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [31], input_sha_func_48[31]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [32], input_sha_func_48[32]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [33], input_sha_func_48[33]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [34], input_sha_func_48[34]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [35], input_sha_func_48[35]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [36], input_sha_func_48[36]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [37], input_sha_func_48[37]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [38], input_sha_func_48[38]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [39], input_sha_func_48[39]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [40], input_sha_func_48[40]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [41], input_sha_func_48[41]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [42], input_sha_func_48[42]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [43], input_sha_func_48[43]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [44], input_sha_func_48[44]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [45], input_sha_func_48[45]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [46], input_sha_func_48[46]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [47], input_sha_func_48[47]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [48], input_sha_func_48[48]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [49], input_sha_func_48[49]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [50], input_sha_func_48[50]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [51], input_sha_func_48[51]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [52], input_sha_func_48[52]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [53], input_sha_func_48[53]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [54], input_sha_func_48[54]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [55], input_sha_func_48[55]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [56], input_sha_func_48[56]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [57], input_sha_func_48[57]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [58], input_sha_func_48[58]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [59], input_sha_func_48[59]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [60], input_sha_func_48[60]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [61], input_sha_func_48[61]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [62], input_sha_func_48[62]);
  buf(\xm8051_golden_model_1.input_sha_func_48 [63], input_sha_func_48[63]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [0], input_sha_func_47[0]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [1], input_sha_func_47[1]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [2], input_sha_func_47[2]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [3], input_sha_func_47[3]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [4], input_sha_func_47[4]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [5], input_sha_func_47[5]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [6], input_sha_func_47[6]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [7], input_sha_func_47[7]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [8], input_sha_func_47[8]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [9], input_sha_func_47[9]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [10], input_sha_func_47[10]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [11], input_sha_func_47[11]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [12], input_sha_func_47[12]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [13], input_sha_func_47[13]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [14], input_sha_func_47[14]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [15], input_sha_func_47[15]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [16], input_sha_func_47[16]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [17], input_sha_func_47[17]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [18], input_sha_func_47[18]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [19], input_sha_func_47[19]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [20], input_sha_func_47[20]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [21], input_sha_func_47[21]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [22], input_sha_func_47[22]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [23], input_sha_func_47[23]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [24], input_sha_func_47[24]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [25], input_sha_func_47[25]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [26], input_sha_func_47[26]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [27], input_sha_func_47[27]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [28], input_sha_func_47[28]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [29], input_sha_func_47[29]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [30], input_sha_func_47[30]);
  buf(\xm8051_golden_model_1.input_sha_func_47 [31], input_sha_func_47[31]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [0], input_sha_func_46[0]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [1], input_sha_func_46[1]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [2], input_sha_func_46[2]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [3], input_sha_func_46[3]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [4], input_sha_func_46[4]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [5], input_sha_func_46[5]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [6], input_sha_func_46[6]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [7], input_sha_func_46[7]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [8], input_sha_func_46[8]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [9], input_sha_func_46[9]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [10], input_sha_func_46[10]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [11], input_sha_func_46[11]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [12], input_sha_func_46[12]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [13], input_sha_func_46[13]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [14], input_sha_func_46[14]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [15], input_sha_func_46[15]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [16], input_sha_func_46[16]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [17], input_sha_func_46[17]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [18], input_sha_func_46[18]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [19], input_sha_func_46[19]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [20], input_sha_func_46[20]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [21], input_sha_func_46[21]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [22], input_sha_func_46[22]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [23], input_sha_func_46[23]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [24], input_sha_func_46[24]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [25], input_sha_func_46[25]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [26], input_sha_func_46[26]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [27], input_sha_func_46[27]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [28], input_sha_func_46[28]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [29], input_sha_func_46[29]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [30], input_sha_func_46[30]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [31], input_sha_func_46[31]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [32], input_sha_func_46[32]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [33], input_sha_func_46[33]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [34], input_sha_func_46[34]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [35], input_sha_func_46[35]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [36], input_sha_func_46[36]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [37], input_sha_func_46[37]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [38], input_sha_func_46[38]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [39], input_sha_func_46[39]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [40], input_sha_func_46[40]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [41], input_sha_func_46[41]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [42], input_sha_func_46[42]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [43], input_sha_func_46[43]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [44], input_sha_func_46[44]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [45], input_sha_func_46[45]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [46], input_sha_func_46[46]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [47], input_sha_func_46[47]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [48], input_sha_func_46[48]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [49], input_sha_func_46[49]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [50], input_sha_func_46[50]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [51], input_sha_func_46[51]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [52], input_sha_func_46[52]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [53], input_sha_func_46[53]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [54], input_sha_func_46[54]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [55], input_sha_func_46[55]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [56], input_sha_func_46[56]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [57], input_sha_func_46[57]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [58], input_sha_func_46[58]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [59], input_sha_func_46[59]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [60], input_sha_func_46[60]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [61], input_sha_func_46[61]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [62], input_sha_func_46[62]);
  buf(\xm8051_golden_model_1.input_sha_func_46 [63], input_sha_func_46[63]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [0], input_sha_func_45[0]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [1], input_sha_func_45[1]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [2], input_sha_func_45[2]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [3], input_sha_func_45[3]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [4], input_sha_func_45[4]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [5], input_sha_func_45[5]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [6], input_sha_func_45[6]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [7], input_sha_func_45[7]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [8], input_sha_func_45[8]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [9], input_sha_func_45[9]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [10], input_sha_func_45[10]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [11], input_sha_func_45[11]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [12], input_sha_func_45[12]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [13], input_sha_func_45[13]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [14], input_sha_func_45[14]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [15], input_sha_func_45[15]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [16], input_sha_func_45[16]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [17], input_sha_func_45[17]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [18], input_sha_func_45[18]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [19], input_sha_func_45[19]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [20], input_sha_func_45[20]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [21], input_sha_func_45[21]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [22], input_sha_func_45[22]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [23], input_sha_func_45[23]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [24], input_sha_func_45[24]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [25], input_sha_func_45[25]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [26], input_sha_func_45[26]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [27], input_sha_func_45[27]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [28], input_sha_func_45[28]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [29], input_sha_func_45[29]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [30], input_sha_func_45[30]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [31], input_sha_func_45[31]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [32], input_sha_func_45[32]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [33], input_sha_func_45[33]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [34], input_sha_func_45[34]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [35], input_sha_func_45[35]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [36], input_sha_func_45[36]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [37], input_sha_func_45[37]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [38], input_sha_func_45[38]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [39], input_sha_func_45[39]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [40], input_sha_func_45[40]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [41], input_sha_func_45[41]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [42], input_sha_func_45[42]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [43], input_sha_func_45[43]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [44], input_sha_func_45[44]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [45], input_sha_func_45[45]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [46], input_sha_func_45[46]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [47], input_sha_func_45[47]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [48], input_sha_func_45[48]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [49], input_sha_func_45[49]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [50], input_sha_func_45[50]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [51], input_sha_func_45[51]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [52], input_sha_func_45[52]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [53], input_sha_func_45[53]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [54], input_sha_func_45[54]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [55], input_sha_func_45[55]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [56], input_sha_func_45[56]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [57], input_sha_func_45[57]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [58], input_sha_func_45[58]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [59], input_sha_func_45[59]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [60], input_sha_func_45[60]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [61], input_sha_func_45[61]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [62], input_sha_func_45[62]);
  buf(\xm8051_golden_model_1.input_sha_func_45 [63], input_sha_func_45[63]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [0], input_sha_func_44[0]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [1], input_sha_func_44[1]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [2], input_sha_func_44[2]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [3], input_sha_func_44[3]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [4], input_sha_func_44[4]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [5], input_sha_func_44[5]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [6], input_sha_func_44[6]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [7], input_sha_func_44[7]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [8], input_sha_func_44[8]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [9], input_sha_func_44[9]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [10], input_sha_func_44[10]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [11], input_sha_func_44[11]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [12], input_sha_func_44[12]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [13], input_sha_func_44[13]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [14], input_sha_func_44[14]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [15], input_sha_func_44[15]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [16], input_sha_func_44[16]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [17], input_sha_func_44[17]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [18], input_sha_func_44[18]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [19], input_sha_func_44[19]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [20], input_sha_func_44[20]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [21], input_sha_func_44[21]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [22], input_sha_func_44[22]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [23], input_sha_func_44[23]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [24], input_sha_func_44[24]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [25], input_sha_func_44[25]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [26], input_sha_func_44[26]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [27], input_sha_func_44[27]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [28], input_sha_func_44[28]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [29], input_sha_func_44[29]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [30], input_sha_func_44[30]);
  buf(\xm8051_golden_model_1.input_sha_func_44 [31], input_sha_func_44[31]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [0], input_sha_func_43[0]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [1], input_sha_func_43[1]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [2], input_sha_func_43[2]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [3], input_sha_func_43[3]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [4], input_sha_func_43[4]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [5], input_sha_func_43[5]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [6], input_sha_func_43[6]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [7], input_sha_func_43[7]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [8], input_sha_func_43[8]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [9], input_sha_func_43[9]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [10], input_sha_func_43[10]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [11], input_sha_func_43[11]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [12], input_sha_func_43[12]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [13], input_sha_func_43[13]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [14], input_sha_func_43[14]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [15], input_sha_func_43[15]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [16], input_sha_func_43[16]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [17], input_sha_func_43[17]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [18], input_sha_func_43[18]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [19], input_sha_func_43[19]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [20], input_sha_func_43[20]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [21], input_sha_func_43[21]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [22], input_sha_func_43[22]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [23], input_sha_func_43[23]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [24], input_sha_func_43[24]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [25], input_sha_func_43[25]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [26], input_sha_func_43[26]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [27], input_sha_func_43[27]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [28], input_sha_func_43[28]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [29], input_sha_func_43[29]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [30], input_sha_func_43[30]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [31], input_sha_func_43[31]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [32], input_sha_func_43[32]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [33], input_sha_func_43[33]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [34], input_sha_func_43[34]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [35], input_sha_func_43[35]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [36], input_sha_func_43[36]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [37], input_sha_func_43[37]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [38], input_sha_func_43[38]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [39], input_sha_func_43[39]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [40], input_sha_func_43[40]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [41], input_sha_func_43[41]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [42], input_sha_func_43[42]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [43], input_sha_func_43[43]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [44], input_sha_func_43[44]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [45], input_sha_func_43[45]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [46], input_sha_func_43[46]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [47], input_sha_func_43[47]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [48], input_sha_func_43[48]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [49], input_sha_func_43[49]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [50], input_sha_func_43[50]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [51], input_sha_func_43[51]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [52], input_sha_func_43[52]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [53], input_sha_func_43[53]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [54], input_sha_func_43[54]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [55], input_sha_func_43[55]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [56], input_sha_func_43[56]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [57], input_sha_func_43[57]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [58], input_sha_func_43[58]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [59], input_sha_func_43[59]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [60], input_sha_func_43[60]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [61], input_sha_func_43[61]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [62], input_sha_func_43[62]);
  buf(\xm8051_golden_model_1.input_sha_func_43 [63], input_sha_func_43[63]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [0], input_sha_func_42[0]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [1], input_sha_func_42[1]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [2], input_sha_func_42[2]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [3], input_sha_func_42[3]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [4], input_sha_func_42[4]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [5], input_sha_func_42[5]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [6], input_sha_func_42[6]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [7], input_sha_func_42[7]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [8], input_sha_func_42[8]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [9], input_sha_func_42[9]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [10], input_sha_func_42[10]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [11], input_sha_func_42[11]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [12], input_sha_func_42[12]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [13], input_sha_func_42[13]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [14], input_sha_func_42[14]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [15], input_sha_func_42[15]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [16], input_sha_func_42[16]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [17], input_sha_func_42[17]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [18], input_sha_func_42[18]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [19], input_sha_func_42[19]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [20], input_sha_func_42[20]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [21], input_sha_func_42[21]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [22], input_sha_func_42[22]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [23], input_sha_func_42[23]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [24], input_sha_func_42[24]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [25], input_sha_func_42[25]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [26], input_sha_func_42[26]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [27], input_sha_func_42[27]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [28], input_sha_func_42[28]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [29], input_sha_func_42[29]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [30], input_sha_func_42[30]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [31], input_sha_func_42[31]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [32], input_sha_func_42[32]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [33], input_sha_func_42[33]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [34], input_sha_func_42[34]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [35], input_sha_func_42[35]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [36], input_sha_func_42[36]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [37], input_sha_func_42[37]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [38], input_sha_func_42[38]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [39], input_sha_func_42[39]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [40], input_sha_func_42[40]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [41], input_sha_func_42[41]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [42], input_sha_func_42[42]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [43], input_sha_func_42[43]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [44], input_sha_func_42[44]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [45], input_sha_func_42[45]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [46], input_sha_func_42[46]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [47], input_sha_func_42[47]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [48], input_sha_func_42[48]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [49], input_sha_func_42[49]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [50], input_sha_func_42[50]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [51], input_sha_func_42[51]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [52], input_sha_func_42[52]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [53], input_sha_func_42[53]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [54], input_sha_func_42[54]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [55], input_sha_func_42[55]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [56], input_sha_func_42[56]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [57], input_sha_func_42[57]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [58], input_sha_func_42[58]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [59], input_sha_func_42[59]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [60], input_sha_func_42[60]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [61], input_sha_func_42[61]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [62], input_sha_func_42[62]);
  buf(\xm8051_golden_model_1.input_sha_func_42 [63], input_sha_func_42[63]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [0], input_sha_func_41[0]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [1], input_sha_func_41[1]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [2], input_sha_func_41[2]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [3], input_sha_func_41[3]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [4], input_sha_func_41[4]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [5], input_sha_func_41[5]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [6], input_sha_func_41[6]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [7], input_sha_func_41[7]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [8], input_sha_func_41[8]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [9], input_sha_func_41[9]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [10], input_sha_func_41[10]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [11], input_sha_func_41[11]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [12], input_sha_func_41[12]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [13], input_sha_func_41[13]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [14], input_sha_func_41[14]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [15], input_sha_func_41[15]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [16], input_sha_func_41[16]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [17], input_sha_func_41[17]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [18], input_sha_func_41[18]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [19], input_sha_func_41[19]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [20], input_sha_func_41[20]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [21], input_sha_func_41[21]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [22], input_sha_func_41[22]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [23], input_sha_func_41[23]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [24], input_sha_func_41[24]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [25], input_sha_func_41[25]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [26], input_sha_func_41[26]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [27], input_sha_func_41[27]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [28], input_sha_func_41[28]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [29], input_sha_func_41[29]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [30], input_sha_func_41[30]);
  buf(\xm8051_golden_model_1.input_sha_func_41 [31], input_sha_func_41[31]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.data_in [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.data_in [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.data_in [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.data_in [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.data_in [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.data_in [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.data_in [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.data_in [7], proc_data_in[7]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.addr , proc_addr[0]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [0], input_sha_func_40[0]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [1], input_sha_func_40[1]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [2], input_sha_func_40[2]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [3], input_sha_func_40[3]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [4], input_sha_func_40[4]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [5], input_sha_func_40[5]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [6], input_sha_func_40[6]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [7], input_sha_func_40[7]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [8], input_sha_func_40[8]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [9], input_sha_func_40[9]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [10], input_sha_func_40[10]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [11], input_sha_func_40[11]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [12], input_sha_func_40[12]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [13], input_sha_func_40[13]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [14], input_sha_func_40[14]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [15], input_sha_func_40[15]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [16], input_sha_func_40[16]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [17], input_sha_func_40[17]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [18], input_sha_func_40[18]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [19], input_sha_func_40[19]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [20], input_sha_func_40[20]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [21], input_sha_func_40[21]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [22], input_sha_func_40[22]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [23], input_sha_func_40[23]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [24], input_sha_func_40[24]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [25], input_sha_func_40[25]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [26], input_sha_func_40[26]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [27], input_sha_func_40[27]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [28], input_sha_func_40[28]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [29], input_sha_func_40[29]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [30], input_sha_func_40[30]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [31], input_sha_func_40[31]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [32], input_sha_func_40[32]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [33], input_sha_func_40[33]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [34], input_sha_func_40[34]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [35], input_sha_func_40[35]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [36], input_sha_func_40[36]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [37], input_sha_func_40[37]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [38], input_sha_func_40[38]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [39], input_sha_func_40[39]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [40], input_sha_func_40[40]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [41], input_sha_func_40[41]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [42], input_sha_func_40[42]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [43], input_sha_func_40[43]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [44], input_sha_func_40[44]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [45], input_sha_func_40[45]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [46], input_sha_func_40[46]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [47], input_sha_func_40[47]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [48], input_sha_func_40[48]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [49], input_sha_func_40[49]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [50], input_sha_func_40[50]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [51], input_sha_func_40[51]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [52], input_sha_func_40[52]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [53], input_sha_func_40[53]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [54], input_sha_func_40[54]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [55], input_sha_func_40[55]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [56], input_sha_func_40[56]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [57], input_sha_func_40[57]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [58], input_sha_func_40[58]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [59], input_sha_func_40[59]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [60], input_sha_func_40[60]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [61], input_sha_func_40[61]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [62], input_sha_func_40[62]);
  buf(\xm8051_golden_model_1.input_sha_func_40 [63], input_sha_func_40[63]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.rst , rst);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_opaddr_i.clk , clk);
  buf(\xm8051_golden_model_1.input_sha_func_39 [0], input_sha_func_39[0]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [1], input_sha_func_39[1]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [2], input_sha_func_39[2]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [3], input_sha_func_39[3]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [4], input_sha_func_39[4]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [5], input_sha_func_39[5]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [6], input_sha_func_39[6]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [7], input_sha_func_39[7]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [8], input_sha_func_39[8]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [9], input_sha_func_39[9]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [10], input_sha_func_39[10]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [11], input_sha_func_39[11]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [12], input_sha_func_39[12]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [13], input_sha_func_39[13]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [14], input_sha_func_39[14]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [15], input_sha_func_39[15]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [16], input_sha_func_39[16]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [17], input_sha_func_39[17]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [18], input_sha_func_39[18]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [19], input_sha_func_39[19]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [20], input_sha_func_39[20]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [21], input_sha_func_39[21]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [22], input_sha_func_39[22]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [23], input_sha_func_39[23]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [24], input_sha_func_39[24]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [25], input_sha_func_39[25]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [26], input_sha_func_39[26]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [27], input_sha_func_39[27]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [28], input_sha_func_39[28]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [29], input_sha_func_39[29]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [30], input_sha_func_39[30]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [31], input_sha_func_39[31]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [32], input_sha_func_39[32]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [33], input_sha_func_39[33]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [34], input_sha_func_39[34]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [35], input_sha_func_39[35]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [36], input_sha_func_39[36]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [37], input_sha_func_39[37]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [38], input_sha_func_39[38]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [39], input_sha_func_39[39]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [40], input_sha_func_39[40]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [41], input_sha_func_39[41]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [42], input_sha_func_39[42]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [43], input_sha_func_39[43]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [44], input_sha_func_39[44]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [45], input_sha_func_39[45]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [46], input_sha_func_39[46]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [47], input_sha_func_39[47]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [48], input_sha_func_39[48]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [49], input_sha_func_39[49]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [50], input_sha_func_39[50]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [51], input_sha_func_39[51]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [52], input_sha_func_39[52]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [53], input_sha_func_39[53]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [54], input_sha_func_39[54]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [55], input_sha_func_39[55]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [56], input_sha_func_39[56]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [57], input_sha_func_39[57]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [58], input_sha_func_39[58]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [59], input_sha_func_39[59]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [60], input_sha_func_39[60]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [61], input_sha_func_39[61]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [62], input_sha_func_39[62]);
  buf(\xm8051_golden_model_1.input_sha_func_39 [63], input_sha_func_39[63]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [0], input_aes_func_38[0]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [1], input_aes_func_38[1]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [2], input_aes_func_38[2]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [3], input_aes_func_38[3]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [4], input_aes_func_38[4]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [5], input_aes_func_38[5]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [6], input_aes_func_38[6]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [7], input_aes_func_38[7]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [8], input_aes_func_38[8]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [9], input_aes_func_38[9]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [10], input_aes_func_38[10]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [11], input_aes_func_38[11]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [12], input_aes_func_38[12]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [13], input_aes_func_38[13]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [14], input_aes_func_38[14]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [15], input_aes_func_38[15]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [16], input_aes_func_38[16]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [17], input_aes_func_38[17]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [18], input_aes_func_38[18]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [19], input_aes_func_38[19]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [20], input_aes_func_38[20]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [21], input_aes_func_38[21]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [22], input_aes_func_38[22]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [23], input_aes_func_38[23]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [24], input_aes_func_38[24]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [25], input_aes_func_38[25]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [26], input_aes_func_38[26]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [27], input_aes_func_38[27]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [28], input_aes_func_38[28]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [29], input_aes_func_38[29]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [30], input_aes_func_38[30]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [31], input_aes_func_38[31]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [32], input_aes_func_38[32]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [33], input_aes_func_38[33]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [34], input_aes_func_38[34]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [35], input_aes_func_38[35]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [36], input_aes_func_38[36]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [37], input_aes_func_38[37]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [38], input_aes_func_38[38]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [39], input_aes_func_38[39]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [40], input_aes_func_38[40]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [41], input_aes_func_38[41]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [42], input_aes_func_38[42]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [43], input_aes_func_38[43]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [44], input_aes_func_38[44]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [45], input_aes_func_38[45]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [46], input_aes_func_38[46]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [47], input_aes_func_38[47]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [48], input_aes_func_38[48]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [49], input_aes_func_38[49]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [50], input_aes_func_38[50]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [51], input_aes_func_38[51]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [52], input_aes_func_38[52]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [53], input_aes_func_38[53]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [54], input_aes_func_38[54]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [55], input_aes_func_38[55]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [56], input_aes_func_38[56]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [57], input_aes_func_38[57]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [58], input_aes_func_38[58]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [59], input_aes_func_38[59]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [60], input_aes_func_38[60]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [61], input_aes_func_38[61]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [62], input_aes_func_38[62]);
  buf(\xm8051_golden_model_1.input_aes_func_38 [63], input_aes_func_38[63]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [0], input_aes_func_37[0]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [1], input_aes_func_37[1]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [2], input_aes_func_37[2]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [3], input_aes_func_37[3]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [4], input_aes_func_37[4]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [5], input_aes_func_37[5]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [6], input_aes_func_37[6]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [7], input_aes_func_37[7]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [8], input_aes_func_37[8]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [9], input_aes_func_37[9]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [10], input_aes_func_37[10]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [11], input_aes_func_37[11]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [12], input_aes_func_37[12]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [13], input_aes_func_37[13]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [14], input_aes_func_37[14]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [15], input_aes_func_37[15]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [16], input_aes_func_37[16]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [17], input_aes_func_37[17]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [18], input_aes_func_37[18]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [19], input_aes_func_37[19]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [20], input_aes_func_37[20]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [21], input_aes_func_37[21]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [22], input_aes_func_37[22]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [23], input_aes_func_37[23]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [24], input_aes_func_37[24]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [25], input_aes_func_37[25]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [26], input_aes_func_37[26]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [27], input_aes_func_37[27]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [28], input_aes_func_37[28]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [29], input_aes_func_37[29]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [30], input_aes_func_37[30]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [31], input_aes_func_37[31]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [32], input_aes_func_37[32]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [33], input_aes_func_37[33]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [34], input_aes_func_37[34]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [35], input_aes_func_37[35]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [36], input_aes_func_37[36]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [37], input_aes_func_37[37]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [38], input_aes_func_37[38]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [39], input_aes_func_37[39]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [40], input_aes_func_37[40]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [41], input_aes_func_37[41]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [42], input_aes_func_37[42]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [43], input_aes_func_37[43]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [44], input_aes_func_37[44]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [45], input_aes_func_37[45]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [46], input_aes_func_37[46]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [47], input_aes_func_37[47]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [48], input_aes_func_37[48]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [49], input_aes_func_37[49]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [50], input_aes_func_37[50]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [51], input_aes_func_37[51]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [52], input_aes_func_37[52]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [53], input_aes_func_37[53]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [54], input_aes_func_37[54]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [55], input_aes_func_37[55]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [56], input_aes_func_37[56]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [57], input_aes_func_37[57]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [58], input_aes_func_37[58]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [59], input_aes_func_37[59]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [60], input_aes_func_37[60]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [61], input_aes_func_37[61]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [62], input_aes_func_37[62]);
  buf(\xm8051_golden_model_1.input_aes_func_37 [63], input_aes_func_37[63]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [0], input_sha_func_36[0]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [1], input_sha_func_36[1]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [2], input_sha_func_36[2]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [3], input_sha_func_36[3]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [4], input_sha_func_36[4]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [5], input_sha_func_36[5]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [6], input_sha_func_36[6]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [7], input_sha_func_36[7]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [8], input_sha_func_36[8]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [9], input_sha_func_36[9]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [10], input_sha_func_36[10]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [11], input_sha_func_36[11]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [12], input_sha_func_36[12]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [13], input_sha_func_36[13]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [14], input_sha_func_36[14]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [15], input_sha_func_36[15]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [16], input_sha_func_36[16]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [17], input_sha_func_36[17]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [18], input_sha_func_36[18]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [19], input_sha_func_36[19]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [20], input_sha_func_36[20]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [21], input_sha_func_36[21]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [22], input_sha_func_36[22]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [23], input_sha_func_36[23]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [24], input_sha_func_36[24]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [25], input_sha_func_36[25]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [26], input_sha_func_36[26]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [27], input_sha_func_36[27]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [28], input_sha_func_36[28]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [29], input_sha_func_36[29]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [30], input_sha_func_36[30]);
  buf(\xm8051_golden_model_1.input_sha_func_36 [31], input_sha_func_36[31]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [0], input_sha_func_35[0]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [1], input_sha_func_35[1]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [2], input_sha_func_35[2]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [3], input_sha_func_35[3]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [4], input_sha_func_35[4]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [5], input_sha_func_35[5]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [6], input_sha_func_35[6]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [7], input_sha_func_35[7]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [8], input_sha_func_35[8]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [9], input_sha_func_35[9]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [10], input_sha_func_35[10]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [11], input_sha_func_35[11]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [12], input_sha_func_35[12]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [13], input_sha_func_35[13]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [14], input_sha_func_35[14]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [15], input_sha_func_35[15]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [16], input_sha_func_35[16]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [17], input_sha_func_35[17]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [18], input_sha_func_35[18]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [19], input_sha_func_35[19]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [20], input_sha_func_35[20]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [21], input_sha_func_35[21]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [22], input_sha_func_35[22]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [23], input_sha_func_35[23]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [24], input_sha_func_35[24]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [25], input_sha_func_35[25]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [26], input_sha_func_35[26]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [27], input_sha_func_35[27]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [28], input_sha_func_35[28]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [29], input_sha_func_35[29]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [30], input_sha_func_35[30]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [31], input_sha_func_35[31]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [32], input_sha_func_35[32]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [33], input_sha_func_35[33]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [34], input_sha_func_35[34]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [35], input_sha_func_35[35]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [36], input_sha_func_35[36]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [37], input_sha_func_35[37]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [38], input_sha_func_35[38]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [39], input_sha_func_35[39]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [40], input_sha_func_35[40]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [41], input_sha_func_35[41]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [42], input_sha_func_35[42]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [43], input_sha_func_35[43]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [44], input_sha_func_35[44]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [45], input_sha_func_35[45]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [46], input_sha_func_35[46]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [47], input_sha_func_35[47]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [48], input_sha_func_35[48]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [49], input_sha_func_35[49]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [50], input_sha_func_35[50]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [51], input_sha_func_35[51]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [52], input_sha_func_35[52]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [53], input_sha_func_35[53]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [54], input_sha_func_35[54]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [55], input_sha_func_35[55]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [56], input_sha_func_35[56]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [57], input_sha_func_35[57]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [58], input_sha_func_35[58]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [59], input_sha_func_35[59]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [60], input_sha_func_35[60]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [61], input_sha_func_35[61]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [62], input_sha_func_35[62]);
  buf(\xm8051_golden_model_1.input_sha_func_35 [63], input_sha_func_35[63]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [0], input_sha_func_34[0]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [1], input_sha_func_34[1]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [2], input_sha_func_34[2]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [3], input_sha_func_34[3]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [4], input_sha_func_34[4]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [5], input_sha_func_34[5]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [6], input_sha_func_34[6]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [7], input_sha_func_34[7]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [8], input_sha_func_34[8]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [9], input_sha_func_34[9]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [10], input_sha_func_34[10]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [11], input_sha_func_34[11]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [12], input_sha_func_34[12]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [13], input_sha_func_34[13]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [14], input_sha_func_34[14]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [15], input_sha_func_34[15]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [16], input_sha_func_34[16]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [17], input_sha_func_34[17]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [18], input_sha_func_34[18]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [19], input_sha_func_34[19]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [20], input_sha_func_34[20]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [21], input_sha_func_34[21]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [22], input_sha_func_34[22]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [23], input_sha_func_34[23]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [24], input_sha_func_34[24]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [25], input_sha_func_34[25]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [26], input_sha_func_34[26]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [27], input_sha_func_34[27]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [28], input_sha_func_34[28]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [29], input_sha_func_34[29]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [30], input_sha_func_34[30]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [31], input_sha_func_34[31]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [32], input_sha_func_34[32]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [33], input_sha_func_34[33]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [34], input_sha_func_34[34]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [35], input_sha_func_34[35]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [36], input_sha_func_34[36]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [37], input_sha_func_34[37]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [38], input_sha_func_34[38]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [39], input_sha_func_34[39]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [40], input_sha_func_34[40]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [41], input_sha_func_34[41]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [42], input_sha_func_34[42]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [43], input_sha_func_34[43]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [44], input_sha_func_34[44]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [45], input_sha_func_34[45]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [46], input_sha_func_34[46]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [47], input_sha_func_34[47]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [48], input_sha_func_34[48]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [49], input_sha_func_34[49]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [50], input_sha_func_34[50]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [51], input_sha_func_34[51]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [52], input_sha_func_34[52]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [53], input_sha_func_34[53]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [54], input_sha_func_34[54]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [55], input_sha_func_34[55]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [56], input_sha_func_34[56]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [57], input_sha_func_34[57]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [58], input_sha_func_34[58]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [59], input_sha_func_34[59]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [60], input_sha_func_34[60]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [61], input_sha_func_34[61]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [62], input_sha_func_34[62]);
  buf(\xm8051_golden_model_1.input_sha_func_34 [63], input_sha_func_34[63]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.data_in [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.data_in [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.data_in [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.data_in [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.data_in [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.data_in [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.data_in [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.data_in [7], proc_data_in[7]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.addr , proc_addr[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.rst , rst);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.clk , clk);
  buf(\xm8051_golden_model_1.input_sha_func_33 [0], input_sha_func_33[0]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [1], input_sha_func_33[1]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [2], input_sha_func_33[2]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [3], input_sha_func_33[3]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [4], input_sha_func_33[4]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [5], input_sha_func_33[5]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [6], input_sha_func_33[6]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [7], input_sha_func_33[7]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [8], input_sha_func_33[8]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [9], input_sha_func_33[9]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [10], input_sha_func_33[10]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [11], input_sha_func_33[11]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [12], input_sha_func_33[12]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [13], input_sha_func_33[13]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [14], input_sha_func_33[14]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [15], input_sha_func_33[15]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [16], input_sha_func_33[16]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [17], input_sha_func_33[17]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [18], input_sha_func_33[18]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [19], input_sha_func_33[19]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [20], input_sha_func_33[20]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [21], input_sha_func_33[21]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [22], input_sha_func_33[22]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [23], input_sha_func_33[23]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [24], input_sha_func_33[24]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [25], input_sha_func_33[25]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [26], input_sha_func_33[26]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [27], input_sha_func_33[27]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [28], input_sha_func_33[28]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [29], input_sha_func_33[29]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [30], input_sha_func_33[30]);
  buf(\xm8051_golden_model_1.input_sha_func_33 [31], input_sha_func_33[31]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [0], input_sha_func_32[0]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [1], input_sha_func_32[1]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [2], input_sha_func_32[2]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [3], input_sha_func_32[3]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [4], input_sha_func_32[4]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [5], input_sha_func_32[5]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [6], input_sha_func_32[6]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [7], input_sha_func_32[7]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [8], input_sha_func_32[8]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [9], input_sha_func_32[9]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [10], input_sha_func_32[10]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [11], input_sha_func_32[11]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [12], input_sha_func_32[12]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [13], input_sha_func_32[13]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [14], input_sha_func_32[14]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [15], input_sha_func_32[15]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [16], input_sha_func_32[16]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [17], input_sha_func_32[17]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [18], input_sha_func_32[18]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [19], input_sha_func_32[19]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [20], input_sha_func_32[20]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [21], input_sha_func_32[21]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [22], input_sha_func_32[22]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [23], input_sha_func_32[23]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [24], input_sha_func_32[24]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [25], input_sha_func_32[25]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [26], input_sha_func_32[26]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [27], input_sha_func_32[27]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [28], input_sha_func_32[28]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [29], input_sha_func_32[29]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [30], input_sha_func_32[30]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [31], input_sha_func_32[31]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [32], input_sha_func_32[32]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [33], input_sha_func_32[33]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [34], input_sha_func_32[34]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [35], input_sha_func_32[35]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [36], input_sha_func_32[36]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [37], input_sha_func_32[37]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [38], input_sha_func_32[38]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [39], input_sha_func_32[39]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [40], input_sha_func_32[40]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [41], input_sha_func_32[41]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [42], input_sha_func_32[42]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [43], input_sha_func_32[43]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [44], input_sha_func_32[44]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [45], input_sha_func_32[45]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [46], input_sha_func_32[46]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [47], input_sha_func_32[47]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [48], input_sha_func_32[48]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [49], input_sha_func_32[49]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [50], input_sha_func_32[50]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [51], input_sha_func_32[51]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [52], input_sha_func_32[52]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [53], input_sha_func_32[53]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [54], input_sha_func_32[54]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [55], input_sha_func_32[55]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [56], input_sha_func_32[56]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [57], input_sha_func_32[57]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [58], input_sha_func_32[58]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [59], input_sha_func_32[59]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [60], input_sha_func_32[60]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [61], input_sha_func_32[61]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [62], input_sha_func_32[62]);
  buf(\xm8051_golden_model_1.input_sha_func_32 [63], input_sha_func_32[63]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [0], input_sha_func_31[0]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [1], input_sha_func_31[1]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [2], input_sha_func_31[2]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [3], input_sha_func_31[3]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [4], input_sha_func_31[4]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [5], input_sha_func_31[5]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [6], input_sha_func_31[6]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [7], input_sha_func_31[7]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [8], input_sha_func_31[8]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [9], input_sha_func_31[9]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [10], input_sha_func_31[10]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [11], input_sha_func_31[11]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [12], input_sha_func_31[12]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [13], input_sha_func_31[13]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [14], input_sha_func_31[14]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [15], input_sha_func_31[15]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [16], input_sha_func_31[16]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [17], input_sha_func_31[17]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [18], input_sha_func_31[18]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [19], input_sha_func_31[19]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [20], input_sha_func_31[20]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [21], input_sha_func_31[21]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [22], input_sha_func_31[22]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [23], input_sha_func_31[23]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [24], input_sha_func_31[24]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [25], input_sha_func_31[25]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [26], input_sha_func_31[26]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [27], input_sha_func_31[27]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [28], input_sha_func_31[28]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [29], input_sha_func_31[29]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [30], input_sha_func_31[30]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [31], input_sha_func_31[31]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [32], input_sha_func_31[32]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [33], input_sha_func_31[33]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [34], input_sha_func_31[34]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [35], input_sha_func_31[35]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [36], input_sha_func_31[36]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [37], input_sha_func_31[37]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [38], input_sha_func_31[38]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [39], input_sha_func_31[39]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [40], input_sha_func_31[40]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [41], input_sha_func_31[41]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [42], input_sha_func_31[42]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [43], input_sha_func_31[43]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [44], input_sha_func_31[44]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [45], input_sha_func_31[45]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [46], input_sha_func_31[46]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [47], input_sha_func_31[47]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [48], input_sha_func_31[48]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [49], input_sha_func_31[49]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [50], input_sha_func_31[50]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [51], input_sha_func_31[51]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [52], input_sha_func_31[52]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [53], input_sha_func_31[53]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [54], input_sha_func_31[54]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [55], input_sha_func_31[55]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [56], input_sha_func_31[56]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [57], input_sha_func_31[57]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [58], input_sha_func_31[58]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [59], input_sha_func_31[59]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [60], input_sha_func_31[60]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [61], input_sha_func_31[61]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [62], input_sha_func_31[62]);
  buf(\xm8051_golden_model_1.input_sha_func_31 [63], input_sha_func_31[63]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [0], input_sha_func_30[0]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [1], input_sha_func_30[1]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [2], input_sha_func_30[2]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [3], input_sha_func_30[3]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [4], input_sha_func_30[4]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [5], input_sha_func_30[5]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [6], input_sha_func_30[6]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [7], input_sha_func_30[7]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [8], input_sha_func_30[8]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [9], input_sha_func_30[9]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [10], input_sha_func_30[10]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [11], input_sha_func_30[11]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [12], input_sha_func_30[12]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [13], input_sha_func_30[13]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [14], input_sha_func_30[14]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [15], input_sha_func_30[15]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [16], input_sha_func_30[16]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [17], input_sha_func_30[17]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [18], input_sha_func_30[18]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [19], input_sha_func_30[19]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [20], input_sha_func_30[20]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [21], input_sha_func_30[21]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [22], input_sha_func_30[22]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [23], input_sha_func_30[23]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [24], input_sha_func_30[24]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [25], input_sha_func_30[25]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [26], input_sha_func_30[26]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [27], input_sha_func_30[27]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [28], input_sha_func_30[28]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [29], input_sha_func_30[29]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [30], input_sha_func_30[30]);
  buf(\xm8051_golden_model_1.input_sha_func_30 [31], input_sha_func_30[31]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [0], input_sha_func_29[0]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [1], input_sha_func_29[1]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [2], input_sha_func_29[2]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [3], input_sha_func_29[3]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [4], input_sha_func_29[4]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [5], input_sha_func_29[5]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [6], input_sha_func_29[6]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [7], input_sha_func_29[7]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [8], input_sha_func_29[8]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [9], input_sha_func_29[9]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [10], input_sha_func_29[10]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [11], input_sha_func_29[11]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [12], input_sha_func_29[12]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [13], input_sha_func_29[13]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [14], input_sha_func_29[14]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [15], input_sha_func_29[15]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [16], input_sha_func_29[16]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [17], input_sha_func_29[17]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [18], input_sha_func_29[18]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [19], input_sha_func_29[19]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [20], input_sha_func_29[20]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [21], input_sha_func_29[21]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [22], input_sha_func_29[22]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [23], input_sha_func_29[23]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [24], input_sha_func_29[24]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [25], input_sha_func_29[25]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [26], input_sha_func_29[26]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [27], input_sha_func_29[27]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [28], input_sha_func_29[28]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [29], input_sha_func_29[29]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [30], input_sha_func_29[30]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [31], input_sha_func_29[31]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [32], input_sha_func_29[32]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [33], input_sha_func_29[33]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [34], input_sha_func_29[34]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [35], input_sha_func_29[35]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [36], input_sha_func_29[36]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [37], input_sha_func_29[37]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [38], input_sha_func_29[38]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [39], input_sha_func_29[39]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [40], input_sha_func_29[40]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [41], input_sha_func_29[41]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [42], input_sha_func_29[42]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [43], input_sha_func_29[43]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [44], input_sha_func_29[44]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [45], input_sha_func_29[45]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [46], input_sha_func_29[46]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [47], input_sha_func_29[47]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [48], input_sha_func_29[48]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [49], input_sha_func_29[49]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [50], input_sha_func_29[50]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [51], input_sha_func_29[51]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [52], input_sha_func_29[52]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [53], input_sha_func_29[53]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [54], input_sha_func_29[54]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [55], input_sha_func_29[55]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [56], input_sha_func_29[56]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [57], input_sha_func_29[57]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [58], input_sha_func_29[58]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [59], input_sha_func_29[59]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [60], input_sha_func_29[60]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [61], input_sha_func_29[61]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [62], input_sha_func_29[62]);
  buf(\xm8051_golden_model_1.input_sha_func_29 [63], input_sha_func_29[63]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [0], input_sha_func_28[0]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [1], input_sha_func_28[1]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [2], input_sha_func_28[2]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [3], input_sha_func_28[3]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [4], input_sha_func_28[4]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [5], input_sha_func_28[5]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [6], input_sha_func_28[6]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [7], input_sha_func_28[7]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [8], input_sha_func_28[8]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [9], input_sha_func_28[9]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [10], input_sha_func_28[10]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [11], input_sha_func_28[11]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [12], input_sha_func_28[12]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [13], input_sha_func_28[13]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [14], input_sha_func_28[14]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [15], input_sha_func_28[15]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [16], input_sha_func_28[16]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [17], input_sha_func_28[17]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [18], input_sha_func_28[18]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [19], input_sha_func_28[19]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [20], input_sha_func_28[20]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [21], input_sha_func_28[21]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [22], input_sha_func_28[22]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [23], input_sha_func_28[23]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [24], input_sha_func_28[24]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [25], input_sha_func_28[25]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [26], input_sha_func_28[26]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [27], input_sha_func_28[27]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [28], input_sha_func_28[28]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [29], input_sha_func_28[29]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [30], input_sha_func_28[30]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [31], input_sha_func_28[31]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [32], input_sha_func_28[32]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [33], input_sha_func_28[33]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [34], input_sha_func_28[34]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [35], input_sha_func_28[35]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [36], input_sha_func_28[36]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [37], input_sha_func_28[37]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [38], input_sha_func_28[38]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [39], input_sha_func_28[39]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [40], input_sha_func_28[40]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [41], input_sha_func_28[41]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [42], input_sha_func_28[42]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [43], input_sha_func_28[43]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [44], input_sha_func_28[44]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [45], input_sha_func_28[45]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [46], input_sha_func_28[46]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [47], input_sha_func_28[47]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [48], input_sha_func_28[48]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [49], input_sha_func_28[49]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [50], input_sha_func_28[50]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [51], input_sha_func_28[51]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [52], input_sha_func_28[52]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [53], input_sha_func_28[53]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [54], input_sha_func_28[54]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [55], input_sha_func_28[55]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [56], input_sha_func_28[56]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [57], input_sha_func_28[57]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [58], input_sha_func_28[58]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [59], input_sha_func_28[59]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [60], input_sha_func_28[60]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [61], input_sha_func_28[61]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [62], input_sha_func_28[62]);
  buf(\xm8051_golden_model_1.input_sha_func_28 [63], input_sha_func_28[63]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [0], input_sha_func_27[0]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [1], input_sha_func_27[1]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [2], input_sha_func_27[2]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [3], input_sha_func_27[3]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [4], input_sha_func_27[4]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [5], input_sha_func_27[5]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [6], input_sha_func_27[6]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [7], input_sha_func_27[7]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [8], input_sha_func_27[8]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [9], input_sha_func_27[9]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [10], input_sha_func_27[10]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [11], input_sha_func_27[11]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [12], input_sha_func_27[12]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [13], input_sha_func_27[13]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [14], input_sha_func_27[14]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [15], input_sha_func_27[15]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [16], input_sha_func_27[16]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [17], input_sha_func_27[17]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [18], input_sha_func_27[18]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [19], input_sha_func_27[19]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [20], input_sha_func_27[20]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [21], input_sha_func_27[21]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [22], input_sha_func_27[22]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [23], input_sha_func_27[23]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [24], input_sha_func_27[24]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [25], input_sha_func_27[25]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [26], input_sha_func_27[26]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [27], input_sha_func_27[27]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [28], input_sha_func_27[28]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [29], input_sha_func_27[29]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [30], input_sha_func_27[30]);
  buf(\xm8051_golden_model_1.input_sha_func_27 [31], input_sha_func_27[31]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [0], input_sha_func_26[0]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [1], input_sha_func_26[1]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [2], input_sha_func_26[2]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [3], input_sha_func_26[3]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [4], input_sha_func_26[4]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [5], input_sha_func_26[5]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [6], input_sha_func_26[6]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [7], input_sha_func_26[7]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [8], input_sha_func_26[8]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [9], input_sha_func_26[9]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [10], input_sha_func_26[10]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [11], input_sha_func_26[11]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [12], input_sha_func_26[12]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [13], input_sha_func_26[13]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [14], input_sha_func_26[14]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [15], input_sha_func_26[15]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [16], input_sha_func_26[16]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [17], input_sha_func_26[17]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [18], input_sha_func_26[18]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [19], input_sha_func_26[19]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [20], input_sha_func_26[20]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [21], input_sha_func_26[21]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [22], input_sha_func_26[22]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [23], input_sha_func_26[23]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [24], input_sha_func_26[24]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [25], input_sha_func_26[25]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [26], input_sha_func_26[26]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [27], input_sha_func_26[27]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [28], input_sha_func_26[28]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [29], input_sha_func_26[29]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [30], input_sha_func_26[30]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [31], input_sha_func_26[31]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [32], input_sha_func_26[32]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [33], input_sha_func_26[33]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [34], input_sha_func_26[34]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [35], input_sha_func_26[35]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [36], input_sha_func_26[36]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [37], input_sha_func_26[37]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [38], input_sha_func_26[38]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [39], input_sha_func_26[39]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [40], input_sha_func_26[40]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [41], input_sha_func_26[41]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [42], input_sha_func_26[42]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [43], input_sha_func_26[43]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [44], input_sha_func_26[44]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [45], input_sha_func_26[45]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [46], input_sha_func_26[46]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [47], input_sha_func_26[47]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [48], input_sha_func_26[48]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [49], input_sha_func_26[49]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [50], input_sha_func_26[50]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [51], input_sha_func_26[51]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [52], input_sha_func_26[52]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [53], input_sha_func_26[53]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [54], input_sha_func_26[54]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [55], input_sha_func_26[55]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [56], input_sha_func_26[56]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [57], input_sha_func_26[57]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [58], input_sha_func_26[58]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [59], input_sha_func_26[59]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [60], input_sha_func_26[60]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [61], input_sha_func_26[61]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [62], input_sha_func_26[62]);
  buf(\xm8051_golden_model_1.input_sha_func_26 [63], input_sha_func_26[63]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [0], input_sha_func_25[0]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [1], input_sha_func_25[1]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [2], input_sha_func_25[2]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [3], input_sha_func_25[3]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [4], input_sha_func_25[4]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [5], input_sha_func_25[5]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [6], input_sha_func_25[6]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [7], input_sha_func_25[7]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [8], input_sha_func_25[8]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [9], input_sha_func_25[9]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [10], input_sha_func_25[10]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [11], input_sha_func_25[11]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [12], input_sha_func_25[12]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [13], input_sha_func_25[13]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [14], input_sha_func_25[14]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [15], input_sha_func_25[15]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [16], input_sha_func_25[16]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [17], input_sha_func_25[17]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [18], input_sha_func_25[18]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [19], input_sha_func_25[19]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [20], input_sha_func_25[20]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [21], input_sha_func_25[21]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [22], input_sha_func_25[22]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [23], input_sha_func_25[23]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [24], input_sha_func_25[24]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [25], input_sha_func_25[25]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [26], input_sha_func_25[26]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [27], input_sha_func_25[27]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [28], input_sha_func_25[28]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [29], input_sha_func_25[29]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [30], input_sha_func_25[30]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [31], input_sha_func_25[31]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [32], input_sha_func_25[32]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [33], input_sha_func_25[33]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [34], input_sha_func_25[34]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [35], input_sha_func_25[35]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [36], input_sha_func_25[36]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [37], input_sha_func_25[37]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [38], input_sha_func_25[38]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [39], input_sha_func_25[39]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [40], input_sha_func_25[40]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [41], input_sha_func_25[41]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [42], input_sha_func_25[42]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [43], input_sha_func_25[43]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [44], input_sha_func_25[44]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [45], input_sha_func_25[45]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [46], input_sha_func_25[46]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [47], input_sha_func_25[47]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [48], input_sha_func_25[48]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [49], input_sha_func_25[49]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [50], input_sha_func_25[50]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [51], input_sha_func_25[51]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [52], input_sha_func_25[52]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [53], input_sha_func_25[53]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [54], input_sha_func_25[54]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [55], input_sha_func_25[55]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [56], input_sha_func_25[56]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [57], input_sha_func_25[57]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [58], input_sha_func_25[58]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [59], input_sha_func_25[59]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [60], input_sha_func_25[60]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [61], input_sha_func_25[61]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [62], input_sha_func_25[62]);
  buf(\xm8051_golden_model_1.input_sha_func_25 [63], input_sha_func_25[63]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [0], input_aes_func_24[0]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [1], input_aes_func_24[1]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [2], input_aes_func_24[2]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [3], input_aes_func_24[3]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [4], input_aes_func_24[4]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [5], input_aes_func_24[5]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [6], input_aes_func_24[6]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [7], input_aes_func_24[7]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [8], input_aes_func_24[8]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [9], input_aes_func_24[9]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [10], input_aes_func_24[10]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [11], input_aes_func_24[11]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [12], input_aes_func_24[12]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [13], input_aes_func_24[13]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [14], input_aes_func_24[14]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [15], input_aes_func_24[15]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [16], input_aes_func_24[16]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [17], input_aes_func_24[17]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [18], input_aes_func_24[18]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [19], input_aes_func_24[19]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [20], input_aes_func_24[20]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [21], input_aes_func_24[21]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [22], input_aes_func_24[22]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [23], input_aes_func_24[23]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [24], input_aes_func_24[24]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [25], input_aes_func_24[25]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [26], input_aes_func_24[26]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [27], input_aes_func_24[27]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [28], input_aes_func_24[28]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [29], input_aes_func_24[29]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [30], input_aes_func_24[30]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [31], input_aes_func_24[31]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [32], input_aes_func_24[32]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [33], input_aes_func_24[33]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [34], input_aes_func_24[34]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [35], input_aes_func_24[35]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [36], input_aes_func_24[36]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [37], input_aes_func_24[37]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [38], input_aes_func_24[38]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [39], input_aes_func_24[39]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [40], input_aes_func_24[40]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [41], input_aes_func_24[41]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [42], input_aes_func_24[42]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [43], input_aes_func_24[43]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [44], input_aes_func_24[44]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [45], input_aes_func_24[45]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [46], input_aes_func_24[46]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [47], input_aes_func_24[47]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [48], input_aes_func_24[48]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [49], input_aes_func_24[49]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [50], input_aes_func_24[50]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [51], input_aes_func_24[51]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [52], input_aes_func_24[52]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [53], input_aes_func_24[53]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [54], input_aes_func_24[54]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [55], input_aes_func_24[55]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [56], input_aes_func_24[56]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [57], input_aes_func_24[57]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [58], input_aes_func_24[58]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [59], input_aes_func_24[59]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [60], input_aes_func_24[60]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [61], input_aes_func_24[61]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [62], input_aes_func_24[62]);
  buf(\xm8051_golden_model_1.input_aes_func_24 [63], input_aes_func_24[63]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [0], input_aes_func_23[0]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [1], input_aes_func_23[1]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [2], input_aes_func_23[2]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [3], input_aes_func_23[3]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [4], input_aes_func_23[4]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [5], input_aes_func_23[5]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [6], input_aes_func_23[6]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [7], input_aes_func_23[7]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [8], input_aes_func_23[8]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [9], input_aes_func_23[9]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [10], input_aes_func_23[10]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [11], input_aes_func_23[11]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [12], input_aes_func_23[12]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [13], input_aes_func_23[13]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [14], input_aes_func_23[14]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [15], input_aes_func_23[15]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [16], input_aes_func_23[16]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [17], input_aes_func_23[17]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [18], input_aes_func_23[18]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [19], input_aes_func_23[19]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [20], input_aes_func_23[20]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [21], input_aes_func_23[21]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [22], input_aes_func_23[22]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [23], input_aes_func_23[23]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [24], input_aes_func_23[24]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [25], input_aes_func_23[25]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [26], input_aes_func_23[26]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [27], input_aes_func_23[27]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [28], input_aes_func_23[28]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [29], input_aes_func_23[29]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [30], input_aes_func_23[30]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [31], input_aes_func_23[31]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [32], input_aes_func_23[32]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [33], input_aes_func_23[33]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [34], input_aes_func_23[34]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [35], input_aes_func_23[35]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [36], input_aes_func_23[36]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [37], input_aes_func_23[37]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [38], input_aes_func_23[38]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [39], input_aes_func_23[39]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [40], input_aes_func_23[40]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [41], input_aes_func_23[41]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [42], input_aes_func_23[42]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [43], input_aes_func_23[43]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [44], input_aes_func_23[44]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [45], input_aes_func_23[45]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [46], input_aes_func_23[46]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [47], input_aes_func_23[47]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [48], input_aes_func_23[48]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [49], input_aes_func_23[49]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [50], input_aes_func_23[50]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [51], input_aes_func_23[51]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [52], input_aes_func_23[52]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [53], input_aes_func_23[53]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [54], input_aes_func_23[54]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [55], input_aes_func_23[55]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [56], input_aes_func_23[56]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [57], input_aes_func_23[57]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [58], input_aes_func_23[58]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [59], input_aes_func_23[59]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [60], input_aes_func_23[60]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [61], input_aes_func_23[61]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [62], input_aes_func_23[62]);
  buf(\xm8051_golden_model_1.input_aes_func_23 [63], input_aes_func_23[63]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [0], input_sha_func_22[0]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [1], input_sha_func_22[1]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [2], input_sha_func_22[2]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [3], input_sha_func_22[3]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [4], input_sha_func_22[4]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [5], input_sha_func_22[5]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [6], input_sha_func_22[6]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [7], input_sha_func_22[7]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [8], input_sha_func_22[8]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [9], input_sha_func_22[9]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [10], input_sha_func_22[10]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [11], input_sha_func_22[11]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [12], input_sha_func_22[12]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [13], input_sha_func_22[13]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [14], input_sha_func_22[14]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [15], input_sha_func_22[15]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [16], input_sha_func_22[16]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [17], input_sha_func_22[17]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [18], input_sha_func_22[18]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [19], input_sha_func_22[19]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [20], input_sha_func_22[20]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [21], input_sha_func_22[21]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [22], input_sha_func_22[22]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [23], input_sha_func_22[23]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [24], input_sha_func_22[24]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [25], input_sha_func_22[25]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [26], input_sha_func_22[26]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [27], input_sha_func_22[27]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [28], input_sha_func_22[28]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [29], input_sha_func_22[29]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [30], input_sha_func_22[30]);
  buf(\xm8051_golden_model_1.input_sha_func_22 [31], input_sha_func_22[31]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [0], input_sha_func_21[0]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [1], input_sha_func_21[1]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [2], input_sha_func_21[2]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [3], input_sha_func_21[3]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [4], input_sha_func_21[4]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [5], input_sha_func_21[5]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [6], input_sha_func_21[6]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [7], input_sha_func_21[7]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [8], input_sha_func_21[8]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [9], input_sha_func_21[9]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [10], input_sha_func_21[10]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [11], input_sha_func_21[11]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [12], input_sha_func_21[12]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [13], input_sha_func_21[13]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [14], input_sha_func_21[14]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [15], input_sha_func_21[15]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [16], input_sha_func_21[16]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [17], input_sha_func_21[17]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [18], input_sha_func_21[18]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [19], input_sha_func_21[19]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [20], input_sha_func_21[20]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [21], input_sha_func_21[21]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [22], input_sha_func_21[22]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [23], input_sha_func_21[23]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [24], input_sha_func_21[24]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [25], input_sha_func_21[25]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [26], input_sha_func_21[26]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [27], input_sha_func_21[27]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [28], input_sha_func_21[28]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [29], input_sha_func_21[29]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [30], input_sha_func_21[30]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [31], input_sha_func_21[31]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [32], input_sha_func_21[32]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [33], input_sha_func_21[33]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [34], input_sha_func_21[34]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [35], input_sha_func_21[35]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [36], input_sha_func_21[36]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [37], input_sha_func_21[37]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [38], input_sha_func_21[38]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [39], input_sha_func_21[39]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [40], input_sha_func_21[40]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [41], input_sha_func_21[41]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [42], input_sha_func_21[42]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [43], input_sha_func_21[43]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [44], input_sha_func_21[44]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [45], input_sha_func_21[45]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [46], input_sha_func_21[46]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [47], input_sha_func_21[47]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [48], input_sha_func_21[48]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [49], input_sha_func_21[49]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [50], input_sha_func_21[50]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [51], input_sha_func_21[51]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [52], input_sha_func_21[52]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [53], input_sha_func_21[53]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [54], input_sha_func_21[54]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [55], input_sha_func_21[55]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [56], input_sha_func_21[56]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [57], input_sha_func_21[57]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [58], input_sha_func_21[58]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [59], input_sha_func_21[59]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [60], input_sha_func_21[60]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [61], input_sha_func_21[61]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [62], input_sha_func_21[62]);
  buf(\xm8051_golden_model_1.input_sha_func_21 [63], input_sha_func_21[63]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [0], input_sha_func_20[0]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [1], input_sha_func_20[1]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [2], input_sha_func_20[2]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [3], input_sha_func_20[3]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [4], input_sha_func_20[4]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [5], input_sha_func_20[5]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [6], input_sha_func_20[6]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [7], input_sha_func_20[7]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [8], input_sha_func_20[8]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [9], input_sha_func_20[9]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [10], input_sha_func_20[10]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [11], input_sha_func_20[11]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [12], input_sha_func_20[12]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [13], input_sha_func_20[13]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [14], input_sha_func_20[14]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [15], input_sha_func_20[15]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [16], input_sha_func_20[16]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [17], input_sha_func_20[17]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [18], input_sha_func_20[18]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [19], input_sha_func_20[19]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [20], input_sha_func_20[20]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [21], input_sha_func_20[21]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [22], input_sha_func_20[22]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [23], input_sha_func_20[23]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [24], input_sha_func_20[24]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [25], input_sha_func_20[25]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [26], input_sha_func_20[26]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [27], input_sha_func_20[27]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [28], input_sha_func_20[28]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [29], input_sha_func_20[29]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [30], input_sha_func_20[30]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [31], input_sha_func_20[31]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [32], input_sha_func_20[32]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [33], input_sha_func_20[33]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [34], input_sha_func_20[34]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [35], input_sha_func_20[35]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [36], input_sha_func_20[36]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [37], input_sha_func_20[37]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [38], input_sha_func_20[38]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [39], input_sha_func_20[39]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [40], input_sha_func_20[40]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [41], input_sha_func_20[41]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [42], input_sha_func_20[42]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [43], input_sha_func_20[43]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [44], input_sha_func_20[44]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [45], input_sha_func_20[45]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [46], input_sha_func_20[46]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [47], input_sha_func_20[47]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [48], input_sha_func_20[48]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [49], input_sha_func_20[49]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [50], input_sha_func_20[50]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [51], input_sha_func_20[51]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [52], input_sha_func_20[52]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [53], input_sha_func_20[53]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [54], input_sha_func_20[54]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [55], input_sha_func_20[55]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [56], input_sha_func_20[56]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [57], input_sha_func_20[57]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [58], input_sha_func_20[58]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [59], input_sha_func_20[59]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [60], input_sha_func_20[60]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [61], input_sha_func_20[61]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [62], input_sha_func_20[62]);
  buf(\xm8051_golden_model_1.input_sha_func_20 [63], input_sha_func_20[63]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [0], input_sha_func_19[0]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [1], input_sha_func_19[1]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [2], input_sha_func_19[2]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [3], input_sha_func_19[3]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [4], input_sha_func_19[4]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [5], input_sha_func_19[5]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [6], input_sha_func_19[6]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [7], input_sha_func_19[7]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [8], input_sha_func_19[8]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [9], input_sha_func_19[9]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [10], input_sha_func_19[10]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [11], input_sha_func_19[11]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [12], input_sha_func_19[12]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [13], input_sha_func_19[13]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [14], input_sha_func_19[14]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [15], input_sha_func_19[15]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [16], input_sha_func_19[16]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [17], input_sha_func_19[17]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [18], input_sha_func_19[18]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [19], input_sha_func_19[19]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [20], input_sha_func_19[20]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [21], input_sha_func_19[21]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [22], input_sha_func_19[22]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [23], input_sha_func_19[23]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [24], input_sha_func_19[24]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [25], input_sha_func_19[25]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [26], input_sha_func_19[26]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [27], input_sha_func_19[27]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [28], input_sha_func_19[28]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [29], input_sha_func_19[29]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [30], input_sha_func_19[30]);
  buf(\xm8051_golden_model_1.input_sha_func_19 [31], input_sha_func_19[31]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [0], input_sha_func_18[0]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [1], input_sha_func_18[1]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [2], input_sha_func_18[2]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [3], input_sha_func_18[3]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [4], input_sha_func_18[4]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [5], input_sha_func_18[5]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [6], input_sha_func_18[6]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [7], input_sha_func_18[7]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [8], input_sha_func_18[8]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [9], input_sha_func_18[9]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [10], input_sha_func_18[10]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [11], input_sha_func_18[11]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [12], input_sha_func_18[12]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [13], input_sha_func_18[13]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [14], input_sha_func_18[14]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [15], input_sha_func_18[15]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [16], input_sha_func_18[16]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [17], input_sha_func_18[17]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [18], input_sha_func_18[18]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [19], input_sha_func_18[19]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [20], input_sha_func_18[20]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [21], input_sha_func_18[21]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [22], input_sha_func_18[22]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [23], input_sha_func_18[23]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [24], input_sha_func_18[24]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [25], input_sha_func_18[25]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [26], input_sha_func_18[26]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [27], input_sha_func_18[27]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [28], input_sha_func_18[28]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [29], input_sha_func_18[29]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [30], input_sha_func_18[30]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [31], input_sha_func_18[31]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [32], input_sha_func_18[32]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [33], input_sha_func_18[33]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [34], input_sha_func_18[34]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [35], input_sha_func_18[35]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [36], input_sha_func_18[36]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [37], input_sha_func_18[37]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [38], input_sha_func_18[38]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [39], input_sha_func_18[39]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [40], input_sha_func_18[40]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [41], input_sha_func_18[41]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [42], input_sha_func_18[42]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [43], input_sha_func_18[43]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [44], input_sha_func_18[44]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [45], input_sha_func_18[45]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [46], input_sha_func_18[46]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [47], input_sha_func_18[47]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [48], input_sha_func_18[48]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [49], input_sha_func_18[49]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [50], input_sha_func_18[50]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [51], input_sha_func_18[51]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [52], input_sha_func_18[52]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [53], input_sha_func_18[53]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [54], input_sha_func_18[54]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [55], input_sha_func_18[55]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [56], input_sha_func_18[56]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [57], input_sha_func_18[57]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [58], input_sha_func_18[58]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [59], input_sha_func_18[59]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [60], input_sha_func_18[60]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [61], input_sha_func_18[61]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [62], input_sha_func_18[62]);
  buf(\xm8051_golden_model_1.input_sha_func_18 [63], input_sha_func_18[63]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [0], input_sha_func_17[0]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [1], input_sha_func_17[1]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [2], input_sha_func_17[2]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [3], input_sha_func_17[3]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [4], input_sha_func_17[4]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [5], input_sha_func_17[5]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [6], input_sha_func_17[6]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [7], input_sha_func_17[7]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [8], input_sha_func_17[8]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [9], input_sha_func_17[9]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [10], input_sha_func_17[10]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [11], input_sha_func_17[11]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [12], input_sha_func_17[12]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [13], input_sha_func_17[13]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [14], input_sha_func_17[14]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [15], input_sha_func_17[15]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [16], input_sha_func_17[16]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [17], input_sha_func_17[17]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [18], input_sha_func_17[18]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [19], input_sha_func_17[19]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [20], input_sha_func_17[20]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [21], input_sha_func_17[21]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [22], input_sha_func_17[22]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [23], input_sha_func_17[23]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [24], input_sha_func_17[24]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [25], input_sha_func_17[25]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [26], input_sha_func_17[26]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [27], input_sha_func_17[27]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [28], input_sha_func_17[28]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [29], input_sha_func_17[29]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [30], input_sha_func_17[30]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [31], input_sha_func_17[31]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [32], input_sha_func_17[32]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [33], input_sha_func_17[33]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [34], input_sha_func_17[34]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [35], input_sha_func_17[35]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [36], input_sha_func_17[36]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [37], input_sha_func_17[37]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [38], input_sha_func_17[38]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [39], input_sha_func_17[39]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [40], input_sha_func_17[40]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [41], input_sha_func_17[41]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [42], input_sha_func_17[42]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [43], input_sha_func_17[43]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [44], input_sha_func_17[44]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [45], input_sha_func_17[45]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [46], input_sha_func_17[46]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [47], input_sha_func_17[47]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [48], input_sha_func_17[48]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [49], input_sha_func_17[49]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [50], input_sha_func_17[50]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [51], input_sha_func_17[51]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [52], input_sha_func_17[52]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [53], input_sha_func_17[53]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [54], input_sha_func_17[54]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [55], input_sha_func_17[55]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [56], input_sha_func_17[56]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [57], input_sha_func_17[57]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [58], input_sha_func_17[58]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [59], input_sha_func_17[59]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [60], input_sha_func_17[60]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [61], input_sha_func_17[61]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [62], input_sha_func_17[62]);
  buf(\xm8051_golden_model_1.input_sha_func_17 [63], input_sha_func_17[63]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [0], input_sha_func_16[0]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [1], input_sha_func_16[1]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [2], input_sha_func_16[2]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [3], input_sha_func_16[3]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [4], input_sha_func_16[4]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [5], input_sha_func_16[5]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [6], input_sha_func_16[6]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [7], input_sha_func_16[7]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [8], input_sha_func_16[8]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [9], input_sha_func_16[9]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [10], input_sha_func_16[10]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [11], input_sha_func_16[11]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [12], input_sha_func_16[12]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [13], input_sha_func_16[13]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [14], input_sha_func_16[14]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [15], input_sha_func_16[15]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [16], input_sha_func_16[16]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [17], input_sha_func_16[17]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [18], input_sha_func_16[18]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [19], input_sha_func_16[19]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [20], input_sha_func_16[20]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [21], input_sha_func_16[21]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [22], input_sha_func_16[22]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [23], input_sha_func_16[23]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [24], input_sha_func_16[24]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [25], input_sha_func_16[25]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [26], input_sha_func_16[26]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [27], input_sha_func_16[27]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [28], input_sha_func_16[28]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [29], input_sha_func_16[29]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [30], input_sha_func_16[30]);
  buf(\xm8051_golden_model_1.input_sha_func_16 [31], input_sha_func_16[31]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [0], input_sha_func_15[0]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [1], input_sha_func_15[1]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [2], input_sha_func_15[2]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [3], input_sha_func_15[3]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [4], input_sha_func_15[4]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [5], input_sha_func_15[5]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [6], input_sha_func_15[6]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [7], input_sha_func_15[7]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [8], input_sha_func_15[8]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [9], input_sha_func_15[9]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [10], input_sha_func_15[10]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [11], input_sha_func_15[11]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [12], input_sha_func_15[12]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [13], input_sha_func_15[13]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [14], input_sha_func_15[14]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [15], input_sha_func_15[15]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [16], input_sha_func_15[16]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [17], input_sha_func_15[17]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [18], input_sha_func_15[18]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [19], input_sha_func_15[19]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [20], input_sha_func_15[20]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [21], input_sha_func_15[21]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [22], input_sha_func_15[22]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [23], input_sha_func_15[23]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [24], input_sha_func_15[24]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [25], input_sha_func_15[25]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [26], input_sha_func_15[26]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [27], input_sha_func_15[27]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [28], input_sha_func_15[28]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [29], input_sha_func_15[29]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [30], input_sha_func_15[30]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [31], input_sha_func_15[31]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [32], input_sha_func_15[32]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [33], input_sha_func_15[33]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [34], input_sha_func_15[34]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [35], input_sha_func_15[35]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [36], input_sha_func_15[36]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [37], input_sha_func_15[37]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [38], input_sha_func_15[38]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [39], input_sha_func_15[39]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [40], input_sha_func_15[40]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [41], input_sha_func_15[41]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [42], input_sha_func_15[42]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [43], input_sha_func_15[43]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [44], input_sha_func_15[44]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [45], input_sha_func_15[45]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [46], input_sha_func_15[46]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [47], input_sha_func_15[47]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [48], input_sha_func_15[48]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [49], input_sha_func_15[49]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [50], input_sha_func_15[50]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [51], input_sha_func_15[51]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [52], input_sha_func_15[52]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [53], input_sha_func_15[53]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [54], input_sha_func_15[54]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [55], input_sha_func_15[55]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [56], input_sha_func_15[56]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [57], input_sha_func_15[57]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [58], input_sha_func_15[58]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [59], input_sha_func_15[59]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [60], input_sha_func_15[60]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [61], input_sha_func_15[61]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [62], input_sha_func_15[62]);
  buf(\xm8051_golden_model_1.input_sha_func_15 [63], input_sha_func_15[63]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [0], input_sha_func_14[0]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [1], input_sha_func_14[1]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [2], input_sha_func_14[2]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [3], input_sha_func_14[3]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [4], input_sha_func_14[4]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [5], input_sha_func_14[5]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [6], input_sha_func_14[6]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [7], input_sha_func_14[7]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [8], input_sha_func_14[8]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [9], input_sha_func_14[9]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [10], input_sha_func_14[10]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [11], input_sha_func_14[11]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [12], input_sha_func_14[12]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [13], input_sha_func_14[13]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [14], input_sha_func_14[14]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [15], input_sha_func_14[15]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [16], input_sha_func_14[16]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [17], input_sha_func_14[17]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [18], input_sha_func_14[18]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [19], input_sha_func_14[19]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [20], input_sha_func_14[20]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [21], input_sha_func_14[21]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [22], input_sha_func_14[22]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [23], input_sha_func_14[23]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [24], input_sha_func_14[24]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [25], input_sha_func_14[25]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [26], input_sha_func_14[26]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [27], input_sha_func_14[27]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [28], input_sha_func_14[28]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [29], input_sha_func_14[29]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [30], input_sha_func_14[30]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [31], input_sha_func_14[31]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [32], input_sha_func_14[32]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [33], input_sha_func_14[33]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [34], input_sha_func_14[34]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [35], input_sha_func_14[35]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [36], input_sha_func_14[36]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [37], input_sha_func_14[37]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [38], input_sha_func_14[38]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [39], input_sha_func_14[39]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [40], input_sha_func_14[40]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [41], input_sha_func_14[41]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [42], input_sha_func_14[42]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [43], input_sha_func_14[43]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [44], input_sha_func_14[44]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [45], input_sha_func_14[45]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [46], input_sha_func_14[46]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [47], input_sha_func_14[47]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [48], input_sha_func_14[48]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [49], input_sha_func_14[49]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [50], input_sha_func_14[50]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [51], input_sha_func_14[51]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [52], input_sha_func_14[52]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [53], input_sha_func_14[53]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [54], input_sha_func_14[54]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [55], input_sha_func_14[55]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [56], input_sha_func_14[56]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [57], input_sha_func_14[57]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [58], input_sha_func_14[58]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [59], input_sha_func_14[59]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [60], input_sha_func_14[60]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [61], input_sha_func_14[61]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [62], input_sha_func_14[62]);
  buf(\xm8051_golden_model_1.input_sha_func_14 [63], input_sha_func_14[63]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [0], input_sha_func_13[0]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [1], input_sha_func_13[1]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [2], input_sha_func_13[2]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [3], input_sha_func_13[3]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [4], input_sha_func_13[4]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [5], input_sha_func_13[5]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [6], input_sha_func_13[6]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [7], input_sha_func_13[7]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [8], input_sha_func_13[8]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [9], input_sha_func_13[9]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [10], input_sha_func_13[10]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [11], input_sha_func_13[11]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [12], input_sha_func_13[12]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [13], input_sha_func_13[13]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [14], input_sha_func_13[14]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [15], input_sha_func_13[15]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [16], input_sha_func_13[16]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [17], input_sha_func_13[17]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [18], input_sha_func_13[18]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [19], input_sha_func_13[19]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [20], input_sha_func_13[20]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [21], input_sha_func_13[21]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [22], input_sha_func_13[22]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [23], input_sha_func_13[23]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [24], input_sha_func_13[24]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [25], input_sha_func_13[25]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [26], input_sha_func_13[26]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [27], input_sha_func_13[27]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [28], input_sha_func_13[28]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [29], input_sha_func_13[29]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [30], input_sha_func_13[30]);
  buf(\xm8051_golden_model_1.input_sha_func_13 [31], input_sha_func_13[31]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [0], input_sha_func_12[0]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [1], input_sha_func_12[1]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [2], input_sha_func_12[2]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [3], input_sha_func_12[3]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [4], input_sha_func_12[4]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [5], input_sha_func_12[5]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [6], input_sha_func_12[6]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [7], input_sha_func_12[7]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [8], input_sha_func_12[8]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [9], input_sha_func_12[9]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [10], input_sha_func_12[10]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [11], input_sha_func_12[11]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [12], input_sha_func_12[12]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [13], input_sha_func_12[13]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [14], input_sha_func_12[14]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [15], input_sha_func_12[15]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [16], input_sha_func_12[16]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [17], input_sha_func_12[17]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [18], input_sha_func_12[18]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [19], input_sha_func_12[19]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [20], input_sha_func_12[20]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [21], input_sha_func_12[21]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [22], input_sha_func_12[22]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [23], input_sha_func_12[23]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [24], input_sha_func_12[24]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [25], input_sha_func_12[25]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [26], input_sha_func_12[26]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [27], input_sha_func_12[27]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [28], input_sha_func_12[28]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [29], input_sha_func_12[29]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [30], input_sha_func_12[30]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [31], input_sha_func_12[31]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [32], input_sha_func_12[32]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [33], input_sha_func_12[33]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [34], input_sha_func_12[34]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [35], input_sha_func_12[35]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [36], input_sha_func_12[36]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [37], input_sha_func_12[37]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [38], input_sha_func_12[38]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [39], input_sha_func_12[39]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [40], input_sha_func_12[40]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [41], input_sha_func_12[41]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [42], input_sha_func_12[42]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [43], input_sha_func_12[43]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [44], input_sha_func_12[44]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [45], input_sha_func_12[45]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [46], input_sha_func_12[46]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [47], input_sha_func_12[47]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [48], input_sha_func_12[48]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [49], input_sha_func_12[49]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [50], input_sha_func_12[50]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [51], input_sha_func_12[51]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [52], input_sha_func_12[52]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [53], input_sha_func_12[53]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [54], input_sha_func_12[54]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [55], input_sha_func_12[55]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [56], input_sha_func_12[56]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [57], input_sha_func_12[57]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [58], input_sha_func_12[58]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [59], input_sha_func_12[59]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [60], input_sha_func_12[60]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [61], input_sha_func_12[61]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [62], input_sha_func_12[62]);
  buf(\xm8051_golden_model_1.input_sha_func_12 [63], input_sha_func_12[63]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [0], input_sha_func_11[0]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [1], input_sha_func_11[1]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [2], input_sha_func_11[2]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [3], input_sha_func_11[3]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [4], input_sha_func_11[4]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [5], input_sha_func_11[5]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [6], input_sha_func_11[6]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [7], input_sha_func_11[7]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [8], input_sha_func_11[8]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [9], input_sha_func_11[9]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [10], input_sha_func_11[10]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [11], input_sha_func_11[11]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [12], input_sha_func_11[12]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [13], input_sha_func_11[13]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [14], input_sha_func_11[14]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [15], input_sha_func_11[15]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [16], input_sha_func_11[16]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [17], input_sha_func_11[17]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [18], input_sha_func_11[18]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [19], input_sha_func_11[19]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [20], input_sha_func_11[20]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [21], input_sha_func_11[21]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [22], input_sha_func_11[22]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [23], input_sha_func_11[23]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [24], input_sha_func_11[24]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [25], input_sha_func_11[25]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [26], input_sha_func_11[26]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [27], input_sha_func_11[27]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [28], input_sha_func_11[28]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [29], input_sha_func_11[29]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [30], input_sha_func_11[30]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [31], input_sha_func_11[31]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [32], input_sha_func_11[32]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [33], input_sha_func_11[33]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [34], input_sha_func_11[34]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [35], input_sha_func_11[35]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [36], input_sha_func_11[36]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [37], input_sha_func_11[37]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [38], input_sha_func_11[38]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [39], input_sha_func_11[39]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [40], input_sha_func_11[40]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [41], input_sha_func_11[41]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [42], input_sha_func_11[42]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [43], input_sha_func_11[43]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [44], input_sha_func_11[44]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [45], input_sha_func_11[45]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [46], input_sha_func_11[46]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [47], input_sha_func_11[47]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [48], input_sha_func_11[48]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [49], input_sha_func_11[49]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [50], input_sha_func_11[50]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [51], input_sha_func_11[51]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [52], input_sha_func_11[52]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [53], input_sha_func_11[53]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [54], input_sha_func_11[54]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [55], input_sha_func_11[55]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [56], input_sha_func_11[56]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [57], input_sha_func_11[57]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [58], input_sha_func_11[58]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [59], input_sha_func_11[59]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [60], input_sha_func_11[60]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [61], input_sha_func_11[61]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [62], input_sha_func_11[62]);
  buf(\xm8051_golden_model_1.input_sha_func_11 [63], input_sha_func_11[63]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [0], input_sha_func_10[0]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [1], input_sha_func_10[1]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [2], input_sha_func_10[2]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [3], input_sha_func_10[3]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [4], input_sha_func_10[4]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [5], input_sha_func_10[5]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [6], input_sha_func_10[6]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [7], input_sha_func_10[7]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [8], input_sha_func_10[8]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [9], input_sha_func_10[9]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [10], input_sha_func_10[10]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [11], input_sha_func_10[11]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [12], input_sha_func_10[12]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [13], input_sha_func_10[13]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [14], input_sha_func_10[14]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [15], input_sha_func_10[15]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [16], input_sha_func_10[16]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [17], input_sha_func_10[17]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [18], input_sha_func_10[18]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [19], input_sha_func_10[19]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [20], input_sha_func_10[20]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [21], input_sha_func_10[21]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [22], input_sha_func_10[22]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [23], input_sha_func_10[23]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [24], input_sha_func_10[24]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [25], input_sha_func_10[25]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [26], input_sha_func_10[26]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [27], input_sha_func_10[27]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [28], input_sha_func_10[28]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [29], input_sha_func_10[29]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [30], input_sha_func_10[30]);
  buf(\xm8051_golden_model_1.input_sha_func_10 [31], input_sha_func_10[31]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [0], input_sha_func_9[0]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [1], input_sha_func_9[1]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [2], input_sha_func_9[2]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [3], input_sha_func_9[3]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [4], input_sha_func_9[4]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [5], input_sha_func_9[5]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [6], input_sha_func_9[6]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [7], input_sha_func_9[7]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [8], input_sha_func_9[8]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [9], input_sha_func_9[9]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [10], input_sha_func_9[10]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [11], input_sha_func_9[11]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [12], input_sha_func_9[12]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [13], input_sha_func_9[13]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [14], input_sha_func_9[14]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [15], input_sha_func_9[15]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [16], input_sha_func_9[16]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [17], input_sha_func_9[17]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [18], input_sha_func_9[18]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [19], input_sha_func_9[19]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [20], input_sha_func_9[20]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [21], input_sha_func_9[21]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [22], input_sha_func_9[22]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [23], input_sha_func_9[23]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [24], input_sha_func_9[24]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [25], input_sha_func_9[25]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [26], input_sha_func_9[26]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [27], input_sha_func_9[27]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [28], input_sha_func_9[28]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [29], input_sha_func_9[29]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [30], input_sha_func_9[30]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [31], input_sha_func_9[31]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [32], input_sha_func_9[32]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [33], input_sha_func_9[33]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [34], input_sha_func_9[34]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [35], input_sha_func_9[35]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [36], input_sha_func_9[36]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [37], input_sha_func_9[37]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [38], input_sha_func_9[38]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [39], input_sha_func_9[39]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [40], input_sha_func_9[40]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [41], input_sha_func_9[41]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [42], input_sha_func_9[42]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [43], input_sha_func_9[43]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [44], input_sha_func_9[44]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [45], input_sha_func_9[45]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [46], input_sha_func_9[46]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [47], input_sha_func_9[47]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [48], input_sha_func_9[48]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [49], input_sha_func_9[49]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [50], input_sha_func_9[50]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [51], input_sha_func_9[51]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [52], input_sha_func_9[52]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [53], input_sha_func_9[53]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [54], input_sha_func_9[54]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [55], input_sha_func_9[55]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [56], input_sha_func_9[56]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [57], input_sha_func_9[57]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [58], input_sha_func_9[58]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [59], input_sha_func_9[59]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [60], input_sha_func_9[60]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [61], input_sha_func_9[61]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [62], input_sha_func_9[62]);
  buf(\xm8051_golden_model_1.input_sha_func_9 [63], input_sha_func_9[63]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [0], input_sha_func_8[0]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [1], input_sha_func_8[1]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [2], input_sha_func_8[2]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [3], input_sha_func_8[3]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [4], input_sha_func_8[4]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [5], input_sha_func_8[5]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [6], input_sha_func_8[6]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [7], input_sha_func_8[7]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [8], input_sha_func_8[8]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [9], input_sha_func_8[9]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [10], input_sha_func_8[10]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [11], input_sha_func_8[11]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [12], input_sha_func_8[12]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [13], input_sha_func_8[13]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [14], input_sha_func_8[14]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [15], input_sha_func_8[15]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [16], input_sha_func_8[16]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [17], input_sha_func_8[17]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [18], input_sha_func_8[18]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [19], input_sha_func_8[19]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [20], input_sha_func_8[20]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [21], input_sha_func_8[21]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [22], input_sha_func_8[22]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [23], input_sha_func_8[23]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [24], input_sha_func_8[24]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [25], input_sha_func_8[25]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [26], input_sha_func_8[26]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [27], input_sha_func_8[27]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [28], input_sha_func_8[28]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [29], input_sha_func_8[29]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [30], input_sha_func_8[30]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [31], input_sha_func_8[31]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [32], input_sha_func_8[32]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [33], input_sha_func_8[33]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [34], input_sha_func_8[34]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [35], input_sha_func_8[35]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [36], input_sha_func_8[36]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [37], input_sha_func_8[37]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [38], input_sha_func_8[38]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [39], input_sha_func_8[39]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [40], input_sha_func_8[40]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [41], input_sha_func_8[41]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [42], input_sha_func_8[42]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [43], input_sha_func_8[43]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [44], input_sha_func_8[44]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [45], input_sha_func_8[45]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [46], input_sha_func_8[46]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [47], input_sha_func_8[47]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [48], input_sha_func_8[48]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [49], input_sha_func_8[49]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [50], input_sha_func_8[50]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [51], input_sha_func_8[51]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [52], input_sha_func_8[52]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [53], input_sha_func_8[53]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [54], input_sha_func_8[54]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [55], input_sha_func_8[55]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [56], input_sha_func_8[56]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [57], input_sha_func_8[57]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [58], input_sha_func_8[58]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [59], input_sha_func_8[59]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [60], input_sha_func_8[60]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [61], input_sha_func_8[61]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [62], input_sha_func_8[62]);
  buf(\xm8051_golden_model_1.input_sha_func_8 [63], input_sha_func_8[63]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [0], input_aes_func_7[0]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [1], input_aes_func_7[1]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [2], input_aes_func_7[2]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [3], input_aes_func_7[3]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [4], input_aes_func_7[4]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [5], input_aes_func_7[5]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [6], input_aes_func_7[6]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [7], input_aes_func_7[7]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [8], input_aes_func_7[8]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [9], input_aes_func_7[9]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [10], input_aes_func_7[10]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [11], input_aes_func_7[11]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [12], input_aes_func_7[12]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [13], input_aes_func_7[13]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [14], input_aes_func_7[14]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [15], input_aes_func_7[15]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [16], input_aes_func_7[16]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [17], input_aes_func_7[17]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [18], input_aes_func_7[18]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [19], input_aes_func_7[19]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [20], input_aes_func_7[20]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [21], input_aes_func_7[21]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [22], input_aes_func_7[22]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [23], input_aes_func_7[23]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [24], input_aes_func_7[24]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [25], input_aes_func_7[25]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [26], input_aes_func_7[26]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [27], input_aes_func_7[27]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [28], input_aes_func_7[28]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [29], input_aes_func_7[29]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [30], input_aes_func_7[30]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [31], input_aes_func_7[31]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [32], input_aes_func_7[32]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [33], input_aes_func_7[33]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [34], input_aes_func_7[34]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [35], input_aes_func_7[35]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [36], input_aes_func_7[36]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [37], input_aes_func_7[37]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [38], input_aes_func_7[38]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [39], input_aes_func_7[39]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [40], input_aes_func_7[40]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [41], input_aes_func_7[41]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [42], input_aes_func_7[42]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [43], input_aes_func_7[43]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [44], input_aes_func_7[44]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [45], input_aes_func_7[45]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [46], input_aes_func_7[46]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [47], input_aes_func_7[47]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [48], input_aes_func_7[48]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [49], input_aes_func_7[49]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [50], input_aes_func_7[50]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [51], input_aes_func_7[51]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [52], input_aes_func_7[52]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [53], input_aes_func_7[53]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [54], input_aes_func_7[54]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [55], input_aes_func_7[55]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [56], input_aes_func_7[56]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [57], input_aes_func_7[57]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [58], input_aes_func_7[58]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [59], input_aes_func_7[59]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [60], input_aes_func_7[60]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [61], input_aes_func_7[61]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [62], input_aes_func_7[62]);
  buf(\xm8051_golden_model_1.input_aes_func_7 [63], input_aes_func_7[63]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [0], input_aes_func_6[0]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [1], input_aes_func_6[1]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [2], input_aes_func_6[2]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [3], input_aes_func_6[3]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [4], input_aes_func_6[4]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [5], input_aes_func_6[5]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [6], input_aes_func_6[6]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [7], input_aes_func_6[7]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [8], input_aes_func_6[8]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [9], input_aes_func_6[9]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [10], input_aes_func_6[10]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [11], input_aes_func_6[11]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [12], input_aes_func_6[12]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [13], input_aes_func_6[13]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [14], input_aes_func_6[14]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [15], input_aes_func_6[15]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [16], input_aes_func_6[16]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [17], input_aes_func_6[17]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [18], input_aes_func_6[18]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [19], input_aes_func_6[19]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [20], input_aes_func_6[20]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [21], input_aes_func_6[21]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [22], input_aes_func_6[22]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [23], input_aes_func_6[23]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [24], input_aes_func_6[24]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [25], input_aes_func_6[25]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [26], input_aes_func_6[26]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [27], input_aes_func_6[27]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [28], input_aes_func_6[28]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [29], input_aes_func_6[29]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [30], input_aes_func_6[30]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [31], input_aes_func_6[31]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [32], input_aes_func_6[32]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [33], input_aes_func_6[33]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [34], input_aes_func_6[34]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [35], input_aes_func_6[35]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [36], input_aes_func_6[36]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [37], input_aes_func_6[37]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [38], input_aes_func_6[38]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [39], input_aes_func_6[39]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [40], input_aes_func_6[40]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [41], input_aes_func_6[41]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [42], input_aes_func_6[42]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [43], input_aes_func_6[43]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [44], input_aes_func_6[44]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [45], input_aes_func_6[45]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [46], input_aes_func_6[46]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [47], input_aes_func_6[47]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [48], input_aes_func_6[48]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [49], input_aes_func_6[49]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [50], input_aes_func_6[50]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [51], input_aes_func_6[51]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [52], input_aes_func_6[52]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [53], input_aes_func_6[53]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [54], input_aes_func_6[54]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [55], input_aes_func_6[55]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [56], input_aes_func_6[56]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [57], input_aes_func_6[57]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [58], input_aes_func_6[58]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [59], input_aes_func_6[59]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [60], input_aes_func_6[60]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [61], input_aes_func_6[61]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [62], input_aes_func_6[62]);
  buf(\xm8051_golden_model_1.input_aes_func_6 [63], input_aes_func_6[63]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [0], input_sha_func_5[0]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [1], input_sha_func_5[1]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [2], input_sha_func_5[2]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [3], input_sha_func_5[3]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [4], input_sha_func_5[4]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [5], input_sha_func_5[5]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [6], input_sha_func_5[6]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [7], input_sha_func_5[7]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [8], input_sha_func_5[8]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [9], input_sha_func_5[9]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [10], input_sha_func_5[10]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [11], input_sha_func_5[11]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [12], input_sha_func_5[12]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [13], input_sha_func_5[13]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [14], input_sha_func_5[14]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [15], input_sha_func_5[15]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [16], input_sha_func_5[16]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [17], input_sha_func_5[17]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [18], input_sha_func_5[18]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [19], input_sha_func_5[19]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [20], input_sha_func_5[20]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [21], input_sha_func_5[21]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [22], input_sha_func_5[22]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [23], input_sha_func_5[23]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [24], input_sha_func_5[24]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [25], input_sha_func_5[25]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [26], input_sha_func_5[26]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [27], input_sha_func_5[27]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [28], input_sha_func_5[28]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [29], input_sha_func_5[29]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [30], input_sha_func_5[30]);
  buf(\xm8051_golden_model_1.input_sha_func_5 [31], input_sha_func_5[31]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [0], input_sha_func_4[0]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [1], input_sha_func_4[1]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [2], input_sha_func_4[2]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [3], input_sha_func_4[3]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [4], input_sha_func_4[4]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [5], input_sha_func_4[5]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [6], input_sha_func_4[6]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [7], input_sha_func_4[7]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [8], input_sha_func_4[8]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [9], input_sha_func_4[9]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [10], input_sha_func_4[10]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [11], input_sha_func_4[11]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [12], input_sha_func_4[12]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [13], input_sha_func_4[13]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [14], input_sha_func_4[14]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [15], input_sha_func_4[15]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [16], input_sha_func_4[16]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [17], input_sha_func_4[17]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [18], input_sha_func_4[18]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [19], input_sha_func_4[19]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [20], input_sha_func_4[20]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [21], input_sha_func_4[21]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [22], input_sha_func_4[22]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [23], input_sha_func_4[23]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [24], input_sha_func_4[24]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [25], input_sha_func_4[25]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [26], input_sha_func_4[26]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [27], input_sha_func_4[27]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [28], input_sha_func_4[28]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [29], input_sha_func_4[29]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [30], input_sha_func_4[30]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [31], input_sha_func_4[31]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [32], input_sha_func_4[32]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [33], input_sha_func_4[33]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [34], input_sha_func_4[34]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [35], input_sha_func_4[35]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [36], input_sha_func_4[36]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [37], input_sha_func_4[37]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [38], input_sha_func_4[38]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [39], input_sha_func_4[39]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [40], input_sha_func_4[40]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [41], input_sha_func_4[41]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [42], input_sha_func_4[42]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [43], input_sha_func_4[43]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [44], input_sha_func_4[44]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [45], input_sha_func_4[45]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [46], input_sha_func_4[46]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [47], input_sha_func_4[47]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [48], input_sha_func_4[48]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [49], input_sha_func_4[49]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [50], input_sha_func_4[50]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [51], input_sha_func_4[51]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [52], input_sha_func_4[52]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [53], input_sha_func_4[53]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [54], input_sha_func_4[54]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [55], input_sha_func_4[55]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [56], input_sha_func_4[56]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [57], input_sha_func_4[57]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [58], input_sha_func_4[58]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [59], input_sha_func_4[59]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [60], input_sha_func_4[60]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [61], input_sha_func_4[61]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [62], input_sha_func_4[62]);
  buf(\xm8051_golden_model_1.input_sha_func_4 [63], input_sha_func_4[63]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [0], input_sha_func_3[0]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [1], input_sha_func_3[1]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [2], input_sha_func_3[2]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [3], input_sha_func_3[3]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [4], input_sha_func_3[4]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [5], input_sha_func_3[5]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [6], input_sha_func_3[6]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [7], input_sha_func_3[7]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [8], input_sha_func_3[8]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [9], input_sha_func_3[9]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [10], input_sha_func_3[10]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [11], input_sha_func_3[11]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [12], input_sha_func_3[12]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [13], input_sha_func_3[13]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [14], input_sha_func_3[14]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [15], input_sha_func_3[15]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [16], input_sha_func_3[16]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [17], input_sha_func_3[17]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [18], input_sha_func_3[18]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [19], input_sha_func_3[19]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [20], input_sha_func_3[20]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [21], input_sha_func_3[21]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [22], input_sha_func_3[22]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [23], input_sha_func_3[23]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [24], input_sha_func_3[24]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [25], input_sha_func_3[25]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [26], input_sha_func_3[26]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [27], input_sha_func_3[27]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [28], input_sha_func_3[28]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [29], input_sha_func_3[29]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [30], input_sha_func_3[30]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [31], input_sha_func_3[31]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [32], input_sha_func_3[32]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [33], input_sha_func_3[33]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [34], input_sha_func_3[34]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [35], input_sha_func_3[35]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [36], input_sha_func_3[36]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [37], input_sha_func_3[37]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [38], input_sha_func_3[38]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [39], input_sha_func_3[39]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [40], input_sha_func_3[40]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [41], input_sha_func_3[41]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [42], input_sha_func_3[42]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [43], input_sha_func_3[43]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [44], input_sha_func_3[44]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [45], input_sha_func_3[45]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [46], input_sha_func_3[46]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [47], input_sha_func_3[47]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [48], input_sha_func_3[48]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [49], input_sha_func_3[49]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [50], input_sha_func_3[50]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [51], input_sha_func_3[51]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [52], input_sha_func_3[52]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [53], input_sha_func_3[53]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [54], input_sha_func_3[54]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [55], input_sha_func_3[55]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [56], input_sha_func_3[56]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [57], input_sha_func_3[57]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [58], input_sha_func_3[58]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [59], input_sha_func_3[59]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [60], input_sha_func_3[60]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [61], input_sha_func_3[61]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [62], input_sha_func_3[62]);
  buf(\xm8051_golden_model_1.input_sha_func_3 [63], input_sha_func_3[63]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [0], input_sha_func_2[0]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [1], input_sha_func_2[1]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [2], input_sha_func_2[2]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [3], input_sha_func_2[3]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [4], input_sha_func_2[4]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [5], input_sha_func_2[5]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [6], input_sha_func_2[6]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [7], input_sha_func_2[7]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [8], input_sha_func_2[8]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [9], input_sha_func_2[9]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [10], input_sha_func_2[10]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [11], input_sha_func_2[11]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [12], input_sha_func_2[12]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [13], input_sha_func_2[13]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [14], input_sha_func_2[14]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [15], input_sha_func_2[15]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [16], input_sha_func_2[16]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [17], input_sha_func_2[17]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [18], input_sha_func_2[18]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [19], input_sha_func_2[19]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [20], input_sha_func_2[20]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [21], input_sha_func_2[21]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [22], input_sha_func_2[22]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [23], input_sha_func_2[23]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [24], input_sha_func_2[24]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [25], input_sha_func_2[25]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [26], input_sha_func_2[26]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [27], input_sha_func_2[27]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [28], input_sha_func_2[28]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [29], input_sha_func_2[29]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [30], input_sha_func_2[30]);
  buf(\xm8051_golden_model_1.input_sha_func_2 [31], input_sha_func_2[31]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [0], input_sha_func_1[0]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [1], input_sha_func_1[1]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [2], input_sha_func_1[2]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [3], input_sha_func_1[3]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [4], input_sha_func_1[4]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [5], input_sha_func_1[5]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [6], input_sha_func_1[6]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [7], input_sha_func_1[7]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [8], input_sha_func_1[8]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [9], input_sha_func_1[9]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [10], input_sha_func_1[10]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [11], input_sha_func_1[11]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [12], input_sha_func_1[12]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [13], input_sha_func_1[13]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [14], input_sha_func_1[14]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [15], input_sha_func_1[15]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [16], input_sha_func_1[16]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [17], input_sha_func_1[17]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [18], input_sha_func_1[18]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [19], input_sha_func_1[19]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [20], input_sha_func_1[20]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [21], input_sha_func_1[21]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [22], input_sha_func_1[22]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [23], input_sha_func_1[23]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [24], input_sha_func_1[24]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [25], input_sha_func_1[25]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [26], input_sha_func_1[26]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [27], input_sha_func_1[27]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [28], input_sha_func_1[28]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [29], input_sha_func_1[29]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [30], input_sha_func_1[30]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [31], input_sha_func_1[31]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [32], input_sha_func_1[32]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [33], input_sha_func_1[33]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [34], input_sha_func_1[34]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [35], input_sha_func_1[35]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [36], input_sha_func_1[36]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [37], input_sha_func_1[37]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [38], input_sha_func_1[38]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [39], input_sha_func_1[39]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [40], input_sha_func_1[40]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [41], input_sha_func_1[41]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [42], input_sha_func_1[42]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [43], input_sha_func_1[43]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [44], input_sha_func_1[44]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [45], input_sha_func_1[45]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [46], input_sha_func_1[46]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [47], input_sha_func_1[47]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [48], input_sha_func_1[48]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [49], input_sha_func_1[49]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [50], input_sha_func_1[50]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [51], input_sha_func_1[51]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [52], input_sha_func_1[52]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [53], input_sha_func_1[53]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [54], input_sha_func_1[54]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [55], input_sha_func_1[55]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [56], input_sha_func_1[56]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [57], input_sha_func_1[57]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [58], input_sha_func_1[58]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [59], input_sha_func_1[59]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [60], input_sha_func_1[60]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [61], input_sha_func_1[61]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [62], input_sha_func_1[62]);
  buf(\xm8051_golden_model_1.input_sha_func_1 [63], input_sha_func_1[63]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [0], input_sha_func_0[0]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [1], input_sha_func_0[1]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [2], input_sha_func_0[2]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [3], input_sha_func_0[3]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [4], input_sha_func_0[4]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [5], input_sha_func_0[5]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [6], input_sha_func_0[6]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [7], input_sha_func_0[7]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [8], input_sha_func_0[8]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [9], input_sha_func_0[9]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [10], input_sha_func_0[10]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [11], input_sha_func_0[11]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [12], input_sha_func_0[12]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [13], input_sha_func_0[13]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [14], input_sha_func_0[14]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [15], input_sha_func_0[15]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [16], input_sha_func_0[16]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [17], input_sha_func_0[17]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [18], input_sha_func_0[18]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [19], input_sha_func_0[19]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [20], input_sha_func_0[20]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [21], input_sha_func_0[21]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [22], input_sha_func_0[22]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [23], input_sha_func_0[23]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [24], input_sha_func_0[24]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [25], input_sha_func_0[25]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [26], input_sha_func_0[26]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [27], input_sha_func_0[27]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [28], input_sha_func_0[28]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [29], input_sha_func_0[29]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [30], input_sha_func_0[30]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [31], input_sha_func_0[31]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [32], input_sha_func_0[32]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [33], input_sha_func_0[33]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [34], input_sha_func_0[34]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [35], input_sha_func_0[35]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [36], input_sha_func_0[36]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [37], input_sha_func_0[37]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [38], input_sha_func_0[38]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [39], input_sha_func_0[39]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [40], input_sha_func_0[40]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [41], input_sha_func_0[41]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [42], input_sha_func_0[42]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [43], input_sha_func_0[43]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [44], input_sha_func_0[44]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [45], input_sha_func_0[45]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [46], input_sha_func_0[46]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [47], input_sha_func_0[47]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [48], input_sha_func_0[48]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [49], input_sha_func_0[49]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [50], input_sha_func_0[50]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [51], input_sha_func_0[51]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [52], input_sha_func_0[52]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [53], input_sha_func_0[53]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [54], input_sha_func_0[54]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [55], input_sha_func_0[55]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [56], input_sha_func_0[56]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [57], input_sha_func_0[57]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [58], input_sha_func_0[58]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [59], input_sha_func_0[59]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [60], input_sha_func_0[60]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [61], input_sha_func_0[61]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [62], input_sha_func_0[62]);
  buf(\xm8051_golden_model_1.input_sha_func_0 [63], input_sha_func_0[63]);
  buf(\xm8051_golden_model_1.datain [0], proc_data_in[0]);
  buf(\xm8051_golden_model_1.datain [1], proc_data_in[1]);
  buf(\xm8051_golden_model_1.datain [2], proc_data_in[2]);
  buf(\xm8051_golden_model_1.datain [3], proc_data_in[3]);
  buf(\xm8051_golden_model_1.datain [4], proc_data_in[4]);
  buf(\xm8051_golden_model_1.datain [5], proc_data_in[5]);
  buf(\xm8051_golden_model_1.datain [6], proc_data_in[6]);
  buf(\xm8051_golden_model_1.datain [7], proc_data_in[7]);
  buf(\xm8051_golden_model_1.addrin [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.addrin [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.addrin [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.addrin [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.addrin [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.addrin [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.addrin [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.addrin [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.addrin [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.addrin [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.addrin [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.addrin [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.addrin [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.addrin [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.addrin [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.addrin [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.n0867 [0], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0867 [1], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0867 [2], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0867 [3], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0867 [4], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0867 [5], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0867 [6], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0867 [7], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0867 [8], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0867 [9], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0867 [10], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0867 [11], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0867 [12], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0867 [13], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0867 [14], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0867 [15], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0867 [16], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0867 [17], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0867 [18], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0867 [19], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0867 [20], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0867 [21], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0867 [22], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0867 [23], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0867 [24], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0867 [25], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0867 [26], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0867 [27], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0867 [28], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0867 [29], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0867 [30], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0867 [31], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0867 [32], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0867 [33], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0867 [34], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0867 [35], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0867 [36], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0867 [37], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0867 [38], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0867 [39], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0867 [40], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0867 [41], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0867 [42], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0867 [43], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0867 [44], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0867 [45], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0867 [46], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0867 [47], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0867 [48], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0867 [49], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0867 [50], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0867 [51], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0867 [52], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0867 [53], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0867 [54], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0867 [55], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0867 [56], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0867 [57], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0867 [58], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0867 [59], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0867 [60], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0867 [61], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0867 [62], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0867 [63], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.rst , rst);
  buf(\xm8051_golden_model_1.clk , clk);
  buf(\xm8051_golden_model_1.n0866 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0866 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0866 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0866 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0866 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0866 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0866 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0866 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0866 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0866 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0866 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0866 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0866 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0866 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0866 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0866 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0866 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0866 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0866 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0866 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0866 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0866 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0866 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0866 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0866 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0866 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0866 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0866 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0866 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0866 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0866 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0866 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0866 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0866 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0866 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0866 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0866 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0866 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0866 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0866 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0866 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0866 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0866 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0866 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0866 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0866 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0866 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0866 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0866 [48], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0866 [49], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0866 [50], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0866 [51], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0866 [52], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0866 [53], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0866 [54], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0866 [55], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0866 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0866 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0866 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0866 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0866 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0866 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0866 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0866 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0866 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0866 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0866 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0866 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0866 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0866 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0866 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0866 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0866 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0866 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0866 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0866 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0866 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0866 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0866 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0866 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0866 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0866 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0866 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0866 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0866 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0866 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0866 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0866 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0866 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0866 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0866 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0866 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0866 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0866 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0866 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0866 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0866 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0866 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0866 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0866 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0866 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0866 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0866 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0866 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0866 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0866 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0866 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0866 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0866 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0866 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0866 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0866 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0866 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0866 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0866 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0866 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0866 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0866 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0866 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0866 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0866 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0866 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0866 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0866 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0866 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0866 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0866 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0866 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0865 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0865 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0865 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0865 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0865 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0865 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0865 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0865 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0865 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0865 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0865 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0865 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0865 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0865 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0865 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0865 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0865 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0865 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0865 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0865 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0865 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0865 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0865 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0865 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0865 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0865 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0865 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0865 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0865 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0865 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0865 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0865 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0865 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0865 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0865 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0865 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0865 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0865 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0865 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0865 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0865 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0865 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0865 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0865 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0865 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0865 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0865 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0865 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0864 [0], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0864 [1], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0864 [2], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0864 [3], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0864 [4], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0864 [5], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0864 [6], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0864 [7], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0864 [8], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0864 [9], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0864 [10], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0864 [11], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0864 [12], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0864 [13], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0864 [14], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0864 [15], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0864 [16], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0864 [17], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0864 [18], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0864 [19], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0864 [20], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0864 [21], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0864 [22], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0864 [23], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0864 [24], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0864 [25], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0864 [26], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0864 [27], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0864 [28], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0864 [29], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0864 [30], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0864 [31], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0864 [32], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0864 [33], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0864 [34], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0864 [35], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0864 [36], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0864 [37], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0864 [38], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0864 [39], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0864 [40], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0864 [41], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0864 [42], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0864 [43], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0864 [44], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0864 [45], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0864 [46], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0864 [47], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0864 [48], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0864 [49], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0864 [50], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0864 [51], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0864 [52], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0864 [53], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0864 [54], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0864 [55], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0864 [56], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0864 [57], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0864 [58], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0864 [59], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0864 [60], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0864 [61], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0864 [62], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0864 [63], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0864 [64], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0864 [65], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0864 [66], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0864 [67], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0864 [68], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0864 [69], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0864 [70], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0864 [71], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0863 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0863 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0863 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0863 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0863 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0863 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0863 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0863 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0863 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0863 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0863 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0863 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0863 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0863 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0863 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0863 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0863 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0863 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0863 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0863 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0863 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0863 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0863 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0863 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0863 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0863 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0863 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0863 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0863 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0863 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0863 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0863 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0863 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0863 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0863 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0863 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0863 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0863 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0863 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0863 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0863 [40], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0863 [41], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0863 [42], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0863 [43], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0863 [44], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0863 [45], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0863 [46], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0863 [47], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0863 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0863 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0863 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0863 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0863 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0863 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0863 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0863 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0863 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0863 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0863 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0863 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0863 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0863 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0863 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0863 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0863 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0863 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0863 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0863 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0863 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0863 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0863 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0863 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0863 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0863 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0863 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0863 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0863 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0863 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0863 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0863 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0863 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0863 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0863 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0863 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0863 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0863 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0863 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0863 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0863 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0863 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0863 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0863 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0863 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0863 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0863 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0863 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0863 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0863 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0863 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0863 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0863 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0863 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0863 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0863 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0863 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0863 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0863 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0863 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0863 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0863 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0863 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0863 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0863 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0863 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0863 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0863 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0863 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0863 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0863 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0863 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0863 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0863 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0863 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0863 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0863 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0863 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0863 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0863 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0862 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0862 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0862 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0862 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0862 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0862 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0862 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0862 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0862 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0862 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0862 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0862 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0862 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0862 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0862 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0862 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0862 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0862 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0862 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0862 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0862 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0862 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0862 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0862 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0862 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0862 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0862 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0862 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0862 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0862 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0862 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0862 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0862 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0862 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0862 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0862 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0862 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0862 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0862 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0862 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0433 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0433 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0433 [2], \xm8051_golden_model_1.n0473 [2]);
  buf(\xm8051_golden_model_1.n0861 [0], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0861 [1], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0861 [2], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0861 [3], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0861 [4], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0861 [5], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0861 [6], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0861 [7], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0861 [8], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0861 [9], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0861 [10], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0861 [11], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0861 [12], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0861 [13], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0861 [14], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0861 [15], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0861 [16], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0861 [17], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0861 [18], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0861 [19], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0861 [20], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0861 [21], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0861 [22], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0861 [23], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0861 [24], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0861 [25], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0861 [26], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0861 [27], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0861 [28], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0861 [29], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0861 [30], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0861 [31], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0861 [32], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0861 [33], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0861 [34], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0861 [35], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0861 [36], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0861 [37], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0861 [38], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0861 [39], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0861 [40], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0861 [41], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0861 [42], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0861 [43], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0861 [44], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0861 [45], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0861 [46], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0861 [47], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0861 [48], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0861 [49], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0861 [50], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0861 [51], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0861 [52], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0861 [53], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0861 [54], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0861 [55], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0861 [56], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0861 [57], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0861 [58], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0861 [59], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0861 [60], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0861 [61], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0861 [62], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0861 [63], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0861 [64], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0861 [65], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0861 [66], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0861 [67], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0861 [68], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0861 [69], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0861 [70], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0861 [71], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0861 [72], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0861 [73], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0861 [74], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0861 [75], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0861 [76], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0861 [77], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0861 [78], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0861 [79], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0860 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0860 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0860 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0860 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0860 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0860 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0860 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0860 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0860 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0860 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0860 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0860 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0860 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0860 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0860 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0860 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0860 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0860 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0860 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0860 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0860 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0860 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0860 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0860 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0860 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0860 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0860 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0860 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0860 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0860 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0860 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0860 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0860 [32], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0860 [33], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0860 [34], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0860 [35], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0860 [36], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0860 [37], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0860 [38], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0860 [39], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0860 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0860 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0860 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0860 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0860 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0860 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0860 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0860 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0860 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0860 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0860 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0860 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0860 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0860 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0860 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0860 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0860 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0860 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0860 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0860 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0860 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0860 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0860 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0860 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0860 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0860 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0860 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0860 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0860 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0860 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0860 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0860 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0860 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0860 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0860 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0860 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0860 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0860 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0860 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0860 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0860 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0860 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0860 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0860 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0860 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0860 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0860 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0860 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0860 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0860 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0860 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0860 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0860 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0860 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0860 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0860 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0860 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0860 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0860 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0860 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0860 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0860 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0860 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0860 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0860 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0860 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0860 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0860 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0860 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0860 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0860 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0860 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0860 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0860 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0860 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0860 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0860 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0860 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0860 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0860 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0860 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0860 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0860 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0860 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0860 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0860 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0860 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0860 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0859 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0859 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0859 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0859 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0859 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0859 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0859 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0859 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0859 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0859 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0859 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0859 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0859 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0859 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0859 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0859 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0859 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0859 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0859 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0859 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0859 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0859 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0859 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0859 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0859 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0859 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0859 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0859 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0859 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0859 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0859 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0859 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0858 [0], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0858 [1], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0858 [2], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0858 [3], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0858 [4], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0858 [5], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0858 [6], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0858 [7], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0858 [8], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0858 [9], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0858 [10], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0858 [11], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0858 [12], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0858 [13], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0858 [14], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0858 [15], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0858 [16], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0858 [17], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0858 [18], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0858 [19], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0858 [20], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0858 [21], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0858 [22], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0858 [23], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0858 [24], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0858 [25], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0858 [26], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0858 [27], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0858 [28], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0858 [29], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0858 [30], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0858 [31], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0858 [32], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0858 [33], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0858 [34], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0858 [35], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0858 [36], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0858 [37], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0858 [38], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0858 [39], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0858 [40], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0858 [41], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0858 [42], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0858 [43], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0858 [44], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0858 [45], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0858 [46], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0858 [47], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0858 [48], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0858 [49], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0858 [50], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0858 [51], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0858 [52], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0858 [53], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0858 [54], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0858 [55], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0858 [56], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0858 [57], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0858 [58], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0858 [59], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0858 [60], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0858 [61], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0858 [62], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0858 [63], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0858 [64], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0858 [65], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0858 [66], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0858 [67], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0858 [68], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0858 [69], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0858 [70], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0858 [71], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0858 [72], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0858 [73], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0858 [74], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0858 [75], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0858 [76], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0858 [77], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0858 [78], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0858 [79], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0858 [80], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0858 [81], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0858 [82], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0858 [83], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0858 [84], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0858 [85], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0858 [86], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0858 [87], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0857 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0857 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0857 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0857 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0857 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0857 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0857 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0857 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0857 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0857 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0857 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0857 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0857 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0857 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0857 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0857 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0857 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0857 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0857 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0857 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0857 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0857 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0857 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0857 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0857 [24], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0857 [25], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0857 [26], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0857 [27], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0857 [28], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0857 [29], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0857 [30], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0857 [31], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0857 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0857 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0857 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0857 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0857 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0857 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0857 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0857 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0857 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0857 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0857 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0857 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0857 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0857 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0857 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0857 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0857 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0857 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0857 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0857 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0857 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0857 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0857 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0857 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0857 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0857 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0857 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0857 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0857 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0857 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0857 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0857 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0857 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0857 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0857 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0857 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0857 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0857 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0857 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0857 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0857 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0857 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0857 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0857 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0857 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0857 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0857 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0857 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0857 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0857 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0857 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0857 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0857 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0857 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0857 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0857 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0857 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0857 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0857 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0857 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0857 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0857 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0857 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0857 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0857 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0857 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0857 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0857 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0857 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0857 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0857 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0857 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0857 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0857 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0857 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0857 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0857 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0857 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0857 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0857 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0857 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0857 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0857 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0857 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0857 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0857 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0857 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0857 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0857 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0857 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0857 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0857 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0857 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0857 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0857 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0857 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0856 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0856 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0856 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0856 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0856 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0856 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0856 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0856 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0856 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0856 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0856 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0856 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0856 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0856 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0856 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0856 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0856 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0856 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0856 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0856 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0856 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0856 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0856 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0856 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0855 [0], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0855 [1], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0855 [2], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0855 [3], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0855 [4], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0855 [5], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0855 [6], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0855 [7], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0855 [8], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0855 [9], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0855 [10], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0855 [11], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0855 [12], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0855 [13], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0855 [14], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0855 [15], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0855 [16], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0855 [17], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0855 [18], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0855 [19], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0855 [20], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0855 [21], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0855 [22], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0855 [23], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0855 [24], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0855 [25], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0855 [26], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0855 [27], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0855 [28], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0855 [29], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0855 [30], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0855 [31], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0855 [32], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0855 [33], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0855 [34], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0855 [35], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0855 [36], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0855 [37], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0855 [38], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0855 [39], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0855 [40], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0855 [41], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0855 [42], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0855 [43], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0855 [44], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0855 [45], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0855 [46], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0855 [47], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0855 [48], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0855 [49], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0855 [50], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0855 [51], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0855 [52], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0855 [53], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0855 [54], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0855 [55], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0855 [56], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0855 [57], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0855 [58], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0855 [59], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0855 [60], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0855 [61], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0855 [62], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0855 [63], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0855 [64], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0855 [65], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0855 [66], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0855 [67], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0855 [68], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0855 [69], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0855 [70], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0855 [71], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0855 [72], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0855 [73], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0855 [74], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0855 [75], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0855 [76], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0855 [77], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0855 [78], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0855 [79], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0855 [80], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0855 [81], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0855 [82], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0855 [83], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0855 [84], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0855 [85], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0855 [86], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0855 [87], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0855 [88], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0855 [89], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0855 [90], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0855 [91], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0855 [92], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0855 [93], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0855 [94], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0855 [95], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0854 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0854 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0854 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0854 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0854 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0854 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0854 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0854 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0854 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0854 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0854 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0854 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0854 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0854 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0854 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0854 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0854 [16], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0854 [17], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0854 [18], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0854 [19], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0854 [20], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0854 [21], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0854 [22], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0854 [23], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0854 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0854 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0854 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0854 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0854 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0854 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0854 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0854 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0854 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0854 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0854 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0854 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0854 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0854 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0854 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0854 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0854 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0854 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0854 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0854 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0854 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0854 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0854 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0854 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0854 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0854 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0854 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0854 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0854 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0854 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0854 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0854 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0854 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0854 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0854 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0854 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0854 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0854 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0854 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0854 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0854 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0854 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0854 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0854 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0854 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0854 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0854 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0854 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0854 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0854 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0854 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0854 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0854 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0854 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0854 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0854 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0854 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0854 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0854 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0854 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0854 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0854 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0854 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0854 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0854 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0854 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0854 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0854 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0854 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0854 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0854 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0854 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0854 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0854 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0854 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0854 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0854 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0854 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0854 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0854 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0854 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0854 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0854 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0854 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0854 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0854 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0854 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0854 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0854 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0854 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0854 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0854 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0854 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0854 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0854 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0854 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0854 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0854 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0854 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0854 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0854 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0854 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0854 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0854 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0853 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0853 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0853 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0853 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0853 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0853 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0853 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0853 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0853 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0853 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0853 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0853 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0853 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0853 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0853 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0853 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0423 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0423 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0423 [2], \xm8051_golden_model_1.n0463 [2]);
  buf(\xm8051_golden_model_1.n0852 [0], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0852 [1], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0852 [2], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0852 [3], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0852 [4], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0852 [5], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0852 [6], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0852 [7], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0852 [8], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0852 [9], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0852 [10], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0852 [11], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0852 [12], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0852 [13], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0852 [14], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0852 [15], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0852 [16], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0852 [17], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0852 [18], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0852 [19], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0852 [20], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0852 [21], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0852 [22], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0852 [23], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0852 [24], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0852 [25], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0852 [26], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0852 [27], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0852 [28], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0852 [29], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0852 [30], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0852 [31], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0852 [32], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0852 [33], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0852 [34], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0852 [35], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0852 [36], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0852 [37], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0852 [38], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0852 [39], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0852 [40], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0852 [41], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0852 [42], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0852 [43], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0852 [44], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0852 [45], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0852 [46], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0852 [47], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0852 [48], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0852 [49], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0852 [50], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0852 [51], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0852 [52], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0852 [53], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0852 [54], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0852 [55], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0852 [56], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0852 [57], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0852 [58], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0852 [59], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0852 [60], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0852 [61], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0852 [62], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0852 [63], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0852 [64], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0852 [65], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0852 [66], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0852 [67], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0852 [68], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0852 [69], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0852 [70], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0852 [71], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0852 [72], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0852 [73], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0852 [74], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0852 [75], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0852 [76], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0852 [77], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0852 [78], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0852 [79], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0852 [80], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0852 [81], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0852 [82], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0852 [83], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0852 [84], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0852 [85], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0852 [86], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0852 [87], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0852 [88], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0852 [89], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0852 [90], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0852 [91], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0852 [92], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0852 [93], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0852 [94], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0852 [95], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0852 [96], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0852 [97], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0852 [98], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0852 [99], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0852 [100], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0852 [101], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0852 [102], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0852 [103], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0851 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0851 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0851 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0851 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0851 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0851 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0851 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0851 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0851 [8], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0851 [9], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0851 [10], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0851 [11], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0851 [12], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0851 [13], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0851 [14], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0851 [15], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0851 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0851 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0851 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0851 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0851 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0851 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0851 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0851 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0851 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0851 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0851 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0851 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0851 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0851 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0851 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0851 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0851 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0851 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0851 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0851 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0851 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0851 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0851 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0851 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0851 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0851 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0851 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0851 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0851 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0851 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0851 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0851 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0851 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0851 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0851 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0851 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0851 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0851 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0851 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0851 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0851 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0851 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0851 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0851 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0851 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0851 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0851 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0851 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0851 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0851 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0851 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0851 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0851 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0851 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0851 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0851 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0851 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0851 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0851 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0851 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0851 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0851 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0851 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0851 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0851 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0851 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0851 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0851 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0851 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0851 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0851 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0851 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0851 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0851 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0851 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0851 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0851 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0851 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0851 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0851 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0851 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0851 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0851 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0851 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0851 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0851 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0851 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0851 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0851 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0851 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0851 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0851 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0851 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0851 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0851 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0851 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0851 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0851 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0851 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0851 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0851 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0851 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0851 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0851 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0851 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0851 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0851 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0851 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0851 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0851 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0851 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0851 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0850 [0], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0850 [1], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0850 [2], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0850 [3], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0850 [4], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0850 [5], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0850 [6], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0850 [7], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0850 [8], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0850 [9], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0850 [10], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0850 [11], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0850 [12], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0850 [13], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0850 [14], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0850 [15], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0850 [16], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0850 [17], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0850 [18], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0850 [19], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0850 [20], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0850 [21], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0850 [22], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0850 [23], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0850 [24], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0850 [25], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0850 [26], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0850 [27], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0850 [28], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0850 [29], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0850 [30], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0850 [31], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0850 [32], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0850 [33], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0850 [34], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0850 [35], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0850 [36], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0850 [37], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0850 [38], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0850 [39], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0850 [40], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0850 [41], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0850 [42], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0850 [43], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0850 [44], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0850 [45], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0850 [46], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0850 [47], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0850 [48], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0850 [49], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0850 [50], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0850 [51], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0850 [52], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0850 [53], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0850 [54], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0850 [55], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0850 [56], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0850 [57], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0850 [58], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0850 [59], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0850 [60], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0850 [61], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0850 [62], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0850 [63], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0850 [64], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0850 [65], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0850 [66], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0850 [67], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0850 [68], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0850 [69], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0850 [70], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0850 [71], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0850 [72], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0850 [73], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0850 [74], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0850 [75], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0850 [76], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0850 [77], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0850 [78], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0850 [79], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0850 [80], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0850 [81], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0850 [82], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0850 [83], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0850 [84], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0850 [85], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0850 [86], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0850 [87], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0850 [88], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0850 [89], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0850 [90], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0850 [91], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0850 [92], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0850 [93], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0850 [94], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0850 [95], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0850 [96], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0850 [97], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0850 [98], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0850 [99], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0850 [100], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0850 [101], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0850 [102], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0850 [103], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0850 [104], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0850 [105], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0850 [106], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0850 [107], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0850 [108], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0850 [109], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0850 [110], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0850 [111], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0849 [0], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0849 [1], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0849 [2], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0849 [3], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0849 [4], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0849 [5], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0849 [6], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0849 [7], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0849 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0849 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0849 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0849 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0849 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0849 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0849 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0849 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0849 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0849 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0849 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0849 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0849 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0849 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0849 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0849 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0849 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0849 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0849 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0849 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0849 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0849 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0849 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0849 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0849 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0849 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0849 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0849 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0849 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0849 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0849 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0849 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0849 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0849 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0849 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0849 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0849 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0849 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0849 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0849 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0849 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0849 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0849 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0849 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0849 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0849 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0849 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0849 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0849 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0849 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0849 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0849 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0849 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0849 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0849 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0849 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0849 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0849 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0849 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0849 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0849 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0849 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0849 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0849 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0849 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0849 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0849 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0849 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0849 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0849 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0849 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0849 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0849 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0849 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0849 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0849 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0849 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0849 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0849 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0849 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0849 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0849 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0849 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0849 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0849 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0849 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0849 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0849 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0849 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0849 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0849 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0849 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0849 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0849 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0849 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0849 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0849 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0849 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0849 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0849 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0849 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0849 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0849 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0849 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0849 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0849 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0849 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0849 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0849 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0849 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0849 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0849 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0849 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0849 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0849 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0849 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0849 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0849 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0849 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0849 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n1285 [0], input_sha_func_44[0]);
  buf(\xm8051_golden_model_1.n1285 [1], input_sha_func_44[1]);
  buf(\xm8051_golden_model_1.n1285 [2], input_sha_func_44[2]);
  buf(\xm8051_golden_model_1.n1285 [3], input_sha_func_44[3]);
  buf(\xm8051_golden_model_1.n1285 [4], input_sha_func_44[4]);
  buf(\xm8051_golden_model_1.n1285 [5], input_sha_func_44[5]);
  buf(\xm8051_golden_model_1.n1285 [6], input_sha_func_44[6]);
  buf(\xm8051_golden_model_1.n1285 [7], input_sha_func_44[7]);
  buf(\xm8051_golden_model_1.n1285 [8], input_sha_func_44[8]);
  buf(\xm8051_golden_model_1.n1285 [9], input_sha_func_44[9]);
  buf(\xm8051_golden_model_1.n1285 [10], input_sha_func_44[10]);
  buf(\xm8051_golden_model_1.n1285 [11], input_sha_func_44[11]);
  buf(\xm8051_golden_model_1.n1285 [12], input_sha_func_44[12]);
  buf(\xm8051_golden_model_1.n1285 [13], input_sha_func_44[13]);
  buf(\xm8051_golden_model_1.n1285 [14], input_sha_func_44[14]);
  buf(\xm8051_golden_model_1.n1285 [15], input_sha_func_44[15]);
  buf(\xm8051_golden_model_1.n1285 [16], input_sha_func_44[16]);
  buf(\xm8051_golden_model_1.n1285 [17], input_sha_func_44[17]);
  buf(\xm8051_golden_model_1.n1285 [18], input_sha_func_44[18]);
  buf(\xm8051_golden_model_1.n1285 [19], input_sha_func_44[19]);
  buf(\xm8051_golden_model_1.n1285 [20], input_sha_func_44[20]);
  buf(\xm8051_golden_model_1.n1285 [21], input_sha_func_44[21]);
  buf(\xm8051_golden_model_1.n1285 [22], input_sha_func_44[22]);
  buf(\xm8051_golden_model_1.n1285 [23], input_sha_func_44[23]);
  buf(\xm8051_golden_model_1.n1285 [24], input_sha_func_44[24]);
  buf(\xm8051_golden_model_1.n1285 [25], input_sha_func_44[25]);
  buf(\xm8051_golden_model_1.n1285 [26], input_sha_func_44[26]);
  buf(\xm8051_golden_model_1.n1285 [27], input_sha_func_44[27]);
  buf(\xm8051_golden_model_1.n1285 [28], input_sha_func_44[28]);
  buf(\xm8051_golden_model_1.n1285 [29], input_sha_func_44[29]);
  buf(\xm8051_golden_model_1.n1285 [30], input_sha_func_44[30]);
  buf(\xm8051_golden_model_1.n1285 [31], input_sha_func_44[31]);
  buf(\xm8051_golden_model_1.n1285 [32], input_sha_func_43[0]);
  buf(\xm8051_golden_model_1.n1285 [33], input_sha_func_43[1]);
  buf(\xm8051_golden_model_1.n1285 [34], input_sha_func_43[2]);
  buf(\xm8051_golden_model_1.n1285 [35], input_sha_func_43[3]);
  buf(\xm8051_golden_model_1.n1285 [36], input_sha_func_43[4]);
  buf(\xm8051_golden_model_1.n1285 [37], input_sha_func_43[5]);
  buf(\xm8051_golden_model_1.n1285 [38], input_sha_func_43[6]);
  buf(\xm8051_golden_model_1.n1285 [39], input_sha_func_43[7]);
  buf(\xm8051_golden_model_1.n1285 [40], input_sha_func_43[8]);
  buf(\xm8051_golden_model_1.n1285 [41], input_sha_func_43[9]);
  buf(\xm8051_golden_model_1.n1285 [42], input_sha_func_43[10]);
  buf(\xm8051_golden_model_1.n1285 [43], input_sha_func_43[11]);
  buf(\xm8051_golden_model_1.n1285 [44], input_sha_func_43[12]);
  buf(\xm8051_golden_model_1.n1285 [45], input_sha_func_43[13]);
  buf(\xm8051_golden_model_1.n1285 [46], input_sha_func_43[14]);
  buf(\xm8051_golden_model_1.n1285 [47], input_sha_func_43[15]);
  buf(\xm8051_golden_model_1.n1285 [48], input_sha_func_43[16]);
  buf(\xm8051_golden_model_1.n1285 [49], input_sha_func_43[17]);
  buf(\xm8051_golden_model_1.n1285 [50], input_sha_func_43[18]);
  buf(\xm8051_golden_model_1.n1285 [51], input_sha_func_43[19]);
  buf(\xm8051_golden_model_1.n1285 [52], input_sha_func_43[20]);
  buf(\xm8051_golden_model_1.n1285 [53], input_sha_func_43[21]);
  buf(\xm8051_golden_model_1.n1285 [54], input_sha_func_43[22]);
  buf(\xm8051_golden_model_1.n1285 [55], input_sha_func_43[23]);
  buf(\xm8051_golden_model_1.n1285 [56], input_sha_func_43[24]);
  buf(\xm8051_golden_model_1.n1285 [57], input_sha_func_43[25]);
  buf(\xm8051_golden_model_1.n1285 [58], input_sha_func_43[26]);
  buf(\xm8051_golden_model_1.n1285 [59], input_sha_func_43[27]);
  buf(\xm8051_golden_model_1.n1285 [60], input_sha_func_43[28]);
  buf(\xm8051_golden_model_1.n1285 [61], input_sha_func_43[29]);
  buf(\xm8051_golden_model_1.n1285 [62], input_sha_func_43[30]);
  buf(\xm8051_golden_model_1.n1285 [63], input_sha_func_43[31]);
  buf(\xm8051_golden_model_1.n1285 [64], input_sha_func_43[32]);
  buf(\xm8051_golden_model_1.n1285 [65], input_sha_func_43[33]);
  buf(\xm8051_golden_model_1.n1285 [66], input_sha_func_43[34]);
  buf(\xm8051_golden_model_1.n1285 [67], input_sha_func_43[35]);
  buf(\xm8051_golden_model_1.n1285 [68], input_sha_func_43[36]);
  buf(\xm8051_golden_model_1.n1285 [69], input_sha_func_43[37]);
  buf(\xm8051_golden_model_1.n1285 [70], input_sha_func_43[38]);
  buf(\xm8051_golden_model_1.n1285 [71], input_sha_func_43[39]);
  buf(\xm8051_golden_model_1.n1285 [72], input_sha_func_43[40]);
  buf(\xm8051_golden_model_1.n1285 [73], input_sha_func_43[41]);
  buf(\xm8051_golden_model_1.n1285 [74], input_sha_func_43[42]);
  buf(\xm8051_golden_model_1.n1285 [75], input_sha_func_43[43]);
  buf(\xm8051_golden_model_1.n1285 [76], input_sha_func_43[44]);
  buf(\xm8051_golden_model_1.n1285 [77], input_sha_func_43[45]);
  buf(\xm8051_golden_model_1.n1285 [78], input_sha_func_43[46]);
  buf(\xm8051_golden_model_1.n1285 [79], input_sha_func_43[47]);
  buf(\xm8051_golden_model_1.n1285 [80], input_sha_func_43[48]);
  buf(\xm8051_golden_model_1.n1285 [81], input_sha_func_43[49]);
  buf(\xm8051_golden_model_1.n1285 [82], input_sha_func_43[50]);
  buf(\xm8051_golden_model_1.n1285 [83], input_sha_func_43[51]);
  buf(\xm8051_golden_model_1.n1285 [84], input_sha_func_43[52]);
  buf(\xm8051_golden_model_1.n1285 [85], input_sha_func_43[53]);
  buf(\xm8051_golden_model_1.n1285 [86], input_sha_func_43[54]);
  buf(\xm8051_golden_model_1.n1285 [87], input_sha_func_43[55]);
  buf(\xm8051_golden_model_1.n1285 [88], input_sha_func_43[56]);
  buf(\xm8051_golden_model_1.n1285 [89], input_sha_func_43[57]);
  buf(\xm8051_golden_model_1.n1285 [90], input_sha_func_43[58]);
  buf(\xm8051_golden_model_1.n1285 [91], input_sha_func_43[59]);
  buf(\xm8051_golden_model_1.n1285 [92], input_sha_func_43[60]);
  buf(\xm8051_golden_model_1.n1285 [93], input_sha_func_43[61]);
  buf(\xm8051_golden_model_1.n1285 [94], input_sha_func_43[62]);
  buf(\xm8051_golden_model_1.n1285 [95], input_sha_func_43[63]);
  buf(\xm8051_golden_model_1.n1285 [96], input_sha_func_42[0]);
  buf(\xm8051_golden_model_1.n1285 [97], input_sha_func_42[1]);
  buf(\xm8051_golden_model_1.n1285 [98], input_sha_func_42[2]);
  buf(\xm8051_golden_model_1.n1285 [99], input_sha_func_42[3]);
  buf(\xm8051_golden_model_1.n1285 [100], input_sha_func_42[4]);
  buf(\xm8051_golden_model_1.n1285 [101], input_sha_func_42[5]);
  buf(\xm8051_golden_model_1.n1285 [102], input_sha_func_42[6]);
  buf(\xm8051_golden_model_1.n1285 [103], input_sha_func_42[7]);
  buf(\xm8051_golden_model_1.n1285 [104], input_sha_func_42[8]);
  buf(\xm8051_golden_model_1.n1285 [105], input_sha_func_42[9]);
  buf(\xm8051_golden_model_1.n1285 [106], input_sha_func_42[10]);
  buf(\xm8051_golden_model_1.n1285 [107], input_sha_func_42[11]);
  buf(\xm8051_golden_model_1.n1285 [108], input_sha_func_42[12]);
  buf(\xm8051_golden_model_1.n1285 [109], input_sha_func_42[13]);
  buf(\xm8051_golden_model_1.n1285 [110], input_sha_func_42[14]);
  buf(\xm8051_golden_model_1.n1285 [111], input_sha_func_42[15]);
  buf(\xm8051_golden_model_1.n1285 [112], input_sha_func_42[16]);
  buf(\xm8051_golden_model_1.n1285 [113], input_sha_func_42[17]);
  buf(\xm8051_golden_model_1.n1285 [114], input_sha_func_42[18]);
  buf(\xm8051_golden_model_1.n1285 [115], input_sha_func_42[19]);
  buf(\xm8051_golden_model_1.n1285 [116], input_sha_func_42[20]);
  buf(\xm8051_golden_model_1.n1285 [117], input_sha_func_42[21]);
  buf(\xm8051_golden_model_1.n1285 [118], input_sha_func_42[22]);
  buf(\xm8051_golden_model_1.n1285 [119], input_sha_func_42[23]);
  buf(\xm8051_golden_model_1.n1285 [120], input_sha_func_42[24]);
  buf(\xm8051_golden_model_1.n1285 [121], input_sha_func_42[25]);
  buf(\xm8051_golden_model_1.n1285 [122], input_sha_func_42[26]);
  buf(\xm8051_golden_model_1.n1285 [123], input_sha_func_42[27]);
  buf(\xm8051_golden_model_1.n1285 [124], input_sha_func_42[28]);
  buf(\xm8051_golden_model_1.n1285 [125], input_sha_func_42[29]);
  buf(\xm8051_golden_model_1.n1285 [126], input_sha_func_42[30]);
  buf(\xm8051_golden_model_1.n1285 [127], input_sha_func_42[31]);
  buf(\xm8051_golden_model_1.n1285 [128], input_sha_func_42[32]);
  buf(\xm8051_golden_model_1.n1285 [129], input_sha_func_42[33]);
  buf(\xm8051_golden_model_1.n1285 [130], input_sha_func_42[34]);
  buf(\xm8051_golden_model_1.n1285 [131], input_sha_func_42[35]);
  buf(\xm8051_golden_model_1.n1285 [132], input_sha_func_42[36]);
  buf(\xm8051_golden_model_1.n1285 [133], input_sha_func_42[37]);
  buf(\xm8051_golden_model_1.n1285 [134], input_sha_func_42[38]);
  buf(\xm8051_golden_model_1.n1285 [135], input_sha_func_42[39]);
  buf(\xm8051_golden_model_1.n1285 [136], input_sha_func_42[40]);
  buf(\xm8051_golden_model_1.n1285 [137], input_sha_func_42[41]);
  buf(\xm8051_golden_model_1.n1285 [138], input_sha_func_42[42]);
  buf(\xm8051_golden_model_1.n1285 [139], input_sha_func_42[43]);
  buf(\xm8051_golden_model_1.n1285 [140], input_sha_func_42[44]);
  buf(\xm8051_golden_model_1.n1285 [141], input_sha_func_42[45]);
  buf(\xm8051_golden_model_1.n1285 [142], input_sha_func_42[46]);
  buf(\xm8051_golden_model_1.n1285 [143], input_sha_func_42[47]);
  buf(\xm8051_golden_model_1.n1285 [144], input_sha_func_42[48]);
  buf(\xm8051_golden_model_1.n1285 [145], input_sha_func_42[49]);
  buf(\xm8051_golden_model_1.n1285 [146], input_sha_func_42[50]);
  buf(\xm8051_golden_model_1.n1285 [147], input_sha_func_42[51]);
  buf(\xm8051_golden_model_1.n1285 [148], input_sha_func_42[52]);
  buf(\xm8051_golden_model_1.n1285 [149], input_sha_func_42[53]);
  buf(\xm8051_golden_model_1.n1285 [150], input_sha_func_42[54]);
  buf(\xm8051_golden_model_1.n1285 [151], input_sha_func_42[55]);
  buf(\xm8051_golden_model_1.n1285 [152], input_sha_func_42[56]);
  buf(\xm8051_golden_model_1.n1285 [153], input_sha_func_42[57]);
  buf(\xm8051_golden_model_1.n1285 [154], input_sha_func_42[58]);
  buf(\xm8051_golden_model_1.n1285 [155], input_sha_func_42[59]);
  buf(\xm8051_golden_model_1.n1285 [156], input_sha_func_42[60]);
  buf(\xm8051_golden_model_1.n1285 [157], input_sha_func_42[61]);
  buf(\xm8051_golden_model_1.n1285 [158], input_sha_func_42[62]);
  buf(\xm8051_golden_model_1.n1285 [159], input_sha_func_42[63]);
  buf(\xm8051_golden_model_1.n0413 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0413 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0413 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n0413 [3], \xm8051_golden_model_1.sha_bytes_processed [3]);
  buf(\xm8051_golden_model_1.n0401 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0401 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0401 [2], \xm8051_golden_model_1.n0483 [2]);
  buf(\xm8051_golden_model_1.n0401 [3], \xm8051_golden_model_1.n0483 [3]);
  buf(\xm8051_golden_model_1.n0830 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0830 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0830 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0830 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0830 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0830 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0830 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0830 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0830 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0830 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0830 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0830 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0830 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0830 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0830 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0830 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0830 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0830 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0830 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0830 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0830 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0830 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0830 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0830 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0830 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0830 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0830 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0830 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0830 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0830 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0830 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0830 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0830 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0830 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0830 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0830 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0830 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0830 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0830 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0830 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0830 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0830 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0830 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0830 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0830 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0830 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0830 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0830 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0830 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0830 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0830 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0830 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0830 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0830 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0830 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0830 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0830 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0830 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0830 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0830 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0830 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0830 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0830 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0830 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0830 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0830 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0830 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0830 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0830 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0830 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0830 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0830 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0830 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0830 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0830 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0830 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0830 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0830 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0830 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0830 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0830 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0830 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0830 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0830 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0830 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0830 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0830 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0830 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0830 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0830 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0830 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0830 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0830 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0830 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0830 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0830 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0830 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0830 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0830 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0830 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0830 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0830 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0830 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0830 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0830 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0830 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0830 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0830 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0830 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0830 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0830 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0830 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0830 [120], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0830 [121], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0830 [122], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0830 [123], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0830 [124], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0830 [125], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0830 [126], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0830 [127], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0829 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0829 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0829 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0829 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0829 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0829 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0829 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0829 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0829 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0829 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0829 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0829 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0829 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0829 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0829 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0829 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0829 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0829 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0829 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0829 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0829 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0829 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0829 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0829 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0829 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0829 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0829 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0829 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0829 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0829 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0829 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0829 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0829 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0829 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0829 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0829 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0829 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0829 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0829 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0829 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0829 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0829 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0829 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0829 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0829 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0829 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0829 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0829 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0829 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0829 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0829 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0829 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0829 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0829 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0829 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0829 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0829 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0829 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0829 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0829 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0829 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0829 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0829 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0829 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0829 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0829 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0829 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0829 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0829 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0829 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0829 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0829 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0829 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0829 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0829 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0829 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0829 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0829 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0829 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0829 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0829 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0829 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0829 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0829 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0829 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0829 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0829 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0829 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0829 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0829 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0829 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0829 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0829 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0829 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0829 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0829 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0829 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0829 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0829 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0829 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0829 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0829 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0829 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0829 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0829 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0829 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0829 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0829 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0829 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0829 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0829 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0829 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0829 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0829 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0829 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0829 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0829 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0829 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0829 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0829 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0828 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0828 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0828 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0828 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0828 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0828 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0828 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0828 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0828 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0828 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0828 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0828 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0828 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0828 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0828 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0828 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0828 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0828 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0828 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0828 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0828 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0828 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0828 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0828 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0828 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0828 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0828 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0828 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0828 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0828 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0828 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0828 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0828 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0828 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0828 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0828 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0828 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0828 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0828 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0828 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0828 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0828 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0828 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0828 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0828 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0828 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0828 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0828 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0828 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0828 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0828 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0828 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0828 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0828 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0828 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0828 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0828 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0828 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0828 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0828 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0828 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0828 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0828 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0828 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0828 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0828 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0828 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0828 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0828 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0828 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0828 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0828 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0828 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0828 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0828 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0828 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0828 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0828 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0828 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0828 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0828 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0828 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0828 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0828 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0828 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0828 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0828 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0828 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0828 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0828 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0828 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0828 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0828 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0828 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0828 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0828 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0828 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0828 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0828 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0828 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0828 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0828 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0828 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0828 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0828 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0828 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0828 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0828 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0828 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0828 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0828 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0828 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0828 [112], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0828 [113], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0828 [114], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0828 [115], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0828 [116], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0828 [117], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0828 [118], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0828 [119], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0827 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0827 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0827 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0827 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0827 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0827 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0827 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0827 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0827 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0827 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0827 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0827 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0827 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0827 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0827 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0827 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0827 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0827 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0827 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0827 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0827 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0827 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0827 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0827 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0827 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0827 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0827 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0827 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0827 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0827 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0827 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0827 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0827 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0827 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0827 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0827 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0827 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0827 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0827 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0827 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0827 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0827 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0827 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0827 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0827 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0827 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0827 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0827 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0827 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0827 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0827 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0827 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0827 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0827 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0827 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0827 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0827 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0827 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0827 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0827 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0827 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0827 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0827 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0827 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0827 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0827 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0827 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0827 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0827 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0827 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0827 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0827 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0827 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0827 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0827 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0827 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0827 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0827 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0827 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0827 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0827 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0827 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0827 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0827 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0827 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0827 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0827 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0827 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0827 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0827 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0827 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0827 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0827 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0827 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0827 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0827 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0827 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0827 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0827 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0827 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0827 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0827 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0827 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0827 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0827 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0827 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0827 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0827 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0827 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0827 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0827 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0827 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0826 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0826 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0826 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0826 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0826 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0826 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0826 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0826 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0826 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0826 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0826 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0826 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0826 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0826 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0826 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0826 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0826 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0826 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0826 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0826 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0826 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0826 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0826 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0826 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0826 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0826 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0826 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0826 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0826 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0826 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0826 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0826 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0826 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0826 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0826 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0826 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0826 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0826 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0826 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0826 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0826 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0826 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0826 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0826 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0826 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0826 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0826 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0826 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0826 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0826 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0826 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0826 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0826 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0826 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0826 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0826 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0826 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0826 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0826 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0826 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0826 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0826 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0826 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0826 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0826 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0826 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0826 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0826 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0826 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0826 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0826 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0826 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0826 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0826 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0826 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0826 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0826 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0826 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0826 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0826 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0826 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0826 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0826 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0826 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0826 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0826 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0826 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0826 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0826 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0826 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0826 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0826 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0826 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0826 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0826 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0826 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0826 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0826 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0826 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0826 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0826 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0826 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0826 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0826 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0826 [104], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0826 [105], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0826 [106], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0826 [107], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0826 [108], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0826 [109], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0826 [110], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0826 [111], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0826 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0826 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0826 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0826 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0826 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0826 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0826 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0826 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0826 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0826 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0826 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0826 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0826 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0826 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0826 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0826 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0825 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0825 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0825 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0825 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0825 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0825 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0825 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0825 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0825 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0825 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0825 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0825 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0825 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0825 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0825 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0825 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0825 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0825 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0825 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0825 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0825 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0825 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0825 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0825 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0825 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0825 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0825 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0825 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0825 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0825 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0825 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0825 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0825 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0825 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0825 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0825 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0825 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0825 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0825 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0825 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0825 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0825 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0825 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0825 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0825 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0825 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0825 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0825 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0825 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0825 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0825 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0825 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0825 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0825 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0825 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0825 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0825 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0825 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0825 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0825 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0825 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0825 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0825 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0825 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0825 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0825 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0825 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0825 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0825 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0825 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0825 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0825 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0825 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0825 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0825 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0825 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0825 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0825 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0825 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0825 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0825 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0825 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0825 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0825 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0825 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0825 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0825 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0825 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0825 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0825 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0825 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0825 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0825 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0825 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0825 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0825 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0825 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0825 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0825 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0825 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0825 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0825 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0825 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0825 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0389 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0389 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0389 [2], \xm8051_golden_model_1.n0473 [2]);
  buf(\xm8051_golden_model_1.n0389 [3], \xm8051_golden_model_1.n0473 [3]);
  buf(\xm8051_golden_model_1.n0824 [0], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0824 [1], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0824 [2], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0824 [3], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0824 [4], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0824 [5], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0824 [6], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0824 [7], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0824 [8], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0824 [9], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0824 [10], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0824 [11], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0824 [12], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0824 [13], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0824 [14], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0824 [15], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0823 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0823 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0823 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0823 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0823 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0823 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0823 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0823 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0823 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0823 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0823 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0823 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0823 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0823 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0823 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0823 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0823 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0823 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0823 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0823 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0823 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0823 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0823 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0823 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0823 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0823 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0823 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0823 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0823 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0823 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0823 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0823 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0823 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0823 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0823 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0823 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0823 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0823 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0823 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0823 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0823 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0823 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0823 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0823 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0823 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0823 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0823 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0823 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0823 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0823 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0823 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0823 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0823 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0823 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0823 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0823 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0823 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0823 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0823 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0823 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0823 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0823 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0823 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0823 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0823 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0823 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0823 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0823 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0823 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0823 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0823 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0823 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0823 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0823 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0823 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0823 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0823 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0823 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0823 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0823 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0823 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0823 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0823 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0823 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0823 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0823 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0823 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0823 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0823 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0823 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0823 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0823 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0823 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0823 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0823 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0823 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0823 [96], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0823 [97], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0823 [98], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0823 [99], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0823 [100], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0823 [101], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0823 [102], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0823 [103], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0823 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0823 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0823 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0823 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0823 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0823 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0823 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0823 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0823 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0823 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0823 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0823 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0823 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0823 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0823 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0823 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0823 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0823 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0823 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0823 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0823 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0823 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0823 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0823 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0822 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0822 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0822 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0822 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0822 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0822 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0822 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0822 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0822 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0822 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0822 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0822 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0822 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0822 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0822 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0822 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0822 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0822 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0822 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0822 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0822 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0822 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0822 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0822 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0822 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0822 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0822 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0822 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0822 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0822 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0822 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0822 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0822 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0822 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0822 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0822 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0822 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0822 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0822 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0822 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0822 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0822 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0822 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0822 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0822 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0822 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0822 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0822 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0822 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0822 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0822 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0822 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0822 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0822 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0822 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0822 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0822 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0822 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0822 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0822 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0822 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0822 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0822 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0822 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0822 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0822 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0822 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0822 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0822 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0822 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0822 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0822 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0822 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0822 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0822 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0822 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0822 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0822 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0822 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0822 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0822 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0822 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0822 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0822 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0822 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0822 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0822 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0822 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0822 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0822 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0822 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0822 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0822 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0822 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0822 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0822 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0821 [0], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0821 [1], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0821 [2], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0821 [3], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0821 [4], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0821 [5], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0821 [6], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0821 [7], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0821 [8], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0821 [9], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0821 [10], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0821 [11], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0821 [12], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0821 [13], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0821 [14], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0821 [15], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0821 [16], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0821 [17], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0821 [18], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0821 [19], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0821 [20], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0821 [21], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0821 [22], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0821 [23], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0820 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0820 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0820 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0820 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0820 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0820 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0820 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0820 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0820 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0820 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0820 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0820 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0820 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0820 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0820 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0820 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0820 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0820 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0820 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0820 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0820 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0820 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0820 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0820 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0820 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0820 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0820 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0820 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0820 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0820 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0820 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0820 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0820 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0820 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0820 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0820 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0820 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0820 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0820 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0820 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0820 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0820 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0820 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0820 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0820 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0820 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0820 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0820 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0820 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0820 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0820 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0820 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0820 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0820 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0820 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0820 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0820 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0820 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0820 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0820 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0820 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0820 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0820 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0820 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0820 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0820 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0820 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0820 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0820 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0820 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0820 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0820 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0820 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0820 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0820 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0820 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0820 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0820 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0820 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0820 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0820 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0820 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0820 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0820 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0820 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0820 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0820 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0820 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0820 [88], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0820 [89], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0820 [90], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0820 [91], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0820 [92], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0820 [93], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0820 [94], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0820 [95], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0820 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0820 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0820 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0820 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0820 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0820 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0820 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0820 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0820 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0820 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0820 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0820 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0820 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0820 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0820 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0820 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0820 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0820 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0820 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0820 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0820 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0820 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0820 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0820 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0820 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0820 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0820 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0820 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0820 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0820 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0820 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0820 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0819 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0819 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0819 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0819 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0819 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0819 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0819 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0819 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0819 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0819 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0819 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0819 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0819 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0819 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0819 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0819 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0819 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0819 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0819 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0819 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0819 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0819 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0819 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0819 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0819 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0819 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0819 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0819 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0819 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0819 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0819 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0819 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0819 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0819 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0819 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0819 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0819 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0819 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0819 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0819 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0819 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0819 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0819 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0819 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0819 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0819 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0819 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0819 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0819 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0819 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0819 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0819 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0819 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0819 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0819 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0819 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0819 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0819 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0819 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0819 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0819 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0819 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0819 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0819 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0819 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0819 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0819 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0819 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0819 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0819 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0819 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0819 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0819 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0819 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0819 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0819 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0819 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0819 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0819 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0819 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0819 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0819 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0819 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0819 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0819 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0819 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0819 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0819 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0818 [0], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0818 [1], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0818 [2], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0818 [3], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0818 [4], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0818 [5], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0818 [6], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0818 [7], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0818 [8], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0818 [9], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0818 [10], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0818 [11], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0818 [12], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0818 [13], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0818 [14], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0818 [15], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0818 [16], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0818 [17], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0818 [18], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0818 [19], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0818 [20], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0818 [21], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0818 [22], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0818 [23], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0818 [24], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0818 [25], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0818 [26], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0818 [27], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0818 [28], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0818 [29], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0818 [30], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0818 [31], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0817 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0817 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0817 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0817 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0817 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0817 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0817 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0817 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0817 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0817 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0817 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0817 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0817 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0817 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0817 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0817 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0817 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0817 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0817 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0817 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0817 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0817 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0817 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0817 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0817 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0817 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0817 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0817 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0817 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0817 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0817 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0817 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0817 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0817 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0817 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0817 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0817 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0817 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0817 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0817 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0817 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0817 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0817 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0817 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0817 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0817 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0817 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0817 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0817 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0817 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0817 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0817 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0817 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0817 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0817 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0817 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0817 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0817 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0817 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0817 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0817 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0817 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0817 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0817 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0817 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0817 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0817 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0817 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0817 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0817 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0817 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0817 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0817 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0817 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0817 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0817 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0817 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0817 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0817 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0817 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0817 [80], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0817 [81], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0817 [82], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0817 [83], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0817 [84], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0817 [85], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0817 [86], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0817 [87], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0817 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0817 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0817 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0817 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0817 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0817 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0817 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0817 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0817 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0817 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0817 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0817 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0817 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0817 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0817 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0817 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0817 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0817 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0817 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0817 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0817 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0817 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0817 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0817 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0817 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0817 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0817 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0817 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0817 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0817 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0817 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0817 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0817 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0817 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0817 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0817 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0817 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0817 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0817 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0817 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0816 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0816 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0816 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0816 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0816 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0816 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0816 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0816 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0816 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0816 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0816 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0816 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0816 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0816 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0816 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0816 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0816 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0816 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0816 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0816 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0816 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0816 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0816 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0816 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0816 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0816 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0816 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0816 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0816 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0816 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0816 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0816 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0816 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0816 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0816 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0816 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0816 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0816 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0816 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0816 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0816 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0816 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0816 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0816 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0816 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0816 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0816 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0816 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0816 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0816 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0816 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0816 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0816 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0816 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0816 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0816 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0816 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0816 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0816 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0816 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0816 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0816 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0816 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0816 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0816 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0816 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0816 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0816 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0816 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0816 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0816 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0816 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0816 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0816 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0816 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0816 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0816 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0816 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0816 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0816 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0815 [0], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0815 [1], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0815 [2], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0815 [3], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0815 [4], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0815 [5], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0815 [6], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0815 [7], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0815 [8], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0815 [9], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0815 [10], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0815 [11], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0815 [12], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0815 [13], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0815 [14], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0815 [15], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0815 [16], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0815 [17], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0815 [18], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0815 [19], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0815 [20], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0815 [21], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0815 [22], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0815 [23], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0815 [24], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0815 [25], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0815 [26], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0815 [27], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0815 [28], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0815 [29], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0815 [30], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0815 [31], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0815 [32], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0815 [33], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0815 [34], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0815 [35], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0815 [36], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0815 [37], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0815 [38], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0815 [39], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0377 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0377 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0377 [2], \xm8051_golden_model_1.n0463 [2]);
  buf(\xm8051_golden_model_1.n0377 [3], \xm8051_golden_model_1.n0463 [3]);
  buf(\xm8051_golden_model_1.n0814 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0814 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0814 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0814 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0814 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0814 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0814 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0814 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0814 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0814 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0814 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0814 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0814 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0814 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0814 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0814 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0814 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0814 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0814 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0814 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0814 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0814 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0814 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0814 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0814 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0814 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0814 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0814 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0814 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0814 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0814 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0814 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0814 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0814 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0814 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0814 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0814 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0814 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0814 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0814 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0814 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0814 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0814 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0814 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0814 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0814 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0814 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0814 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0814 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0814 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0814 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0814 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0814 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0814 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0814 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0814 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0814 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0814 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0814 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0814 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0814 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0814 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0814 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0814 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0814 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0814 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0814 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0814 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0814 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0814 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0814 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0814 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0814 [72], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0814 [73], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0814 [74], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0814 [75], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0814 [76], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0814 [77], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0814 [78], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0814 [79], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0814 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0814 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0814 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0814 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0814 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0814 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0814 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0814 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0814 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0814 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0814 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0814 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0814 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0814 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0814 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0814 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0814 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0814 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0814 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0814 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0814 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0814 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0814 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0814 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0814 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0814 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0814 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0814 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0814 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0814 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0814 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0814 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0814 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0814 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0814 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0814 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0814 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0814 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0814 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0814 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0814 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0814 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0814 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0814 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0814 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0814 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0814 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0814 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0813 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0813 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0813 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0813 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0813 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0813 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0813 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0813 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0813 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0813 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0813 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0813 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0813 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0813 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0813 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0813 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0813 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0813 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0813 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0813 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0813 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0813 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0813 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0813 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0813 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0813 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0813 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0813 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0813 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0813 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0813 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0813 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0813 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0813 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0813 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0813 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0813 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0813 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0813 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0813 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0813 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0813 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0813 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0813 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0813 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0813 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0813 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0813 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0813 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0813 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0813 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0813 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0813 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0813 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0813 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0813 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0813 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0813 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0813 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0813 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0813 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0813 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0813 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0813 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0813 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0813 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0813 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0813 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0813 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0813 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0813 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0813 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0812 [0], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0812 [1], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0812 [2], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0812 [3], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0812 [4], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0812 [5], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0812 [6], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0812 [7], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0812 [8], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0812 [9], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0812 [10], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0812 [11], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0812 [12], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0812 [13], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0812 [14], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0812 [15], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0812 [16], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0812 [17], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0812 [18], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0812 [19], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0812 [20], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0812 [21], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0812 [22], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0812 [23], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0812 [24], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0812 [25], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0812 [26], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0812 [27], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0812 [28], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0812 [29], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0812 [30], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0812 [31], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0812 [32], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0812 [33], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0812 [34], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0812 [35], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0812 [36], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0812 [37], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0812 [38], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0812 [39], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0812 [40], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0812 [41], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0812 [42], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0812 [43], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0812 [44], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0812 [45], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0812 [46], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0812 [47], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0811 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0811 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0811 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0811 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0811 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0811 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0811 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0811 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0811 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0811 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0811 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0811 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0811 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0811 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0811 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0811 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0811 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0811 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0811 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0811 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0811 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0811 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0811 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0811 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0811 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0811 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0811 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0811 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0811 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0811 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0811 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0811 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0811 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0811 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0811 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0811 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0811 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0811 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0811 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0811 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0811 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0811 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0811 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0811 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0811 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0811 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0811 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0811 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0811 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0811 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0811 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0811 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0811 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0811 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0811 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0811 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0811 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0811 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0811 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0811 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0811 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0811 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0811 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0811 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0811 [64], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0811 [65], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0811 [66], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0811 [67], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0811 [68], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0811 [69], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0811 [70], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0811 [71], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0811 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0811 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0811 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0811 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0811 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0811 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0811 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0811 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0811 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0811 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0811 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0811 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0811 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0811 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0811 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0811 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0811 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0811 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0811 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0811 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0811 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0811 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0811 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0811 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0811 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0811 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0811 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0811 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0811 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0811 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0811 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0811 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0811 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0811 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0811 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0811 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0811 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0811 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0811 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0811 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0811 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0811 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0811 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0811 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0811 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0811 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0811 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0811 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0811 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0811 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0811 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0811 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0811 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0811 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0811 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0811 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0810 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0810 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0810 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0810 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0810 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0810 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0810 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0810 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0810 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0810 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0810 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0810 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0810 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0810 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0810 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0810 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0810 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0810 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0810 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0810 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0810 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0810 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0810 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0810 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0810 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0810 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0810 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0810 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0810 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0810 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0810 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0810 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0810 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0810 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0810 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0810 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0810 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0810 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0810 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0810 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0810 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0810 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0810 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0810 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0810 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0810 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0810 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0810 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0810 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0810 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0810 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0810 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0810 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0810 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0810 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0810 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0810 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0810 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0810 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0810 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0810 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0810 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0810 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0810 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0809 [0], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0809 [1], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0809 [2], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0809 [3], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0809 [4], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0809 [5], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0809 [6], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0809 [7], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0809 [8], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0809 [9], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0809 [10], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0809 [11], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0809 [12], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0809 [13], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0809 [14], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0809 [15], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0809 [16], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0809 [17], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0809 [18], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0809 [19], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0809 [20], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0809 [21], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0809 [22], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0809 [23], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0809 [24], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0809 [25], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0809 [26], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0809 [27], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0809 [28], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0809 [29], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0809 [30], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0809 [31], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0809 [32], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0809 [33], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0809 [34], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0809 [35], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0809 [36], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0809 [37], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0809 [38], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0809 [39], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0809 [40], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0809 [41], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0809 [42], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0809 [43], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0809 [44], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0809 [45], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0809 [46], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0809 [47], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0809 [48], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0809 [49], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0809 [50], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0809 [51], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0809 [52], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0809 [53], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0809 [54], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0809 [55], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0808 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0808 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0808 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0808 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0808 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0808 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0808 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0808 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0808 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0808 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0808 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0808 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0808 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0808 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0808 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0808 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0808 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0808 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0808 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0808 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0808 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0808 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0808 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0808 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0808 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0808 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0808 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0808 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0808 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0808 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0808 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0808 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0808 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0808 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0808 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0808 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0808 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0808 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0808 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0808 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0808 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0808 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0808 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0808 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0808 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0808 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0808 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0808 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0808 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0808 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0808 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0808 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0808 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0808 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0808 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0808 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0808 [56], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0808 [57], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0808 [58], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0808 [59], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0808 [60], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0808 [61], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0808 [62], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0808 [63], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0808 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0808 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0808 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0808 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0808 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0808 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0808 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0808 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0808 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0808 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0808 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0808 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0808 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0808 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0808 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0808 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0808 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0808 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0808 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0808 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0808 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0808 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0808 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0808 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0808 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0808 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0808 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0808 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0808 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0808 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0808 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0808 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0808 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0808 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0808 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0808 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0808 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0808 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0808 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0808 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0808 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0808 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0808 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0808 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0808 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0808 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0808 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0808 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0808 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0808 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0808 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0808 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0808 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0808 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0808 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0808 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0808 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0808 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0808 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0808 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0808 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0808 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0808 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0808 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0807 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0807 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0807 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0807 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0807 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0807 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0807 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0807 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0807 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0807 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0807 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0807 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0807 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0807 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0807 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0807 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0807 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0807 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0807 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0807 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0807 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0807 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0807 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0807 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0807 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0807 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0807 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0807 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0807 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0807 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0807 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0807 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0807 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0807 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0807 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0807 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0807 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0807 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0807 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0807 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0807 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0807 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0807 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0807 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0807 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0807 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0807 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0807 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0807 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0807 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0807 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0807 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0807 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0807 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0807 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0807 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0806 [0], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0806 [1], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0806 [2], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0806 [3], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0806 [4], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0806 [5], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0806 [6], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0806 [7], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0806 [8], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0806 [9], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0806 [10], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0806 [11], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0806 [12], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0806 [13], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0806 [14], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0806 [15], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0806 [16], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0806 [17], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0806 [18], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0806 [19], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0806 [20], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0806 [21], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0806 [22], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0806 [23], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0806 [24], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0806 [25], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0806 [26], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0806 [27], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0806 [28], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0806 [29], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0806 [30], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0806 [31], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0806 [32], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0806 [33], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0806 [34], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0806 [35], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0806 [36], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0806 [37], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0806 [38], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0806 [39], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0806 [40], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0806 [41], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0806 [42], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0806 [43], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0806 [44], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0806 [45], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0806 [46], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0806 [47], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0806 [48], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0806 [49], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0806 [50], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0806 [51], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0806 [52], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0806 [53], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0806 [54], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0806 [55], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0806 [56], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0806 [57], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0806 [58], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0806 [59], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0806 [60], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0806 [61], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0806 [62], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0806 [63], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0365 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0365 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0365 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n0365 [3], \xm8051_golden_model_1.n0453 [3]);
  buf(\xm8051_golden_model_1.n0805 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0805 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0805 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0805 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0805 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0805 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0805 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0805 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0805 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0805 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0805 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0805 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0805 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0805 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0805 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0805 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0805 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0805 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0805 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0805 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0805 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0805 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0805 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0805 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0805 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0805 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0805 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0805 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0805 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0805 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0805 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0805 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0805 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0805 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0805 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0805 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0805 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0805 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0805 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0805 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0805 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0805 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0805 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0805 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0805 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0805 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0805 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0805 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0805 [48], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0805 [49], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0805 [50], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0805 [51], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0805 [52], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0805 [53], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0805 [54], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0805 [55], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0805 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0805 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0805 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0805 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0805 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0805 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0805 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0805 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0805 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0805 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0805 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0805 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0805 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0805 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0805 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0805 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0805 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0805 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0805 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0805 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0805 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0805 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0805 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0805 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0805 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0805 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0805 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0805 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0805 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0805 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0805 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0805 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0805 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0805 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0805 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0805 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0805 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0805 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0805 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0805 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0805 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0805 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0805 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0805 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0805 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0805 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0805 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0805 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0805 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0805 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0805 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0805 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0805 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0805 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0805 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0805 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0805 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0805 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0805 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0805 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0805 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0805 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0805 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0805 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0805 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0805 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0805 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0805 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0805 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0805 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0805 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0805 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0804 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0804 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0804 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0804 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0804 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0804 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0804 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0804 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0804 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0804 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0804 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0804 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0804 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0804 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0804 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0804 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0804 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0804 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0804 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0804 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0804 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0804 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0804 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0804 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0804 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0804 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0804 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0804 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0804 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0804 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0804 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0804 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0804 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0804 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0804 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0804 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0804 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0804 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0804 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0804 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0804 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0804 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0804 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0804 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0804 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0804 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0804 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0804 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0803 [0], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0803 [1], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0803 [2], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0803 [3], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0803 [4], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0803 [5], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0803 [6], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0803 [7], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0803 [8], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0803 [9], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0803 [10], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0803 [11], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0803 [12], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0803 [13], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0803 [14], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0803 [15], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0803 [16], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0803 [17], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0803 [18], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0803 [19], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0803 [20], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0803 [21], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0803 [22], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0803 [23], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0803 [24], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0803 [25], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0803 [26], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0803 [27], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0803 [28], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0803 [29], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0803 [30], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0803 [31], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0803 [32], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0803 [33], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0803 [34], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0803 [35], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0803 [36], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0803 [37], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0803 [38], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0803 [39], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0803 [40], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0803 [41], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0803 [42], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0803 [43], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0803 [44], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0803 [45], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0803 [46], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0803 [47], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0803 [48], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0803 [49], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0803 [50], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0803 [51], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0803 [52], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0803 [53], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0803 [54], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0803 [55], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0803 [56], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0803 [57], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0803 [58], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0803 [59], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0803 [60], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0803 [61], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0803 [62], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0803 [63], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0803 [64], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0803 [65], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0803 [66], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0803 [67], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0803 [68], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0803 [69], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0803 [70], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0803 [71], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0802 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0802 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0802 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0802 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0802 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0802 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0802 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0802 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0802 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0802 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0802 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0802 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0802 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0802 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0802 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0802 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0802 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0802 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0802 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0802 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0802 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0802 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0802 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0802 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0802 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0802 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0802 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0802 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0802 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0802 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0802 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0802 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0802 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0802 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0802 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0802 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0802 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0802 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0802 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0802 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0802 [40], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0802 [41], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0802 [42], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0802 [43], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0802 [44], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0802 [45], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0802 [46], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0802 [47], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0802 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0802 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0802 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0802 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0802 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0802 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0802 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0802 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0802 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0802 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0802 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0802 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0802 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0802 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0802 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0802 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0802 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0802 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0802 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0802 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0802 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0802 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0802 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0802 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0802 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0802 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0802 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0802 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0802 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0802 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0802 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0802 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0802 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0802 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0802 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0802 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0802 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0802 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0802 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0802 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0802 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0802 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0802 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0802 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0802 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0802 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0802 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0802 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0802 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0802 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0802 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0802 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0802 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0802 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0802 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0802 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0802 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0802 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0802 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0802 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0802 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0802 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0802 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0802 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0802 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0802 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0802 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0802 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0802 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0802 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0802 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0802 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0802 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0802 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0802 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0802 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0802 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0802 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0802 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0802 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0801 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0801 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0801 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0801 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0801 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0801 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0801 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0801 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0801 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0801 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0801 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0801 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0801 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0801 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0801 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0801 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0801 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0801 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0801 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0801 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0801 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0801 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0801 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0801 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0801 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0801 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0801 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0801 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0801 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0801 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0801 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0801 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0801 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0801 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0801 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0801 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0801 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0801 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0801 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0801 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0800 [0], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0800 [1], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0800 [2], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0800 [3], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0800 [4], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0800 [5], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0800 [6], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0800 [7], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0800 [8], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0800 [9], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0800 [10], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0800 [11], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0800 [12], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0800 [13], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0800 [14], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0800 [15], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0800 [16], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0800 [17], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0800 [18], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0800 [19], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0800 [20], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0800 [21], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0800 [22], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0800 [23], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0800 [24], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0800 [25], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0800 [26], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0800 [27], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0800 [28], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0800 [29], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0800 [30], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0800 [31], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0800 [32], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0800 [33], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0800 [34], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0800 [35], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0800 [36], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0800 [37], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0800 [38], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0800 [39], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0800 [40], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0800 [41], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0800 [42], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0800 [43], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0800 [44], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0800 [45], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0800 [46], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0800 [47], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0800 [48], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0800 [49], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0800 [50], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0800 [51], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0800 [52], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0800 [53], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0800 [54], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0800 [55], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0800 [56], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0800 [57], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0800 [58], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0800 [59], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0800 [60], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0800 [61], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0800 [62], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0800 [63], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0800 [64], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0800 [65], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0800 [66], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0800 [67], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0800 [68], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0800 [69], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0800 [70], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0800 [71], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0800 [72], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0800 [73], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0800 [74], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0800 [75], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0800 [76], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0800 [77], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0800 [78], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0800 [79], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0799 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0799 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0799 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0799 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0799 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0799 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0799 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0799 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0799 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0799 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0799 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0799 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0799 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0799 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0799 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0799 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0799 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0799 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0799 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0799 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0799 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0799 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0799 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0799 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0799 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0799 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0799 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0799 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0799 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0799 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0799 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0799 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0799 [32], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0799 [33], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0799 [34], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0799 [35], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0799 [36], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0799 [37], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0799 [38], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0799 [39], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0799 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0799 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0799 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0799 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0799 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0799 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0799 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0799 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0799 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0799 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0799 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0799 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0799 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0799 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0799 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0799 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0799 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0799 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0799 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0799 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0799 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0799 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0799 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0799 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0799 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0799 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0799 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0799 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0799 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0799 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0799 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0799 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0799 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0799 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0799 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0799 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0799 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0799 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0799 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0799 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0799 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0799 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0799 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0799 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0799 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0799 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0799 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0799 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0799 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0799 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0799 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0799 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0799 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0799 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0799 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0799 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0799 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0799 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0799 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0799 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0799 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0799 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0799 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0799 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0799 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0799 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0799 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0799 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0799 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0799 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0799 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0799 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0799 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0799 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0799 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0799 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0799 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0799 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0799 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0799 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0799 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0799 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0799 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0799 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0799 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0799 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0799 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0799 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0798 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0798 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0798 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0798 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0798 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0798 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0798 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0798 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0798 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0798 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0798 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0798 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0798 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0798 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0798 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0798 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0798 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0798 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0798 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0798 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0798 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0798 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0798 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0798 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0798 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0798 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0798 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0798 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0798 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0798 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0798 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0798 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0797 [0], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0797 [1], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0797 [2], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0797 [3], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0797 [4], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0797 [5], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0797 [6], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0797 [7], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0797 [8], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0797 [9], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0797 [10], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0797 [11], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0797 [12], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0797 [13], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0797 [14], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0797 [15], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0797 [16], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0797 [17], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0797 [18], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0797 [19], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0797 [20], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0797 [21], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0797 [22], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0797 [23], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0797 [24], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0797 [25], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0797 [26], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0797 [27], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0797 [28], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0797 [29], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0797 [30], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0797 [31], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0797 [32], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0797 [33], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0797 [34], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0797 [35], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0797 [36], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0797 [37], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0797 [38], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0797 [39], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0797 [40], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0797 [41], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0797 [42], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0797 [43], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0797 [44], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0797 [45], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0797 [46], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0797 [47], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0797 [48], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0797 [49], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0797 [50], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0797 [51], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0797 [52], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0797 [53], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0797 [54], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0797 [55], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0797 [56], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0797 [57], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0797 [58], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0797 [59], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0797 [60], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0797 [61], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0797 [62], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0797 [63], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0797 [64], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0797 [65], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0797 [66], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0797 [67], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0797 [68], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0797 [69], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0797 [70], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0797 [71], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0797 [72], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0797 [73], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0797 [74], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0797 [75], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0797 [76], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0797 [77], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0797 [78], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0797 [79], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0797 [80], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0797 [81], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0797 [82], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0797 [83], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0797 [84], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0797 [85], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0797 [86], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0797 [87], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0796 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0796 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0796 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0796 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0796 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0796 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0796 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0796 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0796 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0796 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0796 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0796 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0796 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0796 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0796 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0796 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0796 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0796 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0796 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0796 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0796 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0796 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0796 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0796 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0796 [24], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0796 [25], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0796 [26], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0796 [27], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0796 [28], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0796 [29], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0796 [30], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0796 [31], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0796 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0796 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0796 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0796 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0796 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0796 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0796 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0796 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0796 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0796 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0796 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0796 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0796 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0796 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0796 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0796 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0796 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0796 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0796 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0796 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0796 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0796 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0796 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0796 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0796 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0796 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0796 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0796 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0796 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0796 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0796 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0796 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0796 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0796 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0796 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0796 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0796 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0796 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0796 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0796 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0796 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0796 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0796 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0796 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0796 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0796 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0796 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0796 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0796 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0796 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0796 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0796 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0796 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0796 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0796 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0796 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0796 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0796 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0796 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0796 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0796 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0796 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0796 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0796 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0796 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0796 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0796 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0796 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0796 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0796 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0796 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0796 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0796 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0796 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0796 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0796 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0796 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0796 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0796 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0796 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0796 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0796 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0796 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0796 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0796 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0796 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0796 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0796 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0796 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0796 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0796 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0796 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0796 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0796 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0796 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0796 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0353 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0353 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0353 [2], \xm8051_golden_model_1.n0483 [2]);
  buf(\xm8051_golden_model_1.n0353 [3], \xm8051_golden_model_1.n0443 [3]);
  buf(\xm8051_golden_model_1.n0795 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0795 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0795 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0795 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0795 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0795 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0795 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0795 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0795 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0795 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0795 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0795 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0795 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0795 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0795 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0795 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0795 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0795 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0795 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0795 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0795 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0795 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0795 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0795 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0794 [0], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0794 [1], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0794 [2], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0794 [3], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0794 [4], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0794 [5], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0794 [6], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0794 [7], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0794 [8], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0794 [9], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0794 [10], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0794 [11], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0794 [12], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0794 [13], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0794 [14], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0794 [15], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0794 [16], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0794 [17], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0794 [18], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0794 [19], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0794 [20], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0794 [21], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0794 [22], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0794 [23], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0794 [24], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0794 [25], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0794 [26], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0794 [27], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0794 [28], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0794 [29], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0794 [30], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0794 [31], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0794 [32], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0794 [33], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0794 [34], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0794 [35], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0794 [36], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0794 [37], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0794 [38], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0794 [39], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0794 [40], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0794 [41], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0794 [42], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0794 [43], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0794 [44], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0794 [45], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0794 [46], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0794 [47], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0794 [48], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0794 [49], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0794 [50], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0794 [51], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0794 [52], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0794 [53], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0794 [54], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0794 [55], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0794 [56], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0794 [57], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0794 [58], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0794 [59], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0794 [60], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0794 [61], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0794 [62], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0794 [63], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0794 [64], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0794 [65], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0794 [66], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0794 [67], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0794 [68], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0794 [69], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0794 [70], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0794 [71], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0794 [72], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0794 [73], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0794 [74], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0794 [75], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0794 [76], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0794 [77], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0794 [78], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0794 [79], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0794 [80], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0794 [81], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0794 [82], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0794 [83], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0794 [84], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0794 [85], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0794 [86], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0794 [87], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0794 [88], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0794 [89], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0794 [90], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0794 [91], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0794 [92], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0794 [93], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0794 [94], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0794 [95], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0793 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0793 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0793 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0793 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0793 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0793 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0793 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0793 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0793 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0793 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0793 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0793 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0793 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0793 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0793 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0793 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0793 [16], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0793 [17], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0793 [18], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0793 [19], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0793 [20], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0793 [21], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0793 [22], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0793 [23], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0793 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0793 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0793 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0793 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0793 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0793 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0793 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0793 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0793 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0793 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0793 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0793 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0793 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0793 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0793 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0793 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0793 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0793 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0793 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0793 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0793 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0793 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0793 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0793 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0793 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0793 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0793 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0793 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0793 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0793 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0793 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0793 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0793 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0793 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0793 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0793 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0793 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0793 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0793 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0793 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0793 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0793 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0793 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0793 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0793 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0793 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0793 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0793 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0793 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0793 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0793 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0793 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0793 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0793 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0793 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0793 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0793 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0793 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0793 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0793 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0793 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0793 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0793 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0793 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0793 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0793 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0793 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0793 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0793 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0793 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0793 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0793 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0793 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0793 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0793 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0793 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0793 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0793 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0793 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0793 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0793 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0793 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0793 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0793 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0793 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0793 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0793 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0793 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0793 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0793 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0793 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0793 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0793 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0793 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0793 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0793 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0793 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0793 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0793 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0793 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0793 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0793 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0793 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0793 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0792 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0792 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0792 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0792 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0792 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0792 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0792 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0792 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0792 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0792 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0792 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0792 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0792 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0792 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0792 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0792 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0791 [0], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0791 [1], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0791 [2], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0791 [3], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0791 [4], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0791 [5], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0791 [6], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0791 [7], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0791 [8], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0791 [9], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0791 [10], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0791 [11], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0791 [12], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0791 [13], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0791 [14], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0791 [15], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0791 [16], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0791 [17], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0791 [18], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0791 [19], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0791 [20], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0791 [21], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0791 [22], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0791 [23], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0791 [24], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0791 [25], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0791 [26], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0791 [27], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0791 [28], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0791 [29], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0791 [30], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0791 [31], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0791 [32], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0791 [33], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0791 [34], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0791 [35], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0791 [36], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0791 [37], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0791 [38], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0791 [39], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0791 [40], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0791 [41], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0791 [42], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0791 [43], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0791 [44], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0791 [45], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0791 [46], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0791 [47], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0791 [48], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0791 [49], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0791 [50], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0791 [51], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0791 [52], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0791 [53], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0791 [54], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0791 [55], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0791 [56], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0791 [57], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0791 [58], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0791 [59], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0791 [60], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0791 [61], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0791 [62], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0791 [63], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0791 [64], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0791 [65], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0791 [66], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0791 [67], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0791 [68], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0791 [69], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0791 [70], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0791 [71], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0791 [72], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0791 [73], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0791 [74], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0791 [75], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0791 [76], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0791 [77], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0791 [78], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0791 [79], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0791 [80], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0791 [81], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0791 [82], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0791 [83], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0791 [84], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0791 [85], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0791 [86], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0791 [87], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0791 [88], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0791 [89], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0791 [90], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0791 [91], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0791 [92], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0791 [93], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0791 [94], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0791 [95], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0791 [96], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0791 [97], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0791 [98], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0791 [99], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0791 [100], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0791 [101], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0791 [102], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0791 [103], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0790 [0], \xm8051_golden_model_1.n0844 [0]);
  buf(\xm8051_golden_model_1.n0790 [1], \xm8051_golden_model_1.n0844 [1]);
  buf(\xm8051_golden_model_1.n0790 [2], \xm8051_golden_model_1.n0844 [2]);
  buf(\xm8051_golden_model_1.n0790 [3], \xm8051_golden_model_1.n0844 [3]);
  buf(\xm8051_golden_model_1.n0790 [4], \xm8051_golden_model_1.n0844 [4]);
  buf(\xm8051_golden_model_1.n0790 [5], \xm8051_golden_model_1.n0844 [5]);
  buf(\xm8051_golden_model_1.n0790 [6], \xm8051_golden_model_1.n0844 [6]);
  buf(\xm8051_golden_model_1.n0790 [7], \xm8051_golden_model_1.n0844 [7]);
  buf(\xm8051_golden_model_1.n0790 [8], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0790 [9], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0790 [10], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0790 [11], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0790 [12], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0790 [13], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0790 [14], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0790 [15], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0790 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0790 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0790 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0790 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0790 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0790 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0790 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0790 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0790 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0790 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0790 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0790 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0790 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0790 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0790 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0790 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0790 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0790 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0790 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0790 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0790 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0790 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0790 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0790 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0790 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0790 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0790 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0790 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0790 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0790 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0790 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0790 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0790 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0790 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0790 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0790 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0790 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0790 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0790 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0790 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0790 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0790 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0790 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0790 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0790 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0790 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0790 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0790 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0790 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0790 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0790 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0790 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0790 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0790 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0790 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0790 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0790 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0790 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0790 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0790 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0790 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0790 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0790 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0790 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0790 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0790 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0790 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0790 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0790 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0790 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0790 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0790 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0790 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0790 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0790 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0790 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0790 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0790 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0790 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0790 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0790 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0790 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0790 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0790 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0790 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0790 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0790 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0790 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0790 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0790 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0790 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0790 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0790 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0790 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0790 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0790 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0790 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0790 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0790 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0790 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0790 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0790 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0790 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0790 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0790 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0790 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0790 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0790 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0790 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0790 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0790 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0790 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0789 [0], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0789 [1], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0789 [2], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0789 [3], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0789 [4], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0789 [5], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0789 [6], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0789 [7], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0789 [8], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0789 [9], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0789 [10], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0789 [11], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0789 [12], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0789 [13], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0789 [14], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0789 [15], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0789 [16], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0789 [17], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0789 [18], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0789 [19], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0789 [20], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0789 [21], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0789 [22], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0789 [23], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0789 [24], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0789 [25], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0789 [26], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0789 [27], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0789 [28], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0789 [29], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0789 [30], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0789 [31], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0789 [32], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0789 [33], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0789 [34], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0789 [35], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0789 [36], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0789 [37], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0789 [38], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0789 [39], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0789 [40], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0789 [41], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0789 [42], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0789 [43], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0789 [44], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0789 [45], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0789 [46], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0789 [47], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0789 [48], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0789 [49], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0789 [50], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0789 [51], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0789 [52], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0789 [53], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0789 [54], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0789 [55], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0789 [56], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0789 [57], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0789 [58], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0789 [59], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0789 [60], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0789 [61], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0789 [62], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0789 [63], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0789 [64], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0789 [65], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0789 [66], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0789 [67], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0789 [68], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0789 [69], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0789 [70], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0789 [71], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0789 [72], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0789 [73], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0789 [74], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0789 [75], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0789 [76], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0789 [77], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0789 [78], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0789 [79], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0789 [80], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0789 [81], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0789 [82], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0789 [83], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0789 [84], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0789 [85], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0789 [86], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0789 [87], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0789 [88], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0789 [89], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0789 [90], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0789 [91], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0789 [92], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0789 [93], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0789 [94], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0789 [95], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0789 [96], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0789 [97], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0789 [98], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0789 [99], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0789 [100], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0789 [101], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0789 [102], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0789 [103], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0789 [104], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0789 [105], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0789 [106], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0789 [107], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0789 [108], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0789 [109], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0789 [110], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0789 [111], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n0788 [0], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0788 [1], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0788 [2], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0788 [3], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0788 [4], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0788 [5], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0788 [6], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0788 [7], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0788 [8], \xm8051_golden_model_1.n0843 [8]);
  buf(\xm8051_golden_model_1.n0788 [9], \xm8051_golden_model_1.n0843 [9]);
  buf(\xm8051_golden_model_1.n0788 [10], \xm8051_golden_model_1.n0843 [10]);
  buf(\xm8051_golden_model_1.n0788 [11], \xm8051_golden_model_1.n0843 [11]);
  buf(\xm8051_golden_model_1.n0788 [12], \xm8051_golden_model_1.n0843 [12]);
  buf(\xm8051_golden_model_1.n0788 [13], \xm8051_golden_model_1.n0843 [13]);
  buf(\xm8051_golden_model_1.n0788 [14], \xm8051_golden_model_1.n0843 [14]);
  buf(\xm8051_golden_model_1.n0788 [15], \xm8051_golden_model_1.n0843 [15]);
  buf(\xm8051_golden_model_1.n0788 [16], \xm8051_golden_model_1.n0842 [16]);
  buf(\xm8051_golden_model_1.n0788 [17], \xm8051_golden_model_1.n0842 [17]);
  buf(\xm8051_golden_model_1.n0788 [18], \xm8051_golden_model_1.n0842 [18]);
  buf(\xm8051_golden_model_1.n0788 [19], \xm8051_golden_model_1.n0842 [19]);
  buf(\xm8051_golden_model_1.n0788 [20], \xm8051_golden_model_1.n0842 [20]);
  buf(\xm8051_golden_model_1.n0788 [21], \xm8051_golden_model_1.n0842 [21]);
  buf(\xm8051_golden_model_1.n0788 [22], \xm8051_golden_model_1.n0842 [22]);
  buf(\xm8051_golden_model_1.n0788 [23], \xm8051_golden_model_1.n0842 [23]);
  buf(\xm8051_golden_model_1.n0788 [24], \xm8051_golden_model_1.n0841 [24]);
  buf(\xm8051_golden_model_1.n0788 [25], \xm8051_golden_model_1.n0841 [25]);
  buf(\xm8051_golden_model_1.n0788 [26], \xm8051_golden_model_1.n0841 [26]);
  buf(\xm8051_golden_model_1.n0788 [27], \xm8051_golden_model_1.n0841 [27]);
  buf(\xm8051_golden_model_1.n0788 [28], \xm8051_golden_model_1.n0841 [28]);
  buf(\xm8051_golden_model_1.n0788 [29], \xm8051_golden_model_1.n0841 [29]);
  buf(\xm8051_golden_model_1.n0788 [30], \xm8051_golden_model_1.n0841 [30]);
  buf(\xm8051_golden_model_1.n0788 [31], \xm8051_golden_model_1.n0841 [31]);
  buf(\xm8051_golden_model_1.n0788 [32], \xm8051_golden_model_1.n0840 [32]);
  buf(\xm8051_golden_model_1.n0788 [33], \xm8051_golden_model_1.n0840 [33]);
  buf(\xm8051_golden_model_1.n0788 [34], \xm8051_golden_model_1.n0840 [34]);
  buf(\xm8051_golden_model_1.n0788 [35], \xm8051_golden_model_1.n0840 [35]);
  buf(\xm8051_golden_model_1.n0788 [36], \xm8051_golden_model_1.n0840 [36]);
  buf(\xm8051_golden_model_1.n0788 [37], \xm8051_golden_model_1.n0840 [37]);
  buf(\xm8051_golden_model_1.n0788 [38], \xm8051_golden_model_1.n0840 [38]);
  buf(\xm8051_golden_model_1.n0788 [39], \xm8051_golden_model_1.n0840 [39]);
  buf(\xm8051_golden_model_1.n0788 [40], \xm8051_golden_model_1.n0839 [40]);
  buf(\xm8051_golden_model_1.n0788 [41], \xm8051_golden_model_1.n0839 [41]);
  buf(\xm8051_golden_model_1.n0788 [42], \xm8051_golden_model_1.n0839 [42]);
  buf(\xm8051_golden_model_1.n0788 [43], \xm8051_golden_model_1.n0839 [43]);
  buf(\xm8051_golden_model_1.n0788 [44], \xm8051_golden_model_1.n0839 [44]);
  buf(\xm8051_golden_model_1.n0788 [45], \xm8051_golden_model_1.n0839 [45]);
  buf(\xm8051_golden_model_1.n0788 [46], \xm8051_golden_model_1.n0839 [46]);
  buf(\xm8051_golden_model_1.n0788 [47], \xm8051_golden_model_1.n0839 [47]);
  buf(\xm8051_golden_model_1.n0788 [48], \xm8051_golden_model_1.n0838 [48]);
  buf(\xm8051_golden_model_1.n0788 [49], \xm8051_golden_model_1.n0838 [49]);
  buf(\xm8051_golden_model_1.n0788 [50], \xm8051_golden_model_1.n0838 [50]);
  buf(\xm8051_golden_model_1.n0788 [51], \xm8051_golden_model_1.n0838 [51]);
  buf(\xm8051_golden_model_1.n0788 [52], \xm8051_golden_model_1.n0838 [52]);
  buf(\xm8051_golden_model_1.n0788 [53], \xm8051_golden_model_1.n0838 [53]);
  buf(\xm8051_golden_model_1.n0788 [54], \xm8051_golden_model_1.n0838 [54]);
  buf(\xm8051_golden_model_1.n0788 [55], \xm8051_golden_model_1.n0838 [55]);
  buf(\xm8051_golden_model_1.n0788 [56], \xm8051_golden_model_1.n0837 [56]);
  buf(\xm8051_golden_model_1.n0788 [57], \xm8051_golden_model_1.n0837 [57]);
  buf(\xm8051_golden_model_1.n0788 [58], \xm8051_golden_model_1.n0837 [58]);
  buf(\xm8051_golden_model_1.n0788 [59], \xm8051_golden_model_1.n0837 [59]);
  buf(\xm8051_golden_model_1.n0788 [60], \xm8051_golden_model_1.n0837 [60]);
  buf(\xm8051_golden_model_1.n0788 [61], \xm8051_golden_model_1.n0837 [61]);
  buf(\xm8051_golden_model_1.n0788 [62], \xm8051_golden_model_1.n0837 [62]);
  buf(\xm8051_golden_model_1.n0788 [63], \xm8051_golden_model_1.n0837 [63]);
  buf(\xm8051_golden_model_1.n0788 [64], \xm8051_golden_model_1.n0836 [64]);
  buf(\xm8051_golden_model_1.n0788 [65], \xm8051_golden_model_1.n0836 [65]);
  buf(\xm8051_golden_model_1.n0788 [66], \xm8051_golden_model_1.n0836 [66]);
  buf(\xm8051_golden_model_1.n0788 [67], \xm8051_golden_model_1.n0836 [67]);
  buf(\xm8051_golden_model_1.n0788 [68], \xm8051_golden_model_1.n0836 [68]);
  buf(\xm8051_golden_model_1.n0788 [69], \xm8051_golden_model_1.n0836 [69]);
  buf(\xm8051_golden_model_1.n0788 [70], \xm8051_golden_model_1.n0836 [70]);
  buf(\xm8051_golden_model_1.n0788 [71], \xm8051_golden_model_1.n0836 [71]);
  buf(\xm8051_golden_model_1.n0788 [72], \xm8051_golden_model_1.n0835 [72]);
  buf(\xm8051_golden_model_1.n0788 [73], \xm8051_golden_model_1.n0835 [73]);
  buf(\xm8051_golden_model_1.n0788 [74], \xm8051_golden_model_1.n0835 [74]);
  buf(\xm8051_golden_model_1.n0788 [75], \xm8051_golden_model_1.n0835 [75]);
  buf(\xm8051_golden_model_1.n0788 [76], \xm8051_golden_model_1.n0835 [76]);
  buf(\xm8051_golden_model_1.n0788 [77], \xm8051_golden_model_1.n0835 [77]);
  buf(\xm8051_golden_model_1.n0788 [78], \xm8051_golden_model_1.n0835 [78]);
  buf(\xm8051_golden_model_1.n0788 [79], \xm8051_golden_model_1.n0835 [79]);
  buf(\xm8051_golden_model_1.n0788 [80], \xm8051_golden_model_1.n0834 [80]);
  buf(\xm8051_golden_model_1.n0788 [81], \xm8051_golden_model_1.n0834 [81]);
  buf(\xm8051_golden_model_1.n0788 [82], \xm8051_golden_model_1.n0834 [82]);
  buf(\xm8051_golden_model_1.n0788 [83], \xm8051_golden_model_1.n0834 [83]);
  buf(\xm8051_golden_model_1.n0788 [84], \xm8051_golden_model_1.n0834 [84]);
  buf(\xm8051_golden_model_1.n0788 [85], \xm8051_golden_model_1.n0834 [85]);
  buf(\xm8051_golden_model_1.n0788 [86], \xm8051_golden_model_1.n0834 [86]);
  buf(\xm8051_golden_model_1.n0788 [87], \xm8051_golden_model_1.n0834 [87]);
  buf(\xm8051_golden_model_1.n0788 [88], \xm8051_golden_model_1.n0833 [88]);
  buf(\xm8051_golden_model_1.n0788 [89], \xm8051_golden_model_1.n0833 [89]);
  buf(\xm8051_golden_model_1.n0788 [90], \xm8051_golden_model_1.n0833 [90]);
  buf(\xm8051_golden_model_1.n0788 [91], \xm8051_golden_model_1.n0833 [91]);
  buf(\xm8051_golden_model_1.n0788 [92], \xm8051_golden_model_1.n0833 [92]);
  buf(\xm8051_golden_model_1.n0788 [93], \xm8051_golden_model_1.n0833 [93]);
  buf(\xm8051_golden_model_1.n0788 [94], \xm8051_golden_model_1.n0833 [94]);
  buf(\xm8051_golden_model_1.n0788 [95], \xm8051_golden_model_1.n0833 [95]);
  buf(\xm8051_golden_model_1.n0788 [96], \xm8051_golden_model_1.n0832 [96]);
  buf(\xm8051_golden_model_1.n0788 [97], \xm8051_golden_model_1.n0832 [97]);
  buf(\xm8051_golden_model_1.n0788 [98], \xm8051_golden_model_1.n0832 [98]);
  buf(\xm8051_golden_model_1.n0788 [99], \xm8051_golden_model_1.n0832 [99]);
  buf(\xm8051_golden_model_1.n0788 [100], \xm8051_golden_model_1.n0832 [100]);
  buf(\xm8051_golden_model_1.n0788 [101], \xm8051_golden_model_1.n0832 [101]);
  buf(\xm8051_golden_model_1.n0788 [102], \xm8051_golden_model_1.n0832 [102]);
  buf(\xm8051_golden_model_1.n0788 [103], \xm8051_golden_model_1.n0832 [103]);
  buf(\xm8051_golden_model_1.n0788 [104], \xm8051_golden_model_1.n0831 [104]);
  buf(\xm8051_golden_model_1.n0788 [105], \xm8051_golden_model_1.n0831 [105]);
  buf(\xm8051_golden_model_1.n0788 [106], \xm8051_golden_model_1.n0831 [106]);
  buf(\xm8051_golden_model_1.n0788 [107], \xm8051_golden_model_1.n0831 [107]);
  buf(\xm8051_golden_model_1.n0788 [108], \xm8051_golden_model_1.n0831 [108]);
  buf(\xm8051_golden_model_1.n0788 [109], \xm8051_golden_model_1.n0831 [109]);
  buf(\xm8051_golden_model_1.n0788 [110], \xm8051_golden_model_1.n0831 [110]);
  buf(\xm8051_golden_model_1.n0788 [111], \xm8051_golden_model_1.n0831 [111]);
  buf(\xm8051_golden_model_1.n0788 [112], \xm8051_golden_model_1.n0830 [112]);
  buf(\xm8051_golden_model_1.n0788 [113], \xm8051_golden_model_1.n0830 [113]);
  buf(\xm8051_golden_model_1.n0788 [114], \xm8051_golden_model_1.n0830 [114]);
  buf(\xm8051_golden_model_1.n0788 [115], \xm8051_golden_model_1.n0830 [115]);
  buf(\xm8051_golden_model_1.n0788 [116], \xm8051_golden_model_1.n0830 [116]);
  buf(\xm8051_golden_model_1.n0788 [117], \xm8051_golden_model_1.n0830 [117]);
  buf(\xm8051_golden_model_1.n0788 [118], \xm8051_golden_model_1.n0830 [118]);
  buf(\xm8051_golden_model_1.n0788 [119], \xm8051_golden_model_1.n0830 [119]);
  buf(\xm8051_golden_model_1.n0788 [120], \xm8051_golden_model_1.n0828 [120]);
  buf(\xm8051_golden_model_1.n0788 [121], \xm8051_golden_model_1.n0828 [121]);
  buf(\xm8051_golden_model_1.n0788 [122], \xm8051_golden_model_1.n0828 [122]);
  buf(\xm8051_golden_model_1.n0788 [123], \xm8051_golden_model_1.n0828 [123]);
  buf(\xm8051_golden_model_1.n0788 [124], \xm8051_golden_model_1.n0828 [124]);
  buf(\xm8051_golden_model_1.n0788 [125], \xm8051_golden_model_1.n0828 [125]);
  buf(\xm8051_golden_model_1.n0788 [126], \xm8051_golden_model_1.n0828 [126]);
  buf(\xm8051_golden_model_1.n0788 [127], \xm8051_golden_model_1.n0828 [127]);
  buf(\xm8051_golden_model_1.n1281 [0], input_sha_func_41[0]);
  buf(\xm8051_golden_model_1.n1281 [1], input_sha_func_41[1]);
  buf(\xm8051_golden_model_1.n1281 [2], input_sha_func_41[2]);
  buf(\xm8051_golden_model_1.n1281 [3], input_sha_func_41[3]);
  buf(\xm8051_golden_model_1.n1281 [4], input_sha_func_41[4]);
  buf(\xm8051_golden_model_1.n1281 [5], input_sha_func_41[5]);
  buf(\xm8051_golden_model_1.n1281 [6], input_sha_func_41[6]);
  buf(\xm8051_golden_model_1.n1281 [7], input_sha_func_41[7]);
  buf(\xm8051_golden_model_1.n1281 [8], input_sha_func_41[8]);
  buf(\xm8051_golden_model_1.n1281 [9], input_sha_func_41[9]);
  buf(\xm8051_golden_model_1.n1281 [10], input_sha_func_41[10]);
  buf(\xm8051_golden_model_1.n1281 [11], input_sha_func_41[11]);
  buf(\xm8051_golden_model_1.n1281 [12], input_sha_func_41[12]);
  buf(\xm8051_golden_model_1.n1281 [13], input_sha_func_41[13]);
  buf(\xm8051_golden_model_1.n1281 [14], input_sha_func_41[14]);
  buf(\xm8051_golden_model_1.n1281 [15], input_sha_func_41[15]);
  buf(\xm8051_golden_model_1.n1281 [16], input_sha_func_41[16]);
  buf(\xm8051_golden_model_1.n1281 [17], input_sha_func_41[17]);
  buf(\xm8051_golden_model_1.n1281 [18], input_sha_func_41[18]);
  buf(\xm8051_golden_model_1.n1281 [19], input_sha_func_41[19]);
  buf(\xm8051_golden_model_1.n1281 [20], input_sha_func_41[20]);
  buf(\xm8051_golden_model_1.n1281 [21], input_sha_func_41[21]);
  buf(\xm8051_golden_model_1.n1281 [22], input_sha_func_41[22]);
  buf(\xm8051_golden_model_1.n1281 [23], input_sha_func_41[23]);
  buf(\xm8051_golden_model_1.n1281 [24], input_sha_func_41[24]);
  buf(\xm8051_golden_model_1.n1281 [25], input_sha_func_41[25]);
  buf(\xm8051_golden_model_1.n1281 [26], input_sha_func_41[26]);
  buf(\xm8051_golden_model_1.n1281 [27], input_sha_func_41[27]);
  buf(\xm8051_golden_model_1.n1281 [28], input_sha_func_41[28]);
  buf(\xm8051_golden_model_1.n1281 [29], input_sha_func_41[29]);
  buf(\xm8051_golden_model_1.n1281 [30], input_sha_func_41[30]);
  buf(\xm8051_golden_model_1.n1281 [31], input_sha_func_41[31]);
  buf(\xm8051_golden_model_1.n1281 [32], input_sha_func_40[0]);
  buf(\xm8051_golden_model_1.n1281 [33], input_sha_func_40[1]);
  buf(\xm8051_golden_model_1.n1281 [34], input_sha_func_40[2]);
  buf(\xm8051_golden_model_1.n1281 [35], input_sha_func_40[3]);
  buf(\xm8051_golden_model_1.n1281 [36], input_sha_func_40[4]);
  buf(\xm8051_golden_model_1.n1281 [37], input_sha_func_40[5]);
  buf(\xm8051_golden_model_1.n1281 [38], input_sha_func_40[6]);
  buf(\xm8051_golden_model_1.n1281 [39], input_sha_func_40[7]);
  buf(\xm8051_golden_model_1.n1281 [40], input_sha_func_40[8]);
  buf(\xm8051_golden_model_1.n1281 [41], input_sha_func_40[9]);
  buf(\xm8051_golden_model_1.n1281 [42], input_sha_func_40[10]);
  buf(\xm8051_golden_model_1.n1281 [43], input_sha_func_40[11]);
  buf(\xm8051_golden_model_1.n1281 [44], input_sha_func_40[12]);
  buf(\xm8051_golden_model_1.n1281 [45], input_sha_func_40[13]);
  buf(\xm8051_golden_model_1.n1281 [46], input_sha_func_40[14]);
  buf(\xm8051_golden_model_1.n1281 [47], input_sha_func_40[15]);
  buf(\xm8051_golden_model_1.n1281 [48], input_sha_func_40[16]);
  buf(\xm8051_golden_model_1.n1281 [49], input_sha_func_40[17]);
  buf(\xm8051_golden_model_1.n1281 [50], input_sha_func_40[18]);
  buf(\xm8051_golden_model_1.n1281 [51], input_sha_func_40[19]);
  buf(\xm8051_golden_model_1.n1281 [52], input_sha_func_40[20]);
  buf(\xm8051_golden_model_1.n1281 [53], input_sha_func_40[21]);
  buf(\xm8051_golden_model_1.n1281 [54], input_sha_func_40[22]);
  buf(\xm8051_golden_model_1.n1281 [55], input_sha_func_40[23]);
  buf(\xm8051_golden_model_1.n1281 [56], input_sha_func_40[24]);
  buf(\xm8051_golden_model_1.n1281 [57], input_sha_func_40[25]);
  buf(\xm8051_golden_model_1.n1281 [58], input_sha_func_40[26]);
  buf(\xm8051_golden_model_1.n1281 [59], input_sha_func_40[27]);
  buf(\xm8051_golden_model_1.n1281 [60], input_sha_func_40[28]);
  buf(\xm8051_golden_model_1.n1281 [61], input_sha_func_40[29]);
  buf(\xm8051_golden_model_1.n1281 [62], input_sha_func_40[30]);
  buf(\xm8051_golden_model_1.n1281 [63], input_sha_func_40[31]);
  buf(\xm8051_golden_model_1.n1281 [64], input_sha_func_40[32]);
  buf(\xm8051_golden_model_1.n1281 [65], input_sha_func_40[33]);
  buf(\xm8051_golden_model_1.n1281 [66], input_sha_func_40[34]);
  buf(\xm8051_golden_model_1.n1281 [67], input_sha_func_40[35]);
  buf(\xm8051_golden_model_1.n1281 [68], input_sha_func_40[36]);
  buf(\xm8051_golden_model_1.n1281 [69], input_sha_func_40[37]);
  buf(\xm8051_golden_model_1.n1281 [70], input_sha_func_40[38]);
  buf(\xm8051_golden_model_1.n1281 [71], input_sha_func_40[39]);
  buf(\xm8051_golden_model_1.n1281 [72], input_sha_func_40[40]);
  buf(\xm8051_golden_model_1.n1281 [73], input_sha_func_40[41]);
  buf(\xm8051_golden_model_1.n1281 [74], input_sha_func_40[42]);
  buf(\xm8051_golden_model_1.n1281 [75], input_sha_func_40[43]);
  buf(\xm8051_golden_model_1.n1281 [76], input_sha_func_40[44]);
  buf(\xm8051_golden_model_1.n1281 [77], input_sha_func_40[45]);
  buf(\xm8051_golden_model_1.n1281 [78], input_sha_func_40[46]);
  buf(\xm8051_golden_model_1.n1281 [79], input_sha_func_40[47]);
  buf(\xm8051_golden_model_1.n1281 [80], input_sha_func_40[48]);
  buf(\xm8051_golden_model_1.n1281 [81], input_sha_func_40[49]);
  buf(\xm8051_golden_model_1.n1281 [82], input_sha_func_40[50]);
  buf(\xm8051_golden_model_1.n1281 [83], input_sha_func_40[51]);
  buf(\xm8051_golden_model_1.n1281 [84], input_sha_func_40[52]);
  buf(\xm8051_golden_model_1.n1281 [85], input_sha_func_40[53]);
  buf(\xm8051_golden_model_1.n1281 [86], input_sha_func_40[54]);
  buf(\xm8051_golden_model_1.n1281 [87], input_sha_func_40[55]);
  buf(\xm8051_golden_model_1.n1281 [88], input_sha_func_40[56]);
  buf(\xm8051_golden_model_1.n1281 [89], input_sha_func_40[57]);
  buf(\xm8051_golden_model_1.n1281 [90], input_sha_func_40[58]);
  buf(\xm8051_golden_model_1.n1281 [91], input_sha_func_40[59]);
  buf(\xm8051_golden_model_1.n1281 [92], input_sha_func_40[60]);
  buf(\xm8051_golden_model_1.n1281 [93], input_sha_func_40[61]);
  buf(\xm8051_golden_model_1.n1281 [94], input_sha_func_40[62]);
  buf(\xm8051_golden_model_1.n1281 [95], input_sha_func_40[63]);
  buf(\xm8051_golden_model_1.n1281 [96], input_sha_func_39[0]);
  buf(\xm8051_golden_model_1.n1281 [97], input_sha_func_39[1]);
  buf(\xm8051_golden_model_1.n1281 [98], input_sha_func_39[2]);
  buf(\xm8051_golden_model_1.n1281 [99], input_sha_func_39[3]);
  buf(\xm8051_golden_model_1.n1281 [100], input_sha_func_39[4]);
  buf(\xm8051_golden_model_1.n1281 [101], input_sha_func_39[5]);
  buf(\xm8051_golden_model_1.n1281 [102], input_sha_func_39[6]);
  buf(\xm8051_golden_model_1.n1281 [103], input_sha_func_39[7]);
  buf(\xm8051_golden_model_1.n1281 [104], input_sha_func_39[8]);
  buf(\xm8051_golden_model_1.n1281 [105], input_sha_func_39[9]);
  buf(\xm8051_golden_model_1.n1281 [106], input_sha_func_39[10]);
  buf(\xm8051_golden_model_1.n1281 [107], input_sha_func_39[11]);
  buf(\xm8051_golden_model_1.n1281 [108], input_sha_func_39[12]);
  buf(\xm8051_golden_model_1.n1281 [109], input_sha_func_39[13]);
  buf(\xm8051_golden_model_1.n1281 [110], input_sha_func_39[14]);
  buf(\xm8051_golden_model_1.n1281 [111], input_sha_func_39[15]);
  buf(\xm8051_golden_model_1.n1281 [112], input_sha_func_39[16]);
  buf(\xm8051_golden_model_1.n1281 [113], input_sha_func_39[17]);
  buf(\xm8051_golden_model_1.n1281 [114], input_sha_func_39[18]);
  buf(\xm8051_golden_model_1.n1281 [115], input_sha_func_39[19]);
  buf(\xm8051_golden_model_1.n1281 [116], input_sha_func_39[20]);
  buf(\xm8051_golden_model_1.n1281 [117], input_sha_func_39[21]);
  buf(\xm8051_golden_model_1.n1281 [118], input_sha_func_39[22]);
  buf(\xm8051_golden_model_1.n1281 [119], input_sha_func_39[23]);
  buf(\xm8051_golden_model_1.n1281 [120], input_sha_func_39[24]);
  buf(\xm8051_golden_model_1.n1281 [121], input_sha_func_39[25]);
  buf(\xm8051_golden_model_1.n1281 [122], input_sha_func_39[26]);
  buf(\xm8051_golden_model_1.n1281 [123], input_sha_func_39[27]);
  buf(\xm8051_golden_model_1.n1281 [124], input_sha_func_39[28]);
  buf(\xm8051_golden_model_1.n1281 [125], input_sha_func_39[29]);
  buf(\xm8051_golden_model_1.n1281 [126], input_sha_func_39[30]);
  buf(\xm8051_golden_model_1.n1281 [127], input_sha_func_39[31]);
  buf(\xm8051_golden_model_1.n1281 [128], input_sha_func_39[32]);
  buf(\xm8051_golden_model_1.n1281 [129], input_sha_func_39[33]);
  buf(\xm8051_golden_model_1.n1281 [130], input_sha_func_39[34]);
  buf(\xm8051_golden_model_1.n1281 [131], input_sha_func_39[35]);
  buf(\xm8051_golden_model_1.n1281 [132], input_sha_func_39[36]);
  buf(\xm8051_golden_model_1.n1281 [133], input_sha_func_39[37]);
  buf(\xm8051_golden_model_1.n1281 [134], input_sha_func_39[38]);
  buf(\xm8051_golden_model_1.n1281 [135], input_sha_func_39[39]);
  buf(\xm8051_golden_model_1.n1281 [136], input_sha_func_39[40]);
  buf(\xm8051_golden_model_1.n1281 [137], input_sha_func_39[41]);
  buf(\xm8051_golden_model_1.n1281 [138], input_sha_func_39[42]);
  buf(\xm8051_golden_model_1.n1281 [139], input_sha_func_39[43]);
  buf(\xm8051_golden_model_1.n1281 [140], input_sha_func_39[44]);
  buf(\xm8051_golden_model_1.n1281 [141], input_sha_func_39[45]);
  buf(\xm8051_golden_model_1.n1281 [142], input_sha_func_39[46]);
  buf(\xm8051_golden_model_1.n1281 [143], input_sha_func_39[47]);
  buf(\xm8051_golden_model_1.n1281 [144], input_sha_func_39[48]);
  buf(\xm8051_golden_model_1.n1281 [145], input_sha_func_39[49]);
  buf(\xm8051_golden_model_1.n1281 [146], input_sha_func_39[50]);
  buf(\xm8051_golden_model_1.n1281 [147], input_sha_func_39[51]);
  buf(\xm8051_golden_model_1.n1281 [148], input_sha_func_39[52]);
  buf(\xm8051_golden_model_1.n1281 [149], input_sha_func_39[53]);
  buf(\xm8051_golden_model_1.n1281 [150], input_sha_func_39[54]);
  buf(\xm8051_golden_model_1.n1281 [151], input_sha_func_39[55]);
  buf(\xm8051_golden_model_1.n1281 [152], input_sha_func_39[56]);
  buf(\xm8051_golden_model_1.n1281 [153], input_sha_func_39[57]);
  buf(\xm8051_golden_model_1.n1281 [154], input_sha_func_39[58]);
  buf(\xm8051_golden_model_1.n1281 [155], input_sha_func_39[59]);
  buf(\xm8051_golden_model_1.n1281 [156], input_sha_func_39[60]);
  buf(\xm8051_golden_model_1.n1281 [157], input_sha_func_39[61]);
  buf(\xm8051_golden_model_1.n1281 [158], input_sha_func_39[62]);
  buf(\xm8051_golden_model_1.n1281 [159], input_sha_func_39[63]);
  buf(\xm8051_golden_model_1.n0341 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0341 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0341 [2], \xm8051_golden_model_1.n0473 [2]);
  buf(\xm8051_golden_model_1.n0341 [3], \xm8051_golden_model_1.n0433 [3]);
  buf(\xm8051_golden_model_1.n0783 [0], \xm8051_golden_model_1.sha_len [0]);
  buf(\xm8051_golden_model_1.n0783 [1], \xm8051_golden_model_1.sha_len [1]);
  buf(\xm8051_golden_model_1.n0783 [2], \xm8051_golden_model_1.sha_len [2]);
  buf(\xm8051_golden_model_1.n0783 [3], \xm8051_golden_model_1.sha_len [3]);
  buf(\xm8051_golden_model_1.n0783 [4], \xm8051_golden_model_1.sha_len [4]);
  buf(\xm8051_golden_model_1.n0783 [5], \xm8051_golden_model_1.sha_len [5]);
  buf(\xm8051_golden_model_1.n0783 [6], \xm8051_golden_model_1.sha_len [6]);
  buf(\xm8051_golden_model_1.n0783 [7], \xm8051_golden_model_1.sha_len [7]);
  buf(\xm8051_golden_model_1.n0783 [8], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0783 [9], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0783 [10], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0783 [11], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0783 [12], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0783 [13], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0783 [14], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0783 [15], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0782 [0], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0782 [1], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0782 [2], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0782 [3], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0782 [4], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0782 [5], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0782 [6], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0782 [7], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0782 [8], \xm8051_golden_model_1.sha_len [8]);
  buf(\xm8051_golden_model_1.n0782 [9], \xm8051_golden_model_1.sha_len [9]);
  buf(\xm8051_golden_model_1.n0782 [10], \xm8051_golden_model_1.sha_len [10]);
  buf(\xm8051_golden_model_1.n0782 [11], \xm8051_golden_model_1.sha_len [11]);
  buf(\xm8051_golden_model_1.n0782 [12], \xm8051_golden_model_1.sha_len [12]);
  buf(\xm8051_golden_model_1.n0782 [13], \xm8051_golden_model_1.sha_len [13]);
  buf(\xm8051_golden_model_1.n0782 [14], \xm8051_golden_model_1.sha_len [14]);
  buf(\xm8051_golden_model_1.n0782 [15], \xm8051_golden_model_1.sha_len [15]);
  buf(\xm8051_golden_model_1.n0329 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0329 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0329 [2], \xm8051_golden_model_1.n0463 [2]);
  buf(\xm8051_golden_model_1.n0329 [3], \xm8051_golden_model_1.n0423 [3]);
  buf(\xm8051_golden_model_1.n1279 [0], input_aes_func_38[0]);
  buf(\xm8051_golden_model_1.n1279 [1], input_aes_func_38[1]);
  buf(\xm8051_golden_model_1.n1279 [2], input_aes_func_38[2]);
  buf(\xm8051_golden_model_1.n1279 [3], input_aes_func_38[3]);
  buf(\xm8051_golden_model_1.n1279 [4], input_aes_func_38[4]);
  buf(\xm8051_golden_model_1.n1279 [5], input_aes_func_38[5]);
  buf(\xm8051_golden_model_1.n1279 [6], input_aes_func_38[6]);
  buf(\xm8051_golden_model_1.n1279 [7], input_aes_func_38[7]);
  buf(\xm8051_golden_model_1.n1279 [8], input_aes_func_38[8]);
  buf(\xm8051_golden_model_1.n1279 [9], input_aes_func_38[9]);
  buf(\xm8051_golden_model_1.n1279 [10], input_aes_func_38[10]);
  buf(\xm8051_golden_model_1.n1279 [11], input_aes_func_38[11]);
  buf(\xm8051_golden_model_1.n1279 [12], input_aes_func_38[12]);
  buf(\xm8051_golden_model_1.n1279 [13], input_aes_func_38[13]);
  buf(\xm8051_golden_model_1.n1279 [14], input_aes_func_38[14]);
  buf(\xm8051_golden_model_1.n1279 [15], input_aes_func_38[15]);
  buf(\xm8051_golden_model_1.n1279 [16], input_aes_func_38[16]);
  buf(\xm8051_golden_model_1.n1279 [17], input_aes_func_38[17]);
  buf(\xm8051_golden_model_1.n1279 [18], input_aes_func_38[18]);
  buf(\xm8051_golden_model_1.n1279 [19], input_aes_func_38[19]);
  buf(\xm8051_golden_model_1.n1279 [20], input_aes_func_38[20]);
  buf(\xm8051_golden_model_1.n1279 [21], input_aes_func_38[21]);
  buf(\xm8051_golden_model_1.n1279 [22], input_aes_func_38[22]);
  buf(\xm8051_golden_model_1.n1279 [23], input_aes_func_38[23]);
  buf(\xm8051_golden_model_1.n1279 [24], input_aes_func_38[24]);
  buf(\xm8051_golden_model_1.n1279 [25], input_aes_func_38[25]);
  buf(\xm8051_golden_model_1.n1279 [26], input_aes_func_38[26]);
  buf(\xm8051_golden_model_1.n1279 [27], input_aes_func_38[27]);
  buf(\xm8051_golden_model_1.n1279 [28], input_aes_func_38[28]);
  buf(\xm8051_golden_model_1.n1279 [29], input_aes_func_38[29]);
  buf(\xm8051_golden_model_1.n1279 [30], input_aes_func_38[30]);
  buf(\xm8051_golden_model_1.n1279 [31], input_aes_func_38[31]);
  buf(\xm8051_golden_model_1.n1279 [32], input_aes_func_38[32]);
  buf(\xm8051_golden_model_1.n1279 [33], input_aes_func_38[33]);
  buf(\xm8051_golden_model_1.n1279 [34], input_aes_func_38[34]);
  buf(\xm8051_golden_model_1.n1279 [35], input_aes_func_38[35]);
  buf(\xm8051_golden_model_1.n1279 [36], input_aes_func_38[36]);
  buf(\xm8051_golden_model_1.n1279 [37], input_aes_func_38[37]);
  buf(\xm8051_golden_model_1.n1279 [38], input_aes_func_38[38]);
  buf(\xm8051_golden_model_1.n1279 [39], input_aes_func_38[39]);
  buf(\xm8051_golden_model_1.n1279 [40], input_aes_func_38[40]);
  buf(\xm8051_golden_model_1.n1279 [41], input_aes_func_38[41]);
  buf(\xm8051_golden_model_1.n1279 [42], input_aes_func_38[42]);
  buf(\xm8051_golden_model_1.n1279 [43], input_aes_func_38[43]);
  buf(\xm8051_golden_model_1.n1279 [44], input_aes_func_38[44]);
  buf(\xm8051_golden_model_1.n1279 [45], input_aes_func_38[45]);
  buf(\xm8051_golden_model_1.n1279 [46], input_aes_func_38[46]);
  buf(\xm8051_golden_model_1.n1279 [47], input_aes_func_38[47]);
  buf(\xm8051_golden_model_1.n1279 [48], input_aes_func_38[48]);
  buf(\xm8051_golden_model_1.n1279 [49], input_aes_func_38[49]);
  buf(\xm8051_golden_model_1.n1279 [50], input_aes_func_38[50]);
  buf(\xm8051_golden_model_1.n1279 [51], input_aes_func_38[51]);
  buf(\xm8051_golden_model_1.n1279 [52], input_aes_func_38[52]);
  buf(\xm8051_golden_model_1.n1279 [53], input_aes_func_38[53]);
  buf(\xm8051_golden_model_1.n1279 [54], input_aes_func_38[54]);
  buf(\xm8051_golden_model_1.n1279 [55], input_aes_func_38[55]);
  buf(\xm8051_golden_model_1.n1279 [56], input_aes_func_38[56]);
  buf(\xm8051_golden_model_1.n1279 [57], input_aes_func_38[57]);
  buf(\xm8051_golden_model_1.n1279 [58], input_aes_func_38[58]);
  buf(\xm8051_golden_model_1.n1279 [59], input_aes_func_38[59]);
  buf(\xm8051_golden_model_1.n1279 [60], input_aes_func_38[60]);
  buf(\xm8051_golden_model_1.n1279 [61], input_aes_func_38[61]);
  buf(\xm8051_golden_model_1.n1279 [62], input_aes_func_38[62]);
  buf(\xm8051_golden_model_1.n1279 [63], input_aes_func_38[63]);
  buf(\xm8051_golden_model_1.n1279 [64], input_aes_func_37[0]);
  buf(\xm8051_golden_model_1.n1279 [65], input_aes_func_37[1]);
  buf(\xm8051_golden_model_1.n1279 [66], input_aes_func_37[2]);
  buf(\xm8051_golden_model_1.n1279 [67], input_aes_func_37[3]);
  buf(\xm8051_golden_model_1.n1279 [68], input_aes_func_37[4]);
  buf(\xm8051_golden_model_1.n1279 [69], input_aes_func_37[5]);
  buf(\xm8051_golden_model_1.n1279 [70], input_aes_func_37[6]);
  buf(\xm8051_golden_model_1.n1279 [71], input_aes_func_37[7]);
  buf(\xm8051_golden_model_1.n1279 [72], input_aes_func_37[8]);
  buf(\xm8051_golden_model_1.n1279 [73], input_aes_func_37[9]);
  buf(\xm8051_golden_model_1.n1279 [74], input_aes_func_37[10]);
  buf(\xm8051_golden_model_1.n1279 [75], input_aes_func_37[11]);
  buf(\xm8051_golden_model_1.n1279 [76], input_aes_func_37[12]);
  buf(\xm8051_golden_model_1.n1279 [77], input_aes_func_37[13]);
  buf(\xm8051_golden_model_1.n1279 [78], input_aes_func_37[14]);
  buf(\xm8051_golden_model_1.n1279 [79], input_aes_func_37[15]);
  buf(\xm8051_golden_model_1.n1279 [80], input_aes_func_37[16]);
  buf(\xm8051_golden_model_1.n1279 [81], input_aes_func_37[17]);
  buf(\xm8051_golden_model_1.n1279 [82], input_aes_func_37[18]);
  buf(\xm8051_golden_model_1.n1279 [83], input_aes_func_37[19]);
  buf(\xm8051_golden_model_1.n1279 [84], input_aes_func_37[20]);
  buf(\xm8051_golden_model_1.n1279 [85], input_aes_func_37[21]);
  buf(\xm8051_golden_model_1.n1279 [86], input_aes_func_37[22]);
  buf(\xm8051_golden_model_1.n1279 [87], input_aes_func_37[23]);
  buf(\xm8051_golden_model_1.n1279 [88], input_aes_func_37[24]);
  buf(\xm8051_golden_model_1.n1279 [89], input_aes_func_37[25]);
  buf(\xm8051_golden_model_1.n1279 [90], input_aes_func_37[26]);
  buf(\xm8051_golden_model_1.n1279 [91], input_aes_func_37[27]);
  buf(\xm8051_golden_model_1.n1279 [92], input_aes_func_37[28]);
  buf(\xm8051_golden_model_1.n1279 [93], input_aes_func_37[29]);
  buf(\xm8051_golden_model_1.n1279 [94], input_aes_func_37[30]);
  buf(\xm8051_golden_model_1.n1279 [95], input_aes_func_37[31]);
  buf(\xm8051_golden_model_1.n1279 [96], input_aes_func_37[32]);
  buf(\xm8051_golden_model_1.n1279 [97], input_aes_func_37[33]);
  buf(\xm8051_golden_model_1.n1279 [98], input_aes_func_37[34]);
  buf(\xm8051_golden_model_1.n1279 [99], input_aes_func_37[35]);
  buf(\xm8051_golden_model_1.n1279 [100], input_aes_func_37[36]);
  buf(\xm8051_golden_model_1.n1279 [101], input_aes_func_37[37]);
  buf(\xm8051_golden_model_1.n1279 [102], input_aes_func_37[38]);
  buf(\xm8051_golden_model_1.n1279 [103], input_aes_func_37[39]);
  buf(\xm8051_golden_model_1.n1279 [104], input_aes_func_37[40]);
  buf(\xm8051_golden_model_1.n1279 [105], input_aes_func_37[41]);
  buf(\xm8051_golden_model_1.n1279 [106], input_aes_func_37[42]);
  buf(\xm8051_golden_model_1.n1279 [107], input_aes_func_37[43]);
  buf(\xm8051_golden_model_1.n1279 [108], input_aes_func_37[44]);
  buf(\xm8051_golden_model_1.n1279 [109], input_aes_func_37[45]);
  buf(\xm8051_golden_model_1.n1279 [110], input_aes_func_37[46]);
  buf(\xm8051_golden_model_1.n1279 [111], input_aes_func_37[47]);
  buf(\xm8051_golden_model_1.n1279 [112], input_aes_func_37[48]);
  buf(\xm8051_golden_model_1.n1279 [113], input_aes_func_37[49]);
  buf(\xm8051_golden_model_1.n1279 [114], input_aes_func_37[50]);
  buf(\xm8051_golden_model_1.n1279 [115], input_aes_func_37[51]);
  buf(\xm8051_golden_model_1.n1279 [116], input_aes_func_37[52]);
  buf(\xm8051_golden_model_1.n1279 [117], input_aes_func_37[53]);
  buf(\xm8051_golden_model_1.n1279 [118], input_aes_func_37[54]);
  buf(\xm8051_golden_model_1.n1279 [119], input_aes_func_37[55]);
  buf(\xm8051_golden_model_1.n1279 [120], input_aes_func_37[56]);
  buf(\xm8051_golden_model_1.n1279 [121], input_aes_func_37[57]);
  buf(\xm8051_golden_model_1.n1279 [122], input_aes_func_37[58]);
  buf(\xm8051_golden_model_1.n1279 [123], input_aes_func_37[59]);
  buf(\xm8051_golden_model_1.n1279 [124], input_aes_func_37[60]);
  buf(\xm8051_golden_model_1.n1279 [125], input_aes_func_37[61]);
  buf(\xm8051_golden_model_1.n1279 [126], input_aes_func_37[62]);
  buf(\xm8051_golden_model_1.n1279 [127], input_aes_func_37[63]);
  buf(\xm8051_golden_model_1.n0775 , proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0317 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0317 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0317 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n0317 [3], \xm8051_golden_model_1.sha_bytes_processed [3]);
  buf(\xm8051_golden_model_1.n0317 [4], \xm8051_golden_model_1.sha_bytes_processed [4]);
  buf(\xm8051_golden_model_1.n0758 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0758 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0758 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0758 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0758 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0758 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0758 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0758 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0758 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0758 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0758 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0758 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0758 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0758 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0758 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0758 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0758 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0758 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0758 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0758 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0758 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0758 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0758 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0758 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0758 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0758 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0758 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0758 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0758 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0758 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0758 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0758 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0758 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0758 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0758 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0758 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0758 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0758 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0758 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0758 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0758 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0758 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0758 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0758 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0758 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0758 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0758 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0758 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0758 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0758 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0758 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0758 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0758 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0758 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0758 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0758 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0758 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0758 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0758 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0758 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0758 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0758 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0758 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0758 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0758 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0758 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0758 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0758 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0758 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0758 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0758 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0758 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0758 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0758 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0758 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0758 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0758 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0758 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0758 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0758 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0758 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0758 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0758 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0758 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0758 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0758 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0758 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0758 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0758 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0758 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0758 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0758 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0758 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0758 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0758 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0758 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0758 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0758 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0758 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0758 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0758 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0758 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0758 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0758 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0758 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0758 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0758 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0758 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0758 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0758 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0758 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0758 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0758 [120], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0758 [121], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0758 [122], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0758 [123], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0758 [124], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0758 [125], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0758 [126], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0758 [127], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0757 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0757 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0757 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0757 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0757 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0757 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0757 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0757 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0757 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0757 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0757 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0757 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0757 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0757 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0757 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0757 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0757 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0757 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0757 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0757 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0757 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0757 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0757 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0757 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0757 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0757 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0757 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0757 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0757 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0757 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0757 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0757 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0757 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0757 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0757 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0757 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0757 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0757 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0757 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0757 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0757 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0757 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0757 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0757 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0757 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0757 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0757 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0757 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0757 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0757 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0757 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0757 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0757 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0757 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0757 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0757 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0757 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0757 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0757 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0757 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0757 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0757 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0757 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0757 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0757 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0757 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0757 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0757 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0757 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0757 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0757 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0757 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0757 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0757 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0757 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0757 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0757 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0757 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0757 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0757 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0757 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0757 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0757 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0757 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0757 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0757 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0757 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0757 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0757 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0757 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0757 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0757 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0757 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0757 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0757 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0757 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0757 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0757 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0757 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0757 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0757 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0757 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0757 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0757 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0757 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0757 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0757 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0757 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0757 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0757 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0757 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0757 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0757 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0757 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0757 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0757 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0757 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0757 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0757 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0757 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0305 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0305 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0305 [2], \xm8051_golden_model_1.n0483 [2]);
  buf(\xm8051_golden_model_1.n0305 [3], \xm8051_golden_model_1.n0483 [3]);
  buf(\xm8051_golden_model_1.n0305 [4], \xm8051_golden_model_1.n0483 [4]);
  buf(\xm8051_golden_model_1.n0756 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0756 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0756 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0756 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0756 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0756 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0756 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0756 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0756 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0756 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0756 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0756 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0756 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0756 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0756 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0756 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0756 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0756 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0756 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0756 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0756 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0756 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0756 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0756 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0756 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0756 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0756 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0756 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0756 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0756 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0756 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0756 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0756 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0756 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0756 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0756 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0756 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0756 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0756 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0756 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0756 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0756 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0756 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0756 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0756 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0756 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0756 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0756 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0756 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0756 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0756 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0756 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0756 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0756 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0756 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0756 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0756 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0756 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0756 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0756 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0756 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0756 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0756 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0756 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0756 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0756 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0756 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0756 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0756 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0756 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0756 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0756 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0756 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0756 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0756 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0756 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0756 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0756 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0756 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0756 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0756 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0756 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0756 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0756 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0756 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0756 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0756 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0756 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0756 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0756 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0756 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0756 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0756 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0756 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0756 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0756 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0756 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0756 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0756 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0756 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0756 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0756 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0756 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0756 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0756 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0756 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0756 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0756 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0756 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0756 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0756 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0756 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0756 [112], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0756 [113], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0756 [114], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0756 [115], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0756 [116], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0756 [117], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0756 [118], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0756 [119], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0755 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0755 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0755 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0755 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0755 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0755 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0755 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0755 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0755 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0755 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0755 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0755 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0755 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0755 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0755 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0755 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0755 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0755 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0755 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0755 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0755 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0755 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0755 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0755 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0755 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0755 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0755 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0755 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0755 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0755 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0755 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0755 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0755 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0755 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0755 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0755 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0755 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0755 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0755 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0755 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0755 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0755 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0755 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0755 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0755 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0755 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0755 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0755 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0755 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0755 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0755 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0755 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0755 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0755 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0755 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0755 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0755 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0755 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0755 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0755 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0755 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0755 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0755 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0755 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0755 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0755 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0755 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0755 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0755 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0755 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0755 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0755 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0755 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0755 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0755 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0755 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0755 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0755 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0755 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0755 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0755 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0755 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0755 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0755 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0755 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0755 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0755 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0755 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0755 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0755 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0755 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0755 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0755 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0755 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0755 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0755 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0755 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0755 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0755 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0755 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0755 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0755 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0755 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0755 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0755 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0755 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0755 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0755 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0755 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0755 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0755 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0755 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0754 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0754 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0754 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0754 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0754 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0754 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0754 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0754 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0754 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0754 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0754 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0754 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0754 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0754 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0754 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0754 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0754 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0754 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0754 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0754 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0754 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0754 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0754 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0754 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0754 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0754 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0754 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0754 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0754 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0754 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0754 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0754 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0754 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0754 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0754 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0754 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0754 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0754 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0754 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0754 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0754 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0754 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0754 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0754 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0754 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0754 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0754 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0754 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0754 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0754 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0754 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0754 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0754 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0754 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0754 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0754 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0754 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0754 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0754 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0754 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0754 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0754 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0754 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0754 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0754 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0754 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0754 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0754 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0754 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0754 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0754 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0754 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0754 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0754 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0754 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0754 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0754 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0754 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0754 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0754 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0754 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0754 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0754 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0754 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0754 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0754 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0754 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0754 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0754 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0754 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0754 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0754 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0754 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0754 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0754 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0754 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0754 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0754 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0754 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0754 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0754 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0754 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0754 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0754 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0754 [104], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0754 [105], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0754 [106], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0754 [107], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0754 [108], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0754 [109], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0754 [110], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0754 [111], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0754 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0754 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0754 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0754 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0754 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0754 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0754 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0754 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0754 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0754 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0754 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0754 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0754 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0754 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0754 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0754 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0753 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0753 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0753 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0753 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0753 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0753 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0753 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0753 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0753 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0753 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0753 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0753 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0753 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0753 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0753 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0753 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0753 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0753 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0753 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0753 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0753 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0753 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0753 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0753 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0753 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0753 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0753 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0753 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0753 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0753 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0753 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0753 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0753 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0753 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0753 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0753 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0753 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0753 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0753 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0753 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0753 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0753 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0753 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0753 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0753 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0753 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0753 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0753 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0753 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0753 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0753 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0753 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0753 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0753 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0753 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0753 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0753 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0753 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0753 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0753 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0753 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0753 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0753 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0753 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0753 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0753 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0753 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0753 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0753 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0753 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0753 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0753 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0753 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0753 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0753 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0753 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0753 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0753 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0753 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0753 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0753 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0753 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0753 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0753 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0753 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0753 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0753 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0753 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0753 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0753 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0753 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0753 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0753 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0753 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0753 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0753 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0753 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0753 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0753 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0753 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0753 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0753 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0753 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0753 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0752 [0], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0752 [1], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0752 [2], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0752 [3], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0752 [4], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0752 [5], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0752 [6], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0752 [7], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0752 [8], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0752 [9], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0752 [10], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0752 [11], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0752 [12], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0752 [13], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0752 [14], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0752 [15], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0751 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0751 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0751 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0751 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0751 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0751 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0751 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0751 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0751 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0751 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0751 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0751 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0751 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0751 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0751 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0751 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0751 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0751 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0751 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0751 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0751 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0751 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0751 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0751 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0751 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0751 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0751 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0751 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0751 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0751 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0751 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0751 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0751 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0751 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0751 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0751 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0751 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0751 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0751 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0751 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0751 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0751 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0751 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0751 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0751 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0751 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0751 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0751 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0751 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0751 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0751 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0751 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0751 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0751 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0751 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0751 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0751 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0751 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0751 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0751 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0751 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0751 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0751 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0751 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0751 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0751 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0751 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0751 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0751 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0751 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0751 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0751 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0751 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0751 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0751 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0751 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0751 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0751 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0751 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0751 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0751 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0751 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0751 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0751 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0751 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0751 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0751 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0751 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0751 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0751 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0751 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0751 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0751 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0751 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0751 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0751 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0751 [96], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0751 [97], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0751 [98], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0751 [99], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0751 [100], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0751 [101], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0751 [102], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0751 [103], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0751 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0751 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0751 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0751 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0751 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0751 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0751 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0751 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0751 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0751 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0751 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0751 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0751 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0751 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0751 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0751 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0751 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0751 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0751 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0751 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0751 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0751 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0751 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0751 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0750 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0750 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0750 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0750 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0750 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0750 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0750 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0750 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0750 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0750 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0750 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0750 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0750 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0750 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0750 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0750 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0750 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0750 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0750 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0750 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0750 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0750 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0750 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0750 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0750 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0750 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0750 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0750 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0750 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0750 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0750 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0750 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0750 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0750 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0750 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0750 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0750 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0750 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0750 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0750 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0750 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0750 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0750 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0750 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0750 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0750 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0750 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0750 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0750 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0750 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0750 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0750 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0750 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0750 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0750 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0750 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0750 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0750 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0750 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0750 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0750 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0750 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0750 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0750 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0750 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0750 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0750 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0750 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0750 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0750 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0750 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0750 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0750 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0750 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0750 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0750 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0750 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0750 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0750 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0750 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0750 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0750 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0750 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0750 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0750 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0750 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0750 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0750 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0750 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0750 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0750 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0750 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0750 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0750 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0750 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0750 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0749 [0], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0749 [1], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0749 [2], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0749 [3], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0749 [4], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0749 [5], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0749 [6], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0749 [7], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0749 [8], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0749 [9], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0749 [10], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0749 [11], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0749 [12], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0749 [13], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0749 [14], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0749 [15], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0749 [16], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0749 [17], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0749 [18], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0749 [19], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0749 [20], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0749 [21], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0749 [22], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0749 [23], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0748 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0748 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0748 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0748 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0748 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0748 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0748 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0748 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0748 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0748 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0748 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0748 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0748 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0748 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0748 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0748 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0748 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0748 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0748 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0748 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0748 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0748 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0748 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0748 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0748 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0748 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0748 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0748 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0748 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0748 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0748 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0748 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0748 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0748 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0748 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0748 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0748 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0748 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0748 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0748 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0748 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0748 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0748 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0748 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0748 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0748 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0748 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0748 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0748 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0748 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0748 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0748 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0748 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0748 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0748 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0748 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0748 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0748 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0748 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0748 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0748 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0748 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0748 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0748 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0748 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0748 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0748 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0748 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0748 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0748 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0748 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0748 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0748 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0748 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0748 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0748 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0748 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0748 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0748 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0748 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0748 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0748 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0748 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0748 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0748 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0748 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0748 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0748 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0748 [88], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0748 [89], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0748 [90], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0748 [91], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0748 [92], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0748 [93], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0748 [94], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0748 [95], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0748 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0748 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0748 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0748 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0748 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0748 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0748 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0748 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0748 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0748 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0748 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0748 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0748 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0748 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0748 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0748 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0748 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0748 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0748 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0748 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0748 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0748 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0748 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0748 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0748 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0748 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0748 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0748 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0748 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0748 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0748 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0748 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0293 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0293 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0293 [2], \xm8051_golden_model_1.n0473 [2]);
  buf(\xm8051_golden_model_1.n0293 [3], \xm8051_golden_model_1.n0473 [3]);
  buf(\xm8051_golden_model_1.n0293 [4], \xm8051_golden_model_1.n0473 [4]);
  buf(\xm8051_golden_model_1.n0747 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0747 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0747 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0747 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0747 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0747 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0747 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0747 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0747 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0747 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0747 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0747 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0747 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0747 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0747 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0747 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0747 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0747 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0747 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0747 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0747 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0747 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0747 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0747 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0747 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0747 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0747 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0747 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0747 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0747 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0747 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0747 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0747 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0747 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0747 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0747 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0747 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0747 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0747 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0747 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0747 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0747 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0747 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0747 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0747 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0747 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0747 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0747 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0747 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0747 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0747 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0747 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0747 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0747 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0747 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0747 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0747 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0747 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0747 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0747 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0747 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0747 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0747 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0747 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0747 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0747 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0747 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0747 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0747 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0747 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0747 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0747 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0747 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0747 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0747 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0747 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0747 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0747 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0747 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0747 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0747 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0747 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0747 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0747 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0747 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0747 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0747 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0747 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0746 [0], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0746 [1], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0746 [2], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0746 [3], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0746 [4], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0746 [5], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0746 [6], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0746 [7], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0746 [8], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0746 [9], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0746 [10], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0746 [11], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0746 [12], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0746 [13], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0746 [14], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0746 [15], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0746 [16], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0746 [17], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0746 [18], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0746 [19], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0746 [20], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0746 [21], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0746 [22], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0746 [23], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0746 [24], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0746 [25], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0746 [26], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0746 [27], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0746 [28], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0746 [29], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0746 [30], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0746 [31], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0745 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0745 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0745 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0745 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0745 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0745 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0745 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0745 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0745 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0745 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0745 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0745 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0745 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0745 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0745 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0745 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0745 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0745 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0745 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0745 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0745 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0745 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0745 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0745 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0745 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0745 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0745 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0745 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0745 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0745 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0745 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0745 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0745 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0745 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0745 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0745 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0745 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0745 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0745 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0745 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0745 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0745 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0745 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0745 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0745 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0745 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0745 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0745 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0745 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0745 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0745 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0745 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0745 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0745 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0745 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0745 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0745 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0745 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0745 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0745 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0745 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0745 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0745 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0745 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0745 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0745 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0745 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0745 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0745 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0745 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0745 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0745 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0745 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0745 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0745 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0745 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0745 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0745 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0745 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0745 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0745 [80], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0745 [81], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0745 [82], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0745 [83], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0745 [84], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0745 [85], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0745 [86], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0745 [87], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0745 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0745 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0745 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0745 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0745 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0745 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0745 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0745 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0745 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0745 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0745 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0745 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0745 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0745 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0745 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0745 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0745 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0745 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0745 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0745 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0745 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0745 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0745 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0745 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0745 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0745 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0745 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0745 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0745 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0745 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0745 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0745 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0745 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0745 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0745 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0745 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0745 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0745 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0745 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0745 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0744 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0744 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0744 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0744 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0744 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0744 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0744 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0744 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0744 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0744 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0744 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0744 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0744 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0744 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0744 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0744 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0744 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0744 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0744 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0744 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0744 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0744 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0744 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0744 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0744 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0744 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0744 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0744 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0744 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0744 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0744 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0744 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0744 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0744 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0744 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0744 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0744 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0744 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0744 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0744 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0744 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0744 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0744 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0744 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0744 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0744 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0744 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0744 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0744 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0744 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0744 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0744 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0744 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0744 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0744 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0744 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0744 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0744 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0744 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0744 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0744 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0744 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0744 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0744 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0744 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0744 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0744 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0744 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0744 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0744 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0744 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0744 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0744 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0744 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0744 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0744 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0744 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0744 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0744 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0744 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0743 [0], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0743 [1], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0743 [2], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0743 [3], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0743 [4], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0743 [5], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0743 [6], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0743 [7], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0743 [8], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0743 [9], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0743 [10], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0743 [11], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0743 [12], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0743 [13], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0743 [14], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0743 [15], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0743 [16], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0743 [17], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0743 [18], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0743 [19], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0743 [20], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0743 [21], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0743 [22], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0743 [23], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0743 [24], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0743 [25], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0743 [26], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0743 [27], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0743 [28], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0743 [29], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0743 [30], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0743 [31], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0743 [32], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0743 [33], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0743 [34], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0743 [35], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0743 [36], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0743 [37], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0743 [38], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0743 [39], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0742 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0742 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0742 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0742 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0742 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0742 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0742 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0742 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0742 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0742 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0742 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0742 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0742 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0742 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0742 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0742 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0742 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0742 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0742 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0742 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0742 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0742 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0742 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0742 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0742 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0742 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0742 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0742 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0742 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0742 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0742 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0742 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0742 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0742 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0742 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0742 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0742 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0742 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0742 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0742 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0742 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0742 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0742 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0742 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0742 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0742 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0742 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0742 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0742 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0742 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0742 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0742 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0742 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0742 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0742 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0742 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0742 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0742 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0742 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0742 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0742 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0742 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0742 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0742 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0742 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0742 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0742 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0742 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0742 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0742 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0742 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0742 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0742 [72], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0742 [73], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0742 [74], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0742 [75], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0742 [76], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0742 [77], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0742 [78], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0742 [79], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0742 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0742 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0742 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0742 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0742 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0742 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0742 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0742 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0742 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0742 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0742 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0742 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0742 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0742 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0742 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0742 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0742 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0742 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0742 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0742 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0742 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0742 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0742 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0742 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0742 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0742 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0742 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0742 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0742 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0742 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0742 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0742 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0742 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0742 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0742 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0742 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0742 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0742 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0742 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0742 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0742 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0742 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0742 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0742 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0742 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0742 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0742 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0742 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0741 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0741 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0741 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0741 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0741 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0741 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0741 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0741 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0741 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0741 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0741 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0741 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0741 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0741 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0741 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0741 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0741 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0741 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0741 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0741 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0741 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0741 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0741 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0741 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0741 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0741 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0741 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0741 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0741 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0741 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0741 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0741 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0741 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0741 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0741 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0741 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0741 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0741 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0741 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0741 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0741 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0741 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0741 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0741 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0741 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0741 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0741 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0741 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0741 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0741 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0741 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0741 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0741 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0741 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0741 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0741 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0741 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0741 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0741 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0741 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0741 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0741 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0741 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0741 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0741 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0741 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0741 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0741 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0741 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0741 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0741 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0741 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0740 [0], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0740 [1], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0740 [2], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0740 [3], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0740 [4], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0740 [5], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0740 [6], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0740 [7], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0740 [8], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0740 [9], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0740 [10], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0740 [11], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0740 [12], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0740 [13], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0740 [14], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0740 [15], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0740 [16], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0740 [17], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0740 [18], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0740 [19], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0740 [20], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0740 [21], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0740 [22], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0740 [23], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0740 [24], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0740 [25], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0740 [26], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0740 [27], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0740 [28], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0740 [29], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0740 [30], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0740 [31], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0740 [32], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0740 [33], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0740 [34], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0740 [35], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0740 [36], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0740 [37], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0740 [38], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0740 [39], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0740 [40], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0740 [41], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0740 [42], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0740 [43], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0740 [44], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0740 [45], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0740 [46], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0740 [47], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0739 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0739 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0739 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0739 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0739 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0739 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0739 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0739 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0739 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0739 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0739 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0739 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0739 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0739 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0739 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0739 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0739 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0739 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0739 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0739 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0739 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0739 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0739 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0739 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0739 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0739 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0739 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0739 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0739 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0739 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0739 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0739 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0739 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0739 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0739 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0739 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0739 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0739 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0739 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0739 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0739 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0739 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0739 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0739 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0739 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0739 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0739 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0739 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0739 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0739 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0739 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0739 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0739 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0739 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0739 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0739 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0739 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0739 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0739 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0739 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0739 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0739 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0739 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0739 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0739 [64], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0739 [65], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0739 [66], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0739 [67], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0739 [68], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0739 [69], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0739 [70], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0739 [71], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0739 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0739 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0739 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0739 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0739 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0739 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0739 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0739 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0739 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0739 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0739 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0739 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0739 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0739 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0739 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0739 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0739 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0739 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0739 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0739 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0739 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0739 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0739 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0739 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0739 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0739 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0739 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0739 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0739 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0739 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0739 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0739 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0739 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0739 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0739 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0739 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0739 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0739 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0739 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0739 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0739 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0739 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0739 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0739 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0739 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0739 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0739 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0739 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0739 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0739 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0739 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0739 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0739 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0739 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0739 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0739 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0738 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0738 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0738 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0738 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0738 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0738 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0738 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0738 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0738 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0738 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0738 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0738 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0738 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0738 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0738 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0738 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0738 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0738 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0738 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0738 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0738 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0738 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0738 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0738 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0738 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0738 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0738 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0738 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0738 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0738 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0738 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0738 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0738 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0738 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0738 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0738 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0738 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0738 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0738 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0738 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0738 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0738 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0738 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0738 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0738 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0738 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0738 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0738 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0738 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0738 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0738 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0738 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0738 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0738 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0738 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0738 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0738 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0738 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0738 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0738 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0738 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0738 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0738 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0738 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0737 [0], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0737 [1], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0737 [2], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0737 [3], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0737 [4], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0737 [5], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0737 [6], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0737 [7], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0737 [8], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0737 [9], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0737 [10], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0737 [11], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0737 [12], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0737 [13], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0737 [14], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0737 [15], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0737 [16], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0737 [17], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0737 [18], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0737 [19], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0737 [20], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0737 [21], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0737 [22], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0737 [23], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0737 [24], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0737 [25], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0737 [26], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0737 [27], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0737 [28], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0737 [29], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0737 [30], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0737 [31], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0737 [32], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0737 [33], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0737 [34], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0737 [35], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0737 [36], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0737 [37], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0737 [38], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0737 [39], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0737 [40], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0737 [41], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0737 [42], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0737 [43], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0737 [44], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0737 [45], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0737 [46], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0737 [47], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0737 [48], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0737 [49], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0737 [50], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0737 [51], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0737 [52], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0737 [53], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0737 [54], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0737 [55], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0281 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0281 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0281 [2], \xm8051_golden_model_1.n0463 [2]);
  buf(\xm8051_golden_model_1.n0281 [3], \xm8051_golden_model_1.n0463 [3]);
  buf(\xm8051_golden_model_1.n0281 [4], \xm8051_golden_model_1.n0463 [4]);
  buf(\xm8051_golden_model_1.n0736 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0736 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0736 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0736 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0736 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0736 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0736 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0736 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0736 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0736 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0736 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0736 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0736 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0736 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0736 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0736 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0736 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0736 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0736 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0736 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0736 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0736 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0736 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0736 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0736 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0736 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0736 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0736 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0736 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0736 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0736 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0736 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0736 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0736 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0736 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0736 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0736 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0736 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0736 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0736 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0736 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0736 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0736 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0736 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0736 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0736 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0736 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0736 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0736 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0736 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0736 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0736 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0736 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0736 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0736 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0736 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0736 [56], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0736 [57], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0736 [58], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0736 [59], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0736 [60], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0736 [61], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0736 [62], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0736 [63], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0736 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0736 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0736 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0736 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0736 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0736 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0736 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0736 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0736 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0736 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0736 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0736 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0736 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0736 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0736 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0736 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0736 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0736 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0736 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0736 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0736 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0736 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0736 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0736 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0736 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0736 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0736 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0736 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0736 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0736 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0736 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0736 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0736 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0736 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0736 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0736 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0736 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0736 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0736 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0736 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0736 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0736 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0736 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0736 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0736 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0736 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0736 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0736 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0736 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0736 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0736 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0736 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0736 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0736 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0736 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0736 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0736 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0736 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0736 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0736 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0736 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0736 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0736 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0736 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0735 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0735 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0735 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0735 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0735 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0735 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0735 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0735 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0735 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0735 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0735 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0735 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0735 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0735 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0735 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0735 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0735 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0735 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0735 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0735 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0735 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0735 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0735 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0735 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0735 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0735 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0735 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0735 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0735 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0735 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0735 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0735 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0735 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0735 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0735 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0735 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0735 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0735 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0735 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0735 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0735 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0735 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0735 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0735 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0735 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0735 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0735 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0735 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0735 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0735 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0735 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0735 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0735 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0735 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0735 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0735 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0734 [0], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0734 [1], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0734 [2], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0734 [3], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0734 [4], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0734 [5], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0734 [6], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0734 [7], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0734 [8], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0734 [9], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0734 [10], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0734 [11], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0734 [12], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0734 [13], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0734 [14], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0734 [15], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0734 [16], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0734 [17], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0734 [18], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0734 [19], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0734 [20], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0734 [21], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0734 [22], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0734 [23], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0734 [24], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0734 [25], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0734 [26], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0734 [27], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0734 [28], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0734 [29], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0734 [30], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0734 [31], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0734 [32], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0734 [33], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0734 [34], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0734 [35], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0734 [36], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0734 [37], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0734 [38], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0734 [39], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0734 [40], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0734 [41], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0734 [42], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0734 [43], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0734 [44], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0734 [45], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0734 [46], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0734 [47], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0734 [48], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0734 [49], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0734 [50], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0734 [51], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0734 [52], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0734 [53], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0734 [54], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0734 [55], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0734 [56], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0734 [57], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0734 [58], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0734 [59], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0734 [60], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0734 [61], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0734 [62], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0734 [63], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0733 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0733 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0733 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0733 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0733 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0733 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0733 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0733 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0733 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0733 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0733 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0733 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0733 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0733 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0733 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0733 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0733 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0733 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0733 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0733 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0733 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0733 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0733 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0733 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0733 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0733 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0733 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0733 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0733 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0733 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0733 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0733 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0733 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0733 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0733 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0733 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0733 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0733 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0733 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0733 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0733 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0733 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0733 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0733 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0733 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0733 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0733 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0733 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0733 [48], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0733 [49], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0733 [50], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0733 [51], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0733 [52], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0733 [53], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0733 [54], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0733 [55], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0733 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0733 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0733 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0733 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0733 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0733 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0733 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0733 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0733 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0733 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0733 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0733 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0733 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0733 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0733 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0733 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0733 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0733 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0733 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0733 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0733 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0733 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0733 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0733 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0733 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0733 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0733 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0733 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0733 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0733 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0733 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0733 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0733 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0733 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0733 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0733 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0733 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0733 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0733 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0733 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0733 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0733 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0733 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0733 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0733 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0733 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0733 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0733 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0733 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0733 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0733 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0733 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0733 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0733 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0733 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0733 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0733 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0733 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0733 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0733 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0733 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0733 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0733 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0733 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0733 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0733 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0733 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0733 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0733 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0733 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0733 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0733 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0732 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0732 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0732 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0732 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0732 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0732 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0732 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0732 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0732 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0732 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0732 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0732 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0732 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0732 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0732 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0732 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0732 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0732 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0732 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0732 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0732 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0732 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0732 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0732 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0732 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0732 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0732 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0732 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0732 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0732 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0732 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0732 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0732 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0732 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0732 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0732 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0732 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0732 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0732 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0732 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0732 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0732 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0732 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0732 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0732 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0732 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0732 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0732 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0731 [0], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0731 [1], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0731 [2], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0731 [3], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0731 [4], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0731 [5], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0731 [6], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0731 [7], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0731 [8], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0731 [9], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0731 [10], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0731 [11], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0731 [12], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0731 [13], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0731 [14], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0731 [15], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0731 [16], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0731 [17], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0731 [18], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0731 [19], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0731 [20], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0731 [21], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0731 [22], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0731 [23], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0731 [24], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0731 [25], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0731 [26], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0731 [27], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0731 [28], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0731 [29], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0731 [30], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0731 [31], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0731 [32], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0731 [33], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0731 [34], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0731 [35], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0731 [36], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0731 [37], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0731 [38], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0731 [39], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0731 [40], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0731 [41], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0731 [42], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0731 [43], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0731 [44], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0731 [45], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0731 [46], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0731 [47], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0731 [48], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0731 [49], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0731 [50], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0731 [51], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0731 [52], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0731 [53], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0731 [54], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0731 [55], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0731 [56], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0731 [57], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0731 [58], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0731 [59], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0731 [60], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0731 [61], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0731 [62], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0731 [63], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0731 [64], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0731 [65], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0731 [66], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0731 [67], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0731 [68], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0731 [69], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0731 [70], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0731 [71], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0730 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0730 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0730 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0730 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0730 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0730 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0730 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0730 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0730 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0730 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0730 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0730 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0730 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0730 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0730 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0730 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0730 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0730 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0730 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0730 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0730 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0730 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0730 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0730 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0730 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0730 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0730 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0730 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0730 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0730 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0730 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0730 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0730 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0730 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0730 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0730 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0730 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0730 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0730 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0730 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0730 [40], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0730 [41], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0730 [42], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0730 [43], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0730 [44], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0730 [45], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0730 [46], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0730 [47], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0730 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0730 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0730 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0730 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0730 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0730 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0730 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0730 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0730 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0730 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0730 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0730 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0730 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0730 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0730 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0730 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0730 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0730 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0730 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0730 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0730 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0730 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0730 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0730 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0730 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0730 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0730 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0730 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0730 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0730 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0730 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0730 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0730 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0730 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0730 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0730 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0730 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0730 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0730 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0730 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0730 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0730 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0730 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0730 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0730 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0730 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0730 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0730 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0730 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0730 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0730 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0730 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0730 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0730 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0730 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0730 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0730 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0730 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0730 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0730 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0730 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0730 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0730 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0730 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0730 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0730 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0730 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0730 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0730 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0730 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0730 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0730 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0730 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0730 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0730 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0730 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0730 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0730 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0730 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0730 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0729 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0729 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0729 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0729 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0729 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0729 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0729 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0729 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0729 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0729 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0729 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0729 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0729 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0729 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0729 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0729 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0729 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0729 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0729 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0729 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0729 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0729 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0729 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0729 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0729 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0729 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0729 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0729 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0729 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0729 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0729 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0729 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0729 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0729 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0729 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0729 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0729 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0729 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0729 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0729 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0728 [0], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0728 [1], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0728 [2], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0728 [3], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0728 [4], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0728 [5], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0728 [6], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0728 [7], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0728 [8], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0728 [9], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0728 [10], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0728 [11], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0728 [12], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0728 [13], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0728 [14], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0728 [15], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0728 [16], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0728 [17], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0728 [18], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0728 [19], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0728 [20], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0728 [21], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0728 [22], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0728 [23], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0728 [24], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0728 [25], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0728 [26], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0728 [27], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0728 [28], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0728 [29], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0728 [30], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0728 [31], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0728 [32], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0728 [33], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0728 [34], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0728 [35], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0728 [36], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0728 [37], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0728 [38], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0728 [39], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0728 [40], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0728 [41], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0728 [42], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0728 [43], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0728 [44], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0728 [45], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0728 [46], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0728 [47], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0728 [48], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0728 [49], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0728 [50], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0728 [51], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0728 [52], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0728 [53], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0728 [54], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0728 [55], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0728 [56], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0728 [57], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0728 [58], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0728 [59], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0728 [60], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0728 [61], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0728 [62], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0728 [63], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0728 [64], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0728 [65], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0728 [66], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0728 [67], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0728 [68], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0728 [69], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0728 [70], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0728 [71], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0728 [72], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0728 [73], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0728 [74], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0728 [75], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0728 [76], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0728 [77], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0728 [78], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0728 [79], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0727 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0727 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0727 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0727 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0727 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0727 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0727 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0727 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0727 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0727 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0727 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0727 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0727 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0727 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0727 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0727 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0727 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0727 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0727 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0727 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0727 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0727 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0727 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0727 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0727 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0727 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0727 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0727 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0727 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0727 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0727 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0727 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0727 [32], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0727 [33], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0727 [34], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0727 [35], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0727 [36], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0727 [37], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0727 [38], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0727 [39], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0727 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0727 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0727 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0727 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0727 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0727 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0727 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0727 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0727 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0727 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0727 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0727 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0727 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0727 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0727 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0727 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0727 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0727 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0727 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0727 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0727 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0727 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0727 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0727 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0727 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0727 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0727 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0727 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0727 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0727 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0727 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0727 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0727 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0727 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0727 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0727 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0727 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0727 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0727 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0727 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0727 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0727 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0727 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0727 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0727 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0727 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0727 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0727 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0727 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0727 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0727 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0727 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0727 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0727 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0727 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0727 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0727 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0727 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0727 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0727 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0727 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0727 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0727 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0727 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0727 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0727 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0727 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0727 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0727 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0727 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0727 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0727 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0727 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0727 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0727 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0727 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0727 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0727 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0727 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0727 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0727 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0727 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0727 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0727 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0727 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0727 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0727 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0727 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0726 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0726 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0726 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0726 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0726 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0726 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0726 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0726 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0726 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0726 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0726 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0726 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0726 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0726 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0726 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0726 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0726 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0726 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0726 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0726 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0726 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0726 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0726 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0726 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0726 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0726 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0726 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0726 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0726 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0726 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0726 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0726 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0269 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0269 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0269 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n0269 [3], \xm8051_golden_model_1.n0453 [3]);
  buf(\xm8051_golden_model_1.n0269 [4], \xm8051_golden_model_1.n0453 [4]);
  buf(\xm8051_golden_model_1.n0725 [0], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0725 [1], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0725 [2], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0725 [3], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0725 [4], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0725 [5], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0725 [6], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0725 [7], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0725 [8], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0725 [9], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0725 [10], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0725 [11], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0725 [12], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0725 [13], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0725 [14], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0725 [15], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0725 [16], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0725 [17], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0725 [18], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0725 [19], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0725 [20], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0725 [21], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0725 [22], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0725 [23], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0725 [24], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0725 [25], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0725 [26], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0725 [27], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0725 [28], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0725 [29], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0725 [30], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0725 [31], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0725 [32], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0725 [33], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0725 [34], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0725 [35], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0725 [36], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0725 [37], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0725 [38], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0725 [39], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0725 [40], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0725 [41], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0725 [42], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0725 [43], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0725 [44], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0725 [45], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0725 [46], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0725 [47], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0725 [48], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0725 [49], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0725 [50], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0725 [51], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0725 [52], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0725 [53], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0725 [54], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0725 [55], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0725 [56], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0725 [57], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0725 [58], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0725 [59], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0725 [60], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0725 [61], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0725 [62], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0725 [63], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0725 [64], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0725 [65], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0725 [66], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0725 [67], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0725 [68], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0725 [69], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0725 [70], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0725 [71], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0725 [72], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0725 [73], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0725 [74], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0725 [75], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0725 [76], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0725 [77], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0725 [78], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0725 [79], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0725 [80], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0725 [81], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0725 [82], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0725 [83], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0725 [84], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0725 [85], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0725 [86], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0725 [87], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0724 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0724 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0724 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0724 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0724 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0724 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0724 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0724 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0724 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0724 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0724 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0724 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0724 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0724 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0724 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0724 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0724 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0724 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0724 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0724 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0724 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0724 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0724 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0724 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0724 [24], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0724 [25], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0724 [26], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0724 [27], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0724 [28], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0724 [29], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0724 [30], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0724 [31], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0724 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0724 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0724 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0724 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0724 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0724 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0724 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0724 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0724 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0724 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0724 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0724 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0724 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0724 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0724 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0724 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0724 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0724 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0724 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0724 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0724 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0724 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0724 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0724 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0724 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0724 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0724 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0724 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0724 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0724 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0724 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0724 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0724 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0724 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0724 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0724 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0724 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0724 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0724 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0724 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0724 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0724 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0724 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0724 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0724 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0724 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0724 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0724 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0724 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0724 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0724 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0724 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0724 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0724 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0724 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0724 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0724 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0724 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0724 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0724 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0724 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0724 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0724 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0724 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0724 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0724 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0724 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0724 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0724 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0724 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0724 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0724 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0724 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0724 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0724 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0724 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0724 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0724 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0724 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0724 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0724 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0724 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0724 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0724 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0724 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0724 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0724 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0724 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0724 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0724 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0724 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0724 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0724 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0724 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0724 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0724 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0723 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0723 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0723 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0723 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0723 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0723 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0723 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0723 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0723 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0723 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0723 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0723 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0723 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0723 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0723 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0723 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0723 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0723 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0723 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0723 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0723 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0723 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0723 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0723 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0722 [0], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0722 [1], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0722 [2], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0722 [3], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0722 [4], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0722 [5], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0722 [6], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0722 [7], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0722 [8], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0722 [9], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0722 [10], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0722 [11], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0722 [12], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0722 [13], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0722 [14], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0722 [15], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0722 [16], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0722 [17], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0722 [18], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0722 [19], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0722 [20], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0722 [21], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0722 [22], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0722 [23], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0722 [24], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0722 [25], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0722 [26], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0722 [27], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0722 [28], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0722 [29], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0722 [30], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0722 [31], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0722 [32], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0722 [33], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0722 [34], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0722 [35], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0722 [36], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0722 [37], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0722 [38], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0722 [39], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0722 [40], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0722 [41], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0722 [42], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0722 [43], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0722 [44], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0722 [45], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0722 [46], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0722 [47], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0722 [48], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0722 [49], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0722 [50], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0722 [51], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0722 [52], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0722 [53], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0722 [54], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0722 [55], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0722 [56], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0722 [57], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0722 [58], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0722 [59], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0722 [60], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0722 [61], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0722 [62], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0722 [63], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0722 [64], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0722 [65], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0722 [66], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0722 [67], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0722 [68], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0722 [69], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0722 [70], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0722 [71], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0722 [72], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0722 [73], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0722 [74], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0722 [75], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0722 [76], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0722 [77], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0722 [78], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0722 [79], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0722 [80], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0722 [81], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0722 [82], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0722 [83], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0722 [84], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0722 [85], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0722 [86], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0722 [87], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0722 [88], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0722 [89], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0722 [90], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0722 [91], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0722 [92], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0722 [93], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0722 [94], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0722 [95], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0721 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0721 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0721 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0721 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0721 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0721 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0721 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0721 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0721 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0721 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0721 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0721 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0721 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0721 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0721 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0721 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0721 [16], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0721 [17], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0721 [18], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0721 [19], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0721 [20], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0721 [21], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0721 [22], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0721 [23], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0721 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0721 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0721 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0721 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0721 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0721 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0721 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0721 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0721 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0721 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0721 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0721 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0721 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0721 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0721 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0721 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0721 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0721 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0721 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0721 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0721 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0721 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0721 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0721 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0721 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0721 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0721 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0721 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0721 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0721 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0721 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0721 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0721 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0721 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0721 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0721 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0721 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0721 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0721 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0721 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0721 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0721 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0721 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0721 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0721 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0721 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0721 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0721 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0721 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0721 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0721 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0721 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0721 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0721 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0721 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0721 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0721 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0721 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0721 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0721 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0721 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0721 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0721 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0721 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0721 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0721 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0721 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0721 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0721 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0721 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0721 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0721 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0721 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0721 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0721 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0721 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0721 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0721 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0721 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0721 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0721 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0721 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0721 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0721 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0721 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0721 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0721 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0721 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0721 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0721 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0721 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0721 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0721 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0721 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0721 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0721 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0721 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0721 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0721 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0721 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0721 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0721 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0721 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0721 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0720 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0720 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0720 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0720 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0720 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0720 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0720 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0720 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0720 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0720 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0720 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0720 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0720 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0720 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0720 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0720 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0719 [0], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0719 [1], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0719 [2], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0719 [3], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0719 [4], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0719 [5], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0719 [6], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0719 [7], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0719 [8], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0719 [9], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0719 [10], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0719 [11], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0719 [12], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0719 [13], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0719 [14], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0719 [15], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0719 [16], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0719 [17], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0719 [18], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0719 [19], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0719 [20], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0719 [21], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0719 [22], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0719 [23], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0719 [24], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0719 [25], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0719 [26], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0719 [27], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0719 [28], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0719 [29], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0719 [30], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0719 [31], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0719 [32], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0719 [33], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0719 [34], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0719 [35], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0719 [36], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0719 [37], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0719 [38], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0719 [39], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0719 [40], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0719 [41], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0719 [42], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0719 [43], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0719 [44], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0719 [45], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0719 [46], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0719 [47], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0719 [48], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0719 [49], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0719 [50], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0719 [51], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0719 [52], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0719 [53], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0719 [54], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0719 [55], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0719 [56], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0719 [57], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0719 [58], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0719 [59], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0719 [60], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0719 [61], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0719 [62], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0719 [63], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0719 [64], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0719 [65], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0719 [66], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0719 [67], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0719 [68], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0719 [69], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0719 [70], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0719 [71], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0719 [72], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0719 [73], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0719 [74], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0719 [75], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0719 [76], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0719 [77], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0719 [78], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0719 [79], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0719 [80], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0719 [81], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0719 [82], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0719 [83], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0719 [84], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0719 [85], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0719 [86], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0719 [87], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0719 [88], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0719 [89], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0719 [90], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0719 [91], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0719 [92], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0719 [93], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0719 [94], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0719 [95], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0719 [96], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0719 [97], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0719 [98], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0719 [99], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0719 [100], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0719 [101], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0719 [102], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0719 [103], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0718 [0], \xm8051_golden_model_1.n0772 [0]);
  buf(\xm8051_golden_model_1.n0718 [1], \xm8051_golden_model_1.n0772 [1]);
  buf(\xm8051_golden_model_1.n0718 [2], \xm8051_golden_model_1.n0772 [2]);
  buf(\xm8051_golden_model_1.n0718 [3], \xm8051_golden_model_1.n0772 [3]);
  buf(\xm8051_golden_model_1.n0718 [4], \xm8051_golden_model_1.n0772 [4]);
  buf(\xm8051_golden_model_1.n0718 [5], \xm8051_golden_model_1.n0772 [5]);
  buf(\xm8051_golden_model_1.n0718 [6], \xm8051_golden_model_1.n0772 [6]);
  buf(\xm8051_golden_model_1.n0718 [7], \xm8051_golden_model_1.n0772 [7]);
  buf(\xm8051_golden_model_1.n0718 [8], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0718 [9], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0718 [10], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0718 [11], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0718 [12], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0718 [13], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0718 [14], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0718 [15], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0718 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0718 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0718 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0718 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0718 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0718 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0718 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0718 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0718 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0718 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0718 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0718 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0718 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0718 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0718 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0718 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0718 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0718 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0718 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0718 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0718 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0718 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0718 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0718 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0718 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0718 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0718 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0718 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0718 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0718 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0718 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0718 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0718 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0718 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0718 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0718 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0718 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0718 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0718 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0718 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0718 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0718 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0718 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0718 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0718 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0718 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0718 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0718 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0718 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0718 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0718 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0718 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0718 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0718 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0718 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0718 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0718 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0718 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0718 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0718 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0718 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0718 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0718 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0718 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0718 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0718 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0718 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0718 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0718 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0718 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0718 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0718 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0718 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0718 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0718 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0718 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0718 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0718 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0718 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0718 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0718 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0718 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0718 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0718 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0718 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0718 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0718 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0718 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0718 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0718 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0718 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0718 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0718 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0718 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0718 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0718 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0718 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0718 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0718 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0718 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0718 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0718 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0718 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0718 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0718 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0718 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0718 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0718 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0718 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0718 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0718 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0718 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0717 [0], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0717 [1], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0717 [2], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0717 [3], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0717 [4], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0717 [5], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0717 [6], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0717 [7], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0717 [8], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0717 [9], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0717 [10], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0717 [11], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0717 [12], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0717 [13], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0717 [14], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0717 [15], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0717 [16], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0717 [17], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0717 [18], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0717 [19], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0717 [20], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0717 [21], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0717 [22], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0717 [23], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0717 [24], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0717 [25], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0717 [26], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0717 [27], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0717 [28], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0717 [29], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0717 [30], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0717 [31], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0717 [32], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0717 [33], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0717 [34], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0717 [35], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0717 [36], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0717 [37], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0717 [38], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0717 [39], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0717 [40], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0717 [41], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0717 [42], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0717 [43], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0717 [44], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0717 [45], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0717 [46], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0717 [47], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0717 [48], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0717 [49], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0717 [50], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0717 [51], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0717 [52], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0717 [53], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0717 [54], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0717 [55], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0717 [56], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0717 [57], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0717 [58], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0717 [59], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0717 [60], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0717 [61], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0717 [62], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0717 [63], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0717 [64], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0717 [65], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0717 [66], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0717 [67], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0717 [68], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0717 [69], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0717 [70], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0717 [71], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0717 [72], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0717 [73], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0717 [74], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0717 [75], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0717 [76], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0717 [77], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0717 [78], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0717 [79], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0717 [80], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0717 [81], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0717 [82], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0717 [83], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0717 [84], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0717 [85], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0717 [86], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0717 [87], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0717 [88], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0717 [89], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0717 [90], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0717 [91], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0717 [92], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0717 [93], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0717 [94], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0717 [95], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0717 [96], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0717 [97], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0717 [98], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0717 [99], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0717 [100], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0717 [101], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0717 [102], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0717 [103], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0717 [104], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0717 [105], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0717 [106], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0717 [107], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0717 [108], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0717 [109], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0717 [110], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0717 [111], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0716 [0], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0716 [1], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0716 [2], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0716 [3], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0716 [4], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0716 [5], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0716 [6], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0716 [7], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0716 [8], \xm8051_golden_model_1.n0771 [8]);
  buf(\xm8051_golden_model_1.n0716 [9], \xm8051_golden_model_1.n0771 [9]);
  buf(\xm8051_golden_model_1.n0716 [10], \xm8051_golden_model_1.n0771 [10]);
  buf(\xm8051_golden_model_1.n0716 [11], \xm8051_golden_model_1.n0771 [11]);
  buf(\xm8051_golden_model_1.n0716 [12], \xm8051_golden_model_1.n0771 [12]);
  buf(\xm8051_golden_model_1.n0716 [13], \xm8051_golden_model_1.n0771 [13]);
  buf(\xm8051_golden_model_1.n0716 [14], \xm8051_golden_model_1.n0771 [14]);
  buf(\xm8051_golden_model_1.n0716 [15], \xm8051_golden_model_1.n0771 [15]);
  buf(\xm8051_golden_model_1.n0716 [16], \xm8051_golden_model_1.n0770 [16]);
  buf(\xm8051_golden_model_1.n0716 [17], \xm8051_golden_model_1.n0770 [17]);
  buf(\xm8051_golden_model_1.n0716 [18], \xm8051_golden_model_1.n0770 [18]);
  buf(\xm8051_golden_model_1.n0716 [19], \xm8051_golden_model_1.n0770 [19]);
  buf(\xm8051_golden_model_1.n0716 [20], \xm8051_golden_model_1.n0770 [20]);
  buf(\xm8051_golden_model_1.n0716 [21], \xm8051_golden_model_1.n0770 [21]);
  buf(\xm8051_golden_model_1.n0716 [22], \xm8051_golden_model_1.n0770 [22]);
  buf(\xm8051_golden_model_1.n0716 [23], \xm8051_golden_model_1.n0770 [23]);
  buf(\xm8051_golden_model_1.n0716 [24], \xm8051_golden_model_1.n0769 [24]);
  buf(\xm8051_golden_model_1.n0716 [25], \xm8051_golden_model_1.n0769 [25]);
  buf(\xm8051_golden_model_1.n0716 [26], \xm8051_golden_model_1.n0769 [26]);
  buf(\xm8051_golden_model_1.n0716 [27], \xm8051_golden_model_1.n0769 [27]);
  buf(\xm8051_golden_model_1.n0716 [28], \xm8051_golden_model_1.n0769 [28]);
  buf(\xm8051_golden_model_1.n0716 [29], \xm8051_golden_model_1.n0769 [29]);
  buf(\xm8051_golden_model_1.n0716 [30], \xm8051_golden_model_1.n0769 [30]);
  buf(\xm8051_golden_model_1.n0716 [31], \xm8051_golden_model_1.n0769 [31]);
  buf(\xm8051_golden_model_1.n0716 [32], \xm8051_golden_model_1.n0768 [32]);
  buf(\xm8051_golden_model_1.n0716 [33], \xm8051_golden_model_1.n0768 [33]);
  buf(\xm8051_golden_model_1.n0716 [34], \xm8051_golden_model_1.n0768 [34]);
  buf(\xm8051_golden_model_1.n0716 [35], \xm8051_golden_model_1.n0768 [35]);
  buf(\xm8051_golden_model_1.n0716 [36], \xm8051_golden_model_1.n0768 [36]);
  buf(\xm8051_golden_model_1.n0716 [37], \xm8051_golden_model_1.n0768 [37]);
  buf(\xm8051_golden_model_1.n0716 [38], \xm8051_golden_model_1.n0768 [38]);
  buf(\xm8051_golden_model_1.n0716 [39], \xm8051_golden_model_1.n0768 [39]);
  buf(\xm8051_golden_model_1.n0716 [40], \xm8051_golden_model_1.n0767 [40]);
  buf(\xm8051_golden_model_1.n0716 [41], \xm8051_golden_model_1.n0767 [41]);
  buf(\xm8051_golden_model_1.n0716 [42], \xm8051_golden_model_1.n0767 [42]);
  buf(\xm8051_golden_model_1.n0716 [43], \xm8051_golden_model_1.n0767 [43]);
  buf(\xm8051_golden_model_1.n0716 [44], \xm8051_golden_model_1.n0767 [44]);
  buf(\xm8051_golden_model_1.n0716 [45], \xm8051_golden_model_1.n0767 [45]);
  buf(\xm8051_golden_model_1.n0716 [46], \xm8051_golden_model_1.n0767 [46]);
  buf(\xm8051_golden_model_1.n0716 [47], \xm8051_golden_model_1.n0767 [47]);
  buf(\xm8051_golden_model_1.n0716 [48], \xm8051_golden_model_1.n0766 [48]);
  buf(\xm8051_golden_model_1.n0716 [49], \xm8051_golden_model_1.n0766 [49]);
  buf(\xm8051_golden_model_1.n0716 [50], \xm8051_golden_model_1.n0766 [50]);
  buf(\xm8051_golden_model_1.n0716 [51], \xm8051_golden_model_1.n0766 [51]);
  buf(\xm8051_golden_model_1.n0716 [52], \xm8051_golden_model_1.n0766 [52]);
  buf(\xm8051_golden_model_1.n0716 [53], \xm8051_golden_model_1.n0766 [53]);
  buf(\xm8051_golden_model_1.n0716 [54], \xm8051_golden_model_1.n0766 [54]);
  buf(\xm8051_golden_model_1.n0716 [55], \xm8051_golden_model_1.n0766 [55]);
  buf(\xm8051_golden_model_1.n0716 [56], \xm8051_golden_model_1.n0765 [56]);
  buf(\xm8051_golden_model_1.n0716 [57], \xm8051_golden_model_1.n0765 [57]);
  buf(\xm8051_golden_model_1.n0716 [58], \xm8051_golden_model_1.n0765 [58]);
  buf(\xm8051_golden_model_1.n0716 [59], \xm8051_golden_model_1.n0765 [59]);
  buf(\xm8051_golden_model_1.n0716 [60], \xm8051_golden_model_1.n0765 [60]);
  buf(\xm8051_golden_model_1.n0716 [61], \xm8051_golden_model_1.n0765 [61]);
  buf(\xm8051_golden_model_1.n0716 [62], \xm8051_golden_model_1.n0765 [62]);
  buf(\xm8051_golden_model_1.n0716 [63], \xm8051_golden_model_1.n0765 [63]);
  buf(\xm8051_golden_model_1.n0716 [64], \xm8051_golden_model_1.n0764 [64]);
  buf(\xm8051_golden_model_1.n0716 [65], \xm8051_golden_model_1.n0764 [65]);
  buf(\xm8051_golden_model_1.n0716 [66], \xm8051_golden_model_1.n0764 [66]);
  buf(\xm8051_golden_model_1.n0716 [67], \xm8051_golden_model_1.n0764 [67]);
  buf(\xm8051_golden_model_1.n0716 [68], \xm8051_golden_model_1.n0764 [68]);
  buf(\xm8051_golden_model_1.n0716 [69], \xm8051_golden_model_1.n0764 [69]);
  buf(\xm8051_golden_model_1.n0716 [70], \xm8051_golden_model_1.n0764 [70]);
  buf(\xm8051_golden_model_1.n0716 [71], \xm8051_golden_model_1.n0764 [71]);
  buf(\xm8051_golden_model_1.n0716 [72], \xm8051_golden_model_1.n0763 [72]);
  buf(\xm8051_golden_model_1.n0716 [73], \xm8051_golden_model_1.n0763 [73]);
  buf(\xm8051_golden_model_1.n0716 [74], \xm8051_golden_model_1.n0763 [74]);
  buf(\xm8051_golden_model_1.n0716 [75], \xm8051_golden_model_1.n0763 [75]);
  buf(\xm8051_golden_model_1.n0716 [76], \xm8051_golden_model_1.n0763 [76]);
  buf(\xm8051_golden_model_1.n0716 [77], \xm8051_golden_model_1.n0763 [77]);
  buf(\xm8051_golden_model_1.n0716 [78], \xm8051_golden_model_1.n0763 [78]);
  buf(\xm8051_golden_model_1.n0716 [79], \xm8051_golden_model_1.n0763 [79]);
  buf(\xm8051_golden_model_1.n0716 [80], \xm8051_golden_model_1.n0762 [80]);
  buf(\xm8051_golden_model_1.n0716 [81], \xm8051_golden_model_1.n0762 [81]);
  buf(\xm8051_golden_model_1.n0716 [82], \xm8051_golden_model_1.n0762 [82]);
  buf(\xm8051_golden_model_1.n0716 [83], \xm8051_golden_model_1.n0762 [83]);
  buf(\xm8051_golden_model_1.n0716 [84], \xm8051_golden_model_1.n0762 [84]);
  buf(\xm8051_golden_model_1.n0716 [85], \xm8051_golden_model_1.n0762 [85]);
  buf(\xm8051_golden_model_1.n0716 [86], \xm8051_golden_model_1.n0762 [86]);
  buf(\xm8051_golden_model_1.n0716 [87], \xm8051_golden_model_1.n0762 [87]);
  buf(\xm8051_golden_model_1.n0716 [88], \xm8051_golden_model_1.n0761 [88]);
  buf(\xm8051_golden_model_1.n0716 [89], \xm8051_golden_model_1.n0761 [89]);
  buf(\xm8051_golden_model_1.n0716 [90], \xm8051_golden_model_1.n0761 [90]);
  buf(\xm8051_golden_model_1.n0716 [91], \xm8051_golden_model_1.n0761 [91]);
  buf(\xm8051_golden_model_1.n0716 [92], \xm8051_golden_model_1.n0761 [92]);
  buf(\xm8051_golden_model_1.n0716 [93], \xm8051_golden_model_1.n0761 [93]);
  buf(\xm8051_golden_model_1.n0716 [94], \xm8051_golden_model_1.n0761 [94]);
  buf(\xm8051_golden_model_1.n0716 [95], \xm8051_golden_model_1.n0761 [95]);
  buf(\xm8051_golden_model_1.n0716 [96], \xm8051_golden_model_1.n0760 [96]);
  buf(\xm8051_golden_model_1.n0716 [97], \xm8051_golden_model_1.n0760 [97]);
  buf(\xm8051_golden_model_1.n0716 [98], \xm8051_golden_model_1.n0760 [98]);
  buf(\xm8051_golden_model_1.n0716 [99], \xm8051_golden_model_1.n0760 [99]);
  buf(\xm8051_golden_model_1.n0716 [100], \xm8051_golden_model_1.n0760 [100]);
  buf(\xm8051_golden_model_1.n0716 [101], \xm8051_golden_model_1.n0760 [101]);
  buf(\xm8051_golden_model_1.n0716 [102], \xm8051_golden_model_1.n0760 [102]);
  buf(\xm8051_golden_model_1.n0716 [103], \xm8051_golden_model_1.n0760 [103]);
  buf(\xm8051_golden_model_1.n0716 [104], \xm8051_golden_model_1.n0759 [104]);
  buf(\xm8051_golden_model_1.n0716 [105], \xm8051_golden_model_1.n0759 [105]);
  buf(\xm8051_golden_model_1.n0716 [106], \xm8051_golden_model_1.n0759 [106]);
  buf(\xm8051_golden_model_1.n0716 [107], \xm8051_golden_model_1.n0759 [107]);
  buf(\xm8051_golden_model_1.n0716 [108], \xm8051_golden_model_1.n0759 [108]);
  buf(\xm8051_golden_model_1.n0716 [109], \xm8051_golden_model_1.n0759 [109]);
  buf(\xm8051_golden_model_1.n0716 [110], \xm8051_golden_model_1.n0759 [110]);
  buf(\xm8051_golden_model_1.n0716 [111], \xm8051_golden_model_1.n0759 [111]);
  buf(\xm8051_golden_model_1.n0716 [112], \xm8051_golden_model_1.n0758 [112]);
  buf(\xm8051_golden_model_1.n0716 [113], \xm8051_golden_model_1.n0758 [113]);
  buf(\xm8051_golden_model_1.n0716 [114], \xm8051_golden_model_1.n0758 [114]);
  buf(\xm8051_golden_model_1.n0716 [115], \xm8051_golden_model_1.n0758 [115]);
  buf(\xm8051_golden_model_1.n0716 [116], \xm8051_golden_model_1.n0758 [116]);
  buf(\xm8051_golden_model_1.n0716 [117], \xm8051_golden_model_1.n0758 [117]);
  buf(\xm8051_golden_model_1.n0716 [118], \xm8051_golden_model_1.n0758 [118]);
  buf(\xm8051_golden_model_1.n0716 [119], \xm8051_golden_model_1.n0758 [119]);
  buf(\xm8051_golden_model_1.n0716 [120], \xm8051_golden_model_1.n0756 [120]);
  buf(\xm8051_golden_model_1.n0716 [121], \xm8051_golden_model_1.n0756 [121]);
  buf(\xm8051_golden_model_1.n0716 [122], \xm8051_golden_model_1.n0756 [122]);
  buf(\xm8051_golden_model_1.n0716 [123], \xm8051_golden_model_1.n0756 [123]);
  buf(\xm8051_golden_model_1.n0716 [124], \xm8051_golden_model_1.n0756 [124]);
  buf(\xm8051_golden_model_1.n0716 [125], \xm8051_golden_model_1.n0756 [125]);
  buf(\xm8051_golden_model_1.n0716 [126], \xm8051_golden_model_1.n0756 [126]);
  buf(\xm8051_golden_model_1.n0716 [127], \xm8051_golden_model_1.n0756 [127]);
  buf(\xm8051_golden_model_1.n0257 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0257 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0257 [2], \xm8051_golden_model_1.n0483 [2]);
  buf(\xm8051_golden_model_1.n0257 [3], \xm8051_golden_model_1.n0443 [3]);
  buf(\xm8051_golden_model_1.n0257 [4], \xm8051_golden_model_1.n0443 [4]);
  buf(\xm8051_golden_model_1.n1275 [0], input_sha_func_36[0]);
  buf(\xm8051_golden_model_1.n1275 [1], input_sha_func_36[1]);
  buf(\xm8051_golden_model_1.n1275 [2], input_sha_func_36[2]);
  buf(\xm8051_golden_model_1.n1275 [3], input_sha_func_36[3]);
  buf(\xm8051_golden_model_1.n1275 [4], input_sha_func_36[4]);
  buf(\xm8051_golden_model_1.n1275 [5], input_sha_func_36[5]);
  buf(\xm8051_golden_model_1.n1275 [6], input_sha_func_36[6]);
  buf(\xm8051_golden_model_1.n1275 [7], input_sha_func_36[7]);
  buf(\xm8051_golden_model_1.n1275 [8], input_sha_func_36[8]);
  buf(\xm8051_golden_model_1.n1275 [9], input_sha_func_36[9]);
  buf(\xm8051_golden_model_1.n1275 [10], input_sha_func_36[10]);
  buf(\xm8051_golden_model_1.n1275 [11], input_sha_func_36[11]);
  buf(\xm8051_golden_model_1.n1275 [12], input_sha_func_36[12]);
  buf(\xm8051_golden_model_1.n1275 [13], input_sha_func_36[13]);
  buf(\xm8051_golden_model_1.n1275 [14], input_sha_func_36[14]);
  buf(\xm8051_golden_model_1.n1275 [15], input_sha_func_36[15]);
  buf(\xm8051_golden_model_1.n1275 [16], input_sha_func_36[16]);
  buf(\xm8051_golden_model_1.n1275 [17], input_sha_func_36[17]);
  buf(\xm8051_golden_model_1.n1275 [18], input_sha_func_36[18]);
  buf(\xm8051_golden_model_1.n1275 [19], input_sha_func_36[19]);
  buf(\xm8051_golden_model_1.n1275 [20], input_sha_func_36[20]);
  buf(\xm8051_golden_model_1.n1275 [21], input_sha_func_36[21]);
  buf(\xm8051_golden_model_1.n1275 [22], input_sha_func_36[22]);
  buf(\xm8051_golden_model_1.n1275 [23], input_sha_func_36[23]);
  buf(\xm8051_golden_model_1.n1275 [24], input_sha_func_36[24]);
  buf(\xm8051_golden_model_1.n1275 [25], input_sha_func_36[25]);
  buf(\xm8051_golden_model_1.n1275 [26], input_sha_func_36[26]);
  buf(\xm8051_golden_model_1.n1275 [27], input_sha_func_36[27]);
  buf(\xm8051_golden_model_1.n1275 [28], input_sha_func_36[28]);
  buf(\xm8051_golden_model_1.n1275 [29], input_sha_func_36[29]);
  buf(\xm8051_golden_model_1.n1275 [30], input_sha_func_36[30]);
  buf(\xm8051_golden_model_1.n1275 [31], input_sha_func_36[31]);
  buf(\xm8051_golden_model_1.n1275 [32], input_sha_func_35[0]);
  buf(\xm8051_golden_model_1.n1275 [33], input_sha_func_35[1]);
  buf(\xm8051_golden_model_1.n1275 [34], input_sha_func_35[2]);
  buf(\xm8051_golden_model_1.n1275 [35], input_sha_func_35[3]);
  buf(\xm8051_golden_model_1.n1275 [36], input_sha_func_35[4]);
  buf(\xm8051_golden_model_1.n1275 [37], input_sha_func_35[5]);
  buf(\xm8051_golden_model_1.n1275 [38], input_sha_func_35[6]);
  buf(\xm8051_golden_model_1.n1275 [39], input_sha_func_35[7]);
  buf(\xm8051_golden_model_1.n1275 [40], input_sha_func_35[8]);
  buf(\xm8051_golden_model_1.n1275 [41], input_sha_func_35[9]);
  buf(\xm8051_golden_model_1.n1275 [42], input_sha_func_35[10]);
  buf(\xm8051_golden_model_1.n1275 [43], input_sha_func_35[11]);
  buf(\xm8051_golden_model_1.n1275 [44], input_sha_func_35[12]);
  buf(\xm8051_golden_model_1.n1275 [45], input_sha_func_35[13]);
  buf(\xm8051_golden_model_1.n1275 [46], input_sha_func_35[14]);
  buf(\xm8051_golden_model_1.n1275 [47], input_sha_func_35[15]);
  buf(\xm8051_golden_model_1.n1275 [48], input_sha_func_35[16]);
  buf(\xm8051_golden_model_1.n1275 [49], input_sha_func_35[17]);
  buf(\xm8051_golden_model_1.n1275 [50], input_sha_func_35[18]);
  buf(\xm8051_golden_model_1.n1275 [51], input_sha_func_35[19]);
  buf(\xm8051_golden_model_1.n1275 [52], input_sha_func_35[20]);
  buf(\xm8051_golden_model_1.n1275 [53], input_sha_func_35[21]);
  buf(\xm8051_golden_model_1.n1275 [54], input_sha_func_35[22]);
  buf(\xm8051_golden_model_1.n1275 [55], input_sha_func_35[23]);
  buf(\xm8051_golden_model_1.n1275 [56], input_sha_func_35[24]);
  buf(\xm8051_golden_model_1.n1275 [57], input_sha_func_35[25]);
  buf(\xm8051_golden_model_1.n1275 [58], input_sha_func_35[26]);
  buf(\xm8051_golden_model_1.n1275 [59], input_sha_func_35[27]);
  buf(\xm8051_golden_model_1.n1275 [60], input_sha_func_35[28]);
  buf(\xm8051_golden_model_1.n1275 [61], input_sha_func_35[29]);
  buf(\xm8051_golden_model_1.n1275 [62], input_sha_func_35[30]);
  buf(\xm8051_golden_model_1.n1275 [63], input_sha_func_35[31]);
  buf(\xm8051_golden_model_1.n1275 [64], input_sha_func_35[32]);
  buf(\xm8051_golden_model_1.n1275 [65], input_sha_func_35[33]);
  buf(\xm8051_golden_model_1.n1275 [66], input_sha_func_35[34]);
  buf(\xm8051_golden_model_1.n1275 [67], input_sha_func_35[35]);
  buf(\xm8051_golden_model_1.n1275 [68], input_sha_func_35[36]);
  buf(\xm8051_golden_model_1.n1275 [69], input_sha_func_35[37]);
  buf(\xm8051_golden_model_1.n1275 [70], input_sha_func_35[38]);
  buf(\xm8051_golden_model_1.n1275 [71], input_sha_func_35[39]);
  buf(\xm8051_golden_model_1.n1275 [72], input_sha_func_35[40]);
  buf(\xm8051_golden_model_1.n1275 [73], input_sha_func_35[41]);
  buf(\xm8051_golden_model_1.n1275 [74], input_sha_func_35[42]);
  buf(\xm8051_golden_model_1.n1275 [75], input_sha_func_35[43]);
  buf(\xm8051_golden_model_1.n1275 [76], input_sha_func_35[44]);
  buf(\xm8051_golden_model_1.n1275 [77], input_sha_func_35[45]);
  buf(\xm8051_golden_model_1.n1275 [78], input_sha_func_35[46]);
  buf(\xm8051_golden_model_1.n1275 [79], input_sha_func_35[47]);
  buf(\xm8051_golden_model_1.n1275 [80], input_sha_func_35[48]);
  buf(\xm8051_golden_model_1.n1275 [81], input_sha_func_35[49]);
  buf(\xm8051_golden_model_1.n1275 [82], input_sha_func_35[50]);
  buf(\xm8051_golden_model_1.n1275 [83], input_sha_func_35[51]);
  buf(\xm8051_golden_model_1.n1275 [84], input_sha_func_35[52]);
  buf(\xm8051_golden_model_1.n1275 [85], input_sha_func_35[53]);
  buf(\xm8051_golden_model_1.n1275 [86], input_sha_func_35[54]);
  buf(\xm8051_golden_model_1.n1275 [87], input_sha_func_35[55]);
  buf(\xm8051_golden_model_1.n1275 [88], input_sha_func_35[56]);
  buf(\xm8051_golden_model_1.n1275 [89], input_sha_func_35[57]);
  buf(\xm8051_golden_model_1.n1275 [90], input_sha_func_35[58]);
  buf(\xm8051_golden_model_1.n1275 [91], input_sha_func_35[59]);
  buf(\xm8051_golden_model_1.n1275 [92], input_sha_func_35[60]);
  buf(\xm8051_golden_model_1.n1275 [93], input_sha_func_35[61]);
  buf(\xm8051_golden_model_1.n1275 [94], input_sha_func_35[62]);
  buf(\xm8051_golden_model_1.n1275 [95], input_sha_func_35[63]);
  buf(\xm8051_golden_model_1.n1275 [96], input_sha_func_34[0]);
  buf(\xm8051_golden_model_1.n1275 [97], input_sha_func_34[1]);
  buf(\xm8051_golden_model_1.n1275 [98], input_sha_func_34[2]);
  buf(\xm8051_golden_model_1.n1275 [99], input_sha_func_34[3]);
  buf(\xm8051_golden_model_1.n1275 [100], input_sha_func_34[4]);
  buf(\xm8051_golden_model_1.n1275 [101], input_sha_func_34[5]);
  buf(\xm8051_golden_model_1.n1275 [102], input_sha_func_34[6]);
  buf(\xm8051_golden_model_1.n1275 [103], input_sha_func_34[7]);
  buf(\xm8051_golden_model_1.n1275 [104], input_sha_func_34[8]);
  buf(\xm8051_golden_model_1.n1275 [105], input_sha_func_34[9]);
  buf(\xm8051_golden_model_1.n1275 [106], input_sha_func_34[10]);
  buf(\xm8051_golden_model_1.n1275 [107], input_sha_func_34[11]);
  buf(\xm8051_golden_model_1.n1275 [108], input_sha_func_34[12]);
  buf(\xm8051_golden_model_1.n1275 [109], input_sha_func_34[13]);
  buf(\xm8051_golden_model_1.n1275 [110], input_sha_func_34[14]);
  buf(\xm8051_golden_model_1.n1275 [111], input_sha_func_34[15]);
  buf(\xm8051_golden_model_1.n1275 [112], input_sha_func_34[16]);
  buf(\xm8051_golden_model_1.n1275 [113], input_sha_func_34[17]);
  buf(\xm8051_golden_model_1.n1275 [114], input_sha_func_34[18]);
  buf(\xm8051_golden_model_1.n1275 [115], input_sha_func_34[19]);
  buf(\xm8051_golden_model_1.n1275 [116], input_sha_func_34[20]);
  buf(\xm8051_golden_model_1.n1275 [117], input_sha_func_34[21]);
  buf(\xm8051_golden_model_1.n1275 [118], input_sha_func_34[22]);
  buf(\xm8051_golden_model_1.n1275 [119], input_sha_func_34[23]);
  buf(\xm8051_golden_model_1.n1275 [120], input_sha_func_34[24]);
  buf(\xm8051_golden_model_1.n1275 [121], input_sha_func_34[25]);
  buf(\xm8051_golden_model_1.n1275 [122], input_sha_func_34[26]);
  buf(\xm8051_golden_model_1.n1275 [123], input_sha_func_34[27]);
  buf(\xm8051_golden_model_1.n1275 [124], input_sha_func_34[28]);
  buf(\xm8051_golden_model_1.n1275 [125], input_sha_func_34[29]);
  buf(\xm8051_golden_model_1.n1275 [126], input_sha_func_34[30]);
  buf(\xm8051_golden_model_1.n1275 [127], input_sha_func_34[31]);
  buf(\xm8051_golden_model_1.n1275 [128], input_sha_func_34[32]);
  buf(\xm8051_golden_model_1.n1275 [129], input_sha_func_34[33]);
  buf(\xm8051_golden_model_1.n1275 [130], input_sha_func_34[34]);
  buf(\xm8051_golden_model_1.n1275 [131], input_sha_func_34[35]);
  buf(\xm8051_golden_model_1.n1275 [132], input_sha_func_34[36]);
  buf(\xm8051_golden_model_1.n1275 [133], input_sha_func_34[37]);
  buf(\xm8051_golden_model_1.n1275 [134], input_sha_func_34[38]);
  buf(\xm8051_golden_model_1.n1275 [135], input_sha_func_34[39]);
  buf(\xm8051_golden_model_1.n1275 [136], input_sha_func_34[40]);
  buf(\xm8051_golden_model_1.n1275 [137], input_sha_func_34[41]);
  buf(\xm8051_golden_model_1.n1275 [138], input_sha_func_34[42]);
  buf(\xm8051_golden_model_1.n1275 [139], input_sha_func_34[43]);
  buf(\xm8051_golden_model_1.n1275 [140], input_sha_func_34[44]);
  buf(\xm8051_golden_model_1.n1275 [141], input_sha_func_34[45]);
  buf(\xm8051_golden_model_1.n1275 [142], input_sha_func_34[46]);
  buf(\xm8051_golden_model_1.n1275 [143], input_sha_func_34[47]);
  buf(\xm8051_golden_model_1.n1275 [144], input_sha_func_34[48]);
  buf(\xm8051_golden_model_1.n1275 [145], input_sha_func_34[49]);
  buf(\xm8051_golden_model_1.n1275 [146], input_sha_func_34[50]);
  buf(\xm8051_golden_model_1.n1275 [147], input_sha_func_34[51]);
  buf(\xm8051_golden_model_1.n1275 [148], input_sha_func_34[52]);
  buf(\xm8051_golden_model_1.n1275 [149], input_sha_func_34[53]);
  buf(\xm8051_golden_model_1.n1275 [150], input_sha_func_34[54]);
  buf(\xm8051_golden_model_1.n1275 [151], input_sha_func_34[55]);
  buf(\xm8051_golden_model_1.n1275 [152], input_sha_func_34[56]);
  buf(\xm8051_golden_model_1.n1275 [153], input_sha_func_34[57]);
  buf(\xm8051_golden_model_1.n1275 [154], input_sha_func_34[58]);
  buf(\xm8051_golden_model_1.n1275 [155], input_sha_func_34[59]);
  buf(\xm8051_golden_model_1.n1275 [156], input_sha_func_34[60]);
  buf(\xm8051_golden_model_1.n1275 [157], input_sha_func_34[61]);
  buf(\xm8051_golden_model_1.n1275 [158], input_sha_func_34[62]);
  buf(\xm8051_golden_model_1.n1275 [159], input_sha_func_34[63]);
  buf(\xm8051_golden_model_1.n0711 [0], aes_addr_gm[0]);
  buf(\xm8051_golden_model_1.n0711 [1], aes_addr_gm[1]);
  buf(\xm8051_golden_model_1.n0711 [2], aes_addr_gm[2]);
  buf(\xm8051_golden_model_1.n0711 [3], aes_addr_gm[3]);
  buf(\xm8051_golden_model_1.n0711 [4], aes_addr_gm[4]);
  buf(\xm8051_golden_model_1.n0711 [5], aes_addr_gm[5]);
  buf(\xm8051_golden_model_1.n0711 [6], aes_addr_gm[6]);
  buf(\xm8051_golden_model_1.n0711 [7], aes_addr_gm[7]);
  buf(\xm8051_golden_model_1.n0711 [8], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0711 [9], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0711 [10], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0711 [11], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0711 [12], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0711 [13], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0711 [14], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0711 [15], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0710 [0], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0710 [1], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0710 [2], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0710 [3], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0710 [4], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0710 [5], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0710 [6], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0710 [7], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0710 [8], aes_addr_gm[8]);
  buf(\xm8051_golden_model_1.n0710 [9], aes_addr_gm[9]);
  buf(\xm8051_golden_model_1.n0710 [10], aes_addr_gm[10]);
  buf(\xm8051_golden_model_1.n0710 [11], aes_addr_gm[11]);
  buf(\xm8051_golden_model_1.n0710 [12], aes_addr_gm[12]);
  buf(\xm8051_golden_model_1.n0710 [13], aes_addr_gm[13]);
  buf(\xm8051_golden_model_1.n0710 [14], aes_addr_gm[14]);
  buf(\xm8051_golden_model_1.n0710 [15], aes_addr_gm[15]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.data_in [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.data_in [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.data_in [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.data_in [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.data_in [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.data_in [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.data_in [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.data_in [7], proc_data_in[7]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.addr [0], proc_addr[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.addr [1], proc_addr[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.addr [2], proc_addr[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.addr [3], proc_addr[3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.rst , rst);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_ctr_i.clk , clk);
  buf(\xm8051_golden_model_1.n1271 [0], input_sha_func_33[0]);
  buf(\xm8051_golden_model_1.n1271 [1], input_sha_func_33[1]);
  buf(\xm8051_golden_model_1.n1271 [2], input_sha_func_33[2]);
  buf(\xm8051_golden_model_1.n1271 [3], input_sha_func_33[3]);
  buf(\xm8051_golden_model_1.n1271 [4], input_sha_func_33[4]);
  buf(\xm8051_golden_model_1.n1271 [5], input_sha_func_33[5]);
  buf(\xm8051_golden_model_1.n1271 [6], input_sha_func_33[6]);
  buf(\xm8051_golden_model_1.n1271 [7], input_sha_func_33[7]);
  buf(\xm8051_golden_model_1.n1271 [8], input_sha_func_33[8]);
  buf(\xm8051_golden_model_1.n1271 [9], input_sha_func_33[9]);
  buf(\xm8051_golden_model_1.n1271 [10], input_sha_func_33[10]);
  buf(\xm8051_golden_model_1.n1271 [11], input_sha_func_33[11]);
  buf(\xm8051_golden_model_1.n1271 [12], input_sha_func_33[12]);
  buf(\xm8051_golden_model_1.n1271 [13], input_sha_func_33[13]);
  buf(\xm8051_golden_model_1.n1271 [14], input_sha_func_33[14]);
  buf(\xm8051_golden_model_1.n1271 [15], input_sha_func_33[15]);
  buf(\xm8051_golden_model_1.n1271 [16], input_sha_func_33[16]);
  buf(\xm8051_golden_model_1.n1271 [17], input_sha_func_33[17]);
  buf(\xm8051_golden_model_1.n1271 [18], input_sha_func_33[18]);
  buf(\xm8051_golden_model_1.n1271 [19], input_sha_func_33[19]);
  buf(\xm8051_golden_model_1.n1271 [20], input_sha_func_33[20]);
  buf(\xm8051_golden_model_1.n1271 [21], input_sha_func_33[21]);
  buf(\xm8051_golden_model_1.n1271 [22], input_sha_func_33[22]);
  buf(\xm8051_golden_model_1.n1271 [23], input_sha_func_33[23]);
  buf(\xm8051_golden_model_1.n1271 [24], input_sha_func_33[24]);
  buf(\xm8051_golden_model_1.n1271 [25], input_sha_func_33[25]);
  buf(\xm8051_golden_model_1.n1271 [26], input_sha_func_33[26]);
  buf(\xm8051_golden_model_1.n1271 [27], input_sha_func_33[27]);
  buf(\xm8051_golden_model_1.n1271 [28], input_sha_func_33[28]);
  buf(\xm8051_golden_model_1.n1271 [29], input_sha_func_33[29]);
  buf(\xm8051_golden_model_1.n1271 [30], input_sha_func_33[30]);
  buf(\xm8051_golden_model_1.n1271 [31], input_sha_func_33[31]);
  buf(\xm8051_golden_model_1.n1271 [32], input_sha_func_32[0]);
  buf(\xm8051_golden_model_1.n1271 [33], input_sha_func_32[1]);
  buf(\xm8051_golden_model_1.n1271 [34], input_sha_func_32[2]);
  buf(\xm8051_golden_model_1.n1271 [35], input_sha_func_32[3]);
  buf(\xm8051_golden_model_1.n1271 [36], input_sha_func_32[4]);
  buf(\xm8051_golden_model_1.n1271 [37], input_sha_func_32[5]);
  buf(\xm8051_golden_model_1.n1271 [38], input_sha_func_32[6]);
  buf(\xm8051_golden_model_1.n1271 [39], input_sha_func_32[7]);
  buf(\xm8051_golden_model_1.n1271 [40], input_sha_func_32[8]);
  buf(\xm8051_golden_model_1.n1271 [41], input_sha_func_32[9]);
  buf(\xm8051_golden_model_1.n1271 [42], input_sha_func_32[10]);
  buf(\xm8051_golden_model_1.n1271 [43], input_sha_func_32[11]);
  buf(\xm8051_golden_model_1.n1271 [44], input_sha_func_32[12]);
  buf(\xm8051_golden_model_1.n1271 [45], input_sha_func_32[13]);
  buf(\xm8051_golden_model_1.n1271 [46], input_sha_func_32[14]);
  buf(\xm8051_golden_model_1.n1271 [47], input_sha_func_32[15]);
  buf(\xm8051_golden_model_1.n1271 [48], input_sha_func_32[16]);
  buf(\xm8051_golden_model_1.n1271 [49], input_sha_func_32[17]);
  buf(\xm8051_golden_model_1.n1271 [50], input_sha_func_32[18]);
  buf(\xm8051_golden_model_1.n1271 [51], input_sha_func_32[19]);
  buf(\xm8051_golden_model_1.n1271 [52], input_sha_func_32[20]);
  buf(\xm8051_golden_model_1.n1271 [53], input_sha_func_32[21]);
  buf(\xm8051_golden_model_1.n1271 [54], input_sha_func_32[22]);
  buf(\xm8051_golden_model_1.n1271 [55], input_sha_func_32[23]);
  buf(\xm8051_golden_model_1.n1271 [56], input_sha_func_32[24]);
  buf(\xm8051_golden_model_1.n1271 [57], input_sha_func_32[25]);
  buf(\xm8051_golden_model_1.n1271 [58], input_sha_func_32[26]);
  buf(\xm8051_golden_model_1.n1271 [59], input_sha_func_32[27]);
  buf(\xm8051_golden_model_1.n1271 [60], input_sha_func_32[28]);
  buf(\xm8051_golden_model_1.n1271 [61], input_sha_func_32[29]);
  buf(\xm8051_golden_model_1.n1271 [62], input_sha_func_32[30]);
  buf(\xm8051_golden_model_1.n1271 [63], input_sha_func_32[31]);
  buf(\xm8051_golden_model_1.n1271 [64], input_sha_func_32[32]);
  buf(\xm8051_golden_model_1.n1271 [65], input_sha_func_32[33]);
  buf(\xm8051_golden_model_1.n1271 [66], input_sha_func_32[34]);
  buf(\xm8051_golden_model_1.n1271 [67], input_sha_func_32[35]);
  buf(\xm8051_golden_model_1.n1271 [68], input_sha_func_32[36]);
  buf(\xm8051_golden_model_1.n1271 [69], input_sha_func_32[37]);
  buf(\xm8051_golden_model_1.n1271 [70], input_sha_func_32[38]);
  buf(\xm8051_golden_model_1.n1271 [71], input_sha_func_32[39]);
  buf(\xm8051_golden_model_1.n1271 [72], input_sha_func_32[40]);
  buf(\xm8051_golden_model_1.n1271 [73], input_sha_func_32[41]);
  buf(\xm8051_golden_model_1.n1271 [74], input_sha_func_32[42]);
  buf(\xm8051_golden_model_1.n1271 [75], input_sha_func_32[43]);
  buf(\xm8051_golden_model_1.n1271 [76], input_sha_func_32[44]);
  buf(\xm8051_golden_model_1.n1271 [77], input_sha_func_32[45]);
  buf(\xm8051_golden_model_1.n1271 [78], input_sha_func_32[46]);
  buf(\xm8051_golden_model_1.n1271 [79], input_sha_func_32[47]);
  buf(\xm8051_golden_model_1.n1271 [80], input_sha_func_32[48]);
  buf(\xm8051_golden_model_1.n1271 [81], input_sha_func_32[49]);
  buf(\xm8051_golden_model_1.n1271 [82], input_sha_func_32[50]);
  buf(\xm8051_golden_model_1.n1271 [83], input_sha_func_32[51]);
  buf(\xm8051_golden_model_1.n1271 [84], input_sha_func_32[52]);
  buf(\xm8051_golden_model_1.n1271 [85], input_sha_func_32[53]);
  buf(\xm8051_golden_model_1.n1271 [86], input_sha_func_32[54]);
  buf(\xm8051_golden_model_1.n1271 [87], input_sha_func_32[55]);
  buf(\xm8051_golden_model_1.n1271 [88], input_sha_func_32[56]);
  buf(\xm8051_golden_model_1.n1271 [89], input_sha_func_32[57]);
  buf(\xm8051_golden_model_1.n1271 [90], input_sha_func_32[58]);
  buf(\xm8051_golden_model_1.n1271 [91], input_sha_func_32[59]);
  buf(\xm8051_golden_model_1.n1271 [92], input_sha_func_32[60]);
  buf(\xm8051_golden_model_1.n1271 [93], input_sha_func_32[61]);
  buf(\xm8051_golden_model_1.n1271 [94], input_sha_func_32[62]);
  buf(\xm8051_golden_model_1.n1271 [95], input_sha_func_32[63]);
  buf(\xm8051_golden_model_1.n1271 [96], input_sha_func_31[0]);
  buf(\xm8051_golden_model_1.n1271 [97], input_sha_func_31[1]);
  buf(\xm8051_golden_model_1.n1271 [98], input_sha_func_31[2]);
  buf(\xm8051_golden_model_1.n1271 [99], input_sha_func_31[3]);
  buf(\xm8051_golden_model_1.n1271 [100], input_sha_func_31[4]);
  buf(\xm8051_golden_model_1.n1271 [101], input_sha_func_31[5]);
  buf(\xm8051_golden_model_1.n1271 [102], input_sha_func_31[6]);
  buf(\xm8051_golden_model_1.n1271 [103], input_sha_func_31[7]);
  buf(\xm8051_golden_model_1.n1271 [104], input_sha_func_31[8]);
  buf(\xm8051_golden_model_1.n1271 [105], input_sha_func_31[9]);
  buf(\xm8051_golden_model_1.n1271 [106], input_sha_func_31[10]);
  buf(\xm8051_golden_model_1.n1271 [107], input_sha_func_31[11]);
  buf(\xm8051_golden_model_1.n1271 [108], input_sha_func_31[12]);
  buf(\xm8051_golden_model_1.n1271 [109], input_sha_func_31[13]);
  buf(\xm8051_golden_model_1.n1271 [110], input_sha_func_31[14]);
  buf(\xm8051_golden_model_1.n1271 [111], input_sha_func_31[15]);
  buf(\xm8051_golden_model_1.n1271 [112], input_sha_func_31[16]);
  buf(\xm8051_golden_model_1.n1271 [113], input_sha_func_31[17]);
  buf(\xm8051_golden_model_1.n1271 [114], input_sha_func_31[18]);
  buf(\xm8051_golden_model_1.n1271 [115], input_sha_func_31[19]);
  buf(\xm8051_golden_model_1.n1271 [116], input_sha_func_31[20]);
  buf(\xm8051_golden_model_1.n1271 [117], input_sha_func_31[21]);
  buf(\xm8051_golden_model_1.n1271 [118], input_sha_func_31[22]);
  buf(\xm8051_golden_model_1.n1271 [119], input_sha_func_31[23]);
  buf(\xm8051_golden_model_1.n1271 [120], input_sha_func_31[24]);
  buf(\xm8051_golden_model_1.n1271 [121], input_sha_func_31[25]);
  buf(\xm8051_golden_model_1.n1271 [122], input_sha_func_31[26]);
  buf(\xm8051_golden_model_1.n1271 [123], input_sha_func_31[27]);
  buf(\xm8051_golden_model_1.n1271 [124], input_sha_func_31[28]);
  buf(\xm8051_golden_model_1.n1271 [125], input_sha_func_31[29]);
  buf(\xm8051_golden_model_1.n1271 [126], input_sha_func_31[30]);
  buf(\xm8051_golden_model_1.n1271 [127], input_sha_func_31[31]);
  buf(\xm8051_golden_model_1.n1271 [128], input_sha_func_31[32]);
  buf(\xm8051_golden_model_1.n1271 [129], input_sha_func_31[33]);
  buf(\xm8051_golden_model_1.n1271 [130], input_sha_func_31[34]);
  buf(\xm8051_golden_model_1.n1271 [131], input_sha_func_31[35]);
  buf(\xm8051_golden_model_1.n1271 [132], input_sha_func_31[36]);
  buf(\xm8051_golden_model_1.n1271 [133], input_sha_func_31[37]);
  buf(\xm8051_golden_model_1.n1271 [134], input_sha_func_31[38]);
  buf(\xm8051_golden_model_1.n1271 [135], input_sha_func_31[39]);
  buf(\xm8051_golden_model_1.n1271 [136], input_sha_func_31[40]);
  buf(\xm8051_golden_model_1.n1271 [137], input_sha_func_31[41]);
  buf(\xm8051_golden_model_1.n1271 [138], input_sha_func_31[42]);
  buf(\xm8051_golden_model_1.n1271 [139], input_sha_func_31[43]);
  buf(\xm8051_golden_model_1.n1271 [140], input_sha_func_31[44]);
  buf(\xm8051_golden_model_1.n1271 [141], input_sha_func_31[45]);
  buf(\xm8051_golden_model_1.n1271 [142], input_sha_func_31[46]);
  buf(\xm8051_golden_model_1.n1271 [143], input_sha_func_31[47]);
  buf(\xm8051_golden_model_1.n1271 [144], input_sha_func_31[48]);
  buf(\xm8051_golden_model_1.n1271 [145], input_sha_func_31[49]);
  buf(\xm8051_golden_model_1.n1271 [146], input_sha_func_31[50]);
  buf(\xm8051_golden_model_1.n1271 [147], input_sha_func_31[51]);
  buf(\xm8051_golden_model_1.n1271 [148], input_sha_func_31[52]);
  buf(\xm8051_golden_model_1.n1271 [149], input_sha_func_31[53]);
  buf(\xm8051_golden_model_1.n1271 [150], input_sha_func_31[54]);
  buf(\xm8051_golden_model_1.n1271 [151], input_sha_func_31[55]);
  buf(\xm8051_golden_model_1.n1271 [152], input_sha_func_31[56]);
  buf(\xm8051_golden_model_1.n1271 [153], input_sha_func_31[57]);
  buf(\xm8051_golden_model_1.n1271 [154], input_sha_func_31[58]);
  buf(\xm8051_golden_model_1.n1271 [155], input_sha_func_31[59]);
  buf(\xm8051_golden_model_1.n1271 [156], input_sha_func_31[60]);
  buf(\xm8051_golden_model_1.n1271 [157], input_sha_func_31[61]);
  buf(\xm8051_golden_model_1.n1271 [158], input_sha_func_31[62]);
  buf(\xm8051_golden_model_1.n1271 [159], input_sha_func_31[63]);
  buf(\xm8051_golden_model_1.n0704 [0], sha_rdaddr_gm[0]);
  buf(\xm8051_golden_model_1.n0704 [1], sha_rdaddr_gm[1]);
  buf(\xm8051_golden_model_1.n0704 [2], sha_rdaddr_gm[2]);
  buf(\xm8051_golden_model_1.n0704 [3], sha_rdaddr_gm[3]);
  buf(\xm8051_golden_model_1.n0704 [4], sha_rdaddr_gm[4]);
  buf(\xm8051_golden_model_1.n0704 [5], sha_rdaddr_gm[5]);
  buf(\xm8051_golden_model_1.n0704 [6], sha_rdaddr_gm[6]);
  buf(\xm8051_golden_model_1.n0704 [7], sha_rdaddr_gm[7]);
  buf(\xm8051_golden_model_1.n0704 [8], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0704 [9], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0704 [10], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0704 [11], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0704 [12], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0704 [13], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0704 [14], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0704 [15], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0245 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0245 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0245 [2], \xm8051_golden_model_1.n0473 [2]);
  buf(\xm8051_golden_model_1.n0245 [3], \xm8051_golden_model_1.n0433 [3]);
  buf(\xm8051_golden_model_1.n0245 [4], \xm8051_golden_model_1.n0433 [4]);
  buf(\xm8051_golden_model_1.n0703 [0], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0703 [1], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0703 [2], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0703 [3], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0703 [4], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0703 [5], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0703 [6], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0703 [7], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0703 [8], sha_rdaddr_gm[8]);
  buf(\xm8051_golden_model_1.n0703 [9], sha_rdaddr_gm[9]);
  buf(\xm8051_golden_model_1.n0703 [10], sha_rdaddr_gm[10]);
  buf(\xm8051_golden_model_1.n0703 [11], sha_rdaddr_gm[11]);
  buf(\xm8051_golden_model_1.n0703 [12], sha_rdaddr_gm[12]);
  buf(\xm8051_golden_model_1.n0703 [13], sha_rdaddr_gm[13]);
  buf(\xm8051_golden_model_1.n0703 [14], sha_rdaddr_gm[14]);
  buf(\xm8051_golden_model_1.n0703 [15], sha_rdaddr_gm[15]);
  buf(\xm8051_golden_model_1.n1267 [0], input_sha_func_30[0]);
  buf(\xm8051_golden_model_1.n1267 [1], input_sha_func_30[1]);
  buf(\xm8051_golden_model_1.n1267 [2], input_sha_func_30[2]);
  buf(\xm8051_golden_model_1.n1267 [3], input_sha_func_30[3]);
  buf(\xm8051_golden_model_1.n1267 [4], input_sha_func_30[4]);
  buf(\xm8051_golden_model_1.n1267 [5], input_sha_func_30[5]);
  buf(\xm8051_golden_model_1.n1267 [6], input_sha_func_30[6]);
  buf(\xm8051_golden_model_1.n1267 [7], input_sha_func_30[7]);
  buf(\xm8051_golden_model_1.n1267 [8], input_sha_func_30[8]);
  buf(\xm8051_golden_model_1.n1267 [9], input_sha_func_30[9]);
  buf(\xm8051_golden_model_1.n1267 [10], input_sha_func_30[10]);
  buf(\xm8051_golden_model_1.n1267 [11], input_sha_func_30[11]);
  buf(\xm8051_golden_model_1.n1267 [12], input_sha_func_30[12]);
  buf(\xm8051_golden_model_1.n1267 [13], input_sha_func_30[13]);
  buf(\xm8051_golden_model_1.n1267 [14], input_sha_func_30[14]);
  buf(\xm8051_golden_model_1.n1267 [15], input_sha_func_30[15]);
  buf(\xm8051_golden_model_1.n1267 [16], input_sha_func_30[16]);
  buf(\xm8051_golden_model_1.n1267 [17], input_sha_func_30[17]);
  buf(\xm8051_golden_model_1.n1267 [18], input_sha_func_30[18]);
  buf(\xm8051_golden_model_1.n1267 [19], input_sha_func_30[19]);
  buf(\xm8051_golden_model_1.n1267 [20], input_sha_func_30[20]);
  buf(\xm8051_golden_model_1.n1267 [21], input_sha_func_30[21]);
  buf(\xm8051_golden_model_1.n1267 [22], input_sha_func_30[22]);
  buf(\xm8051_golden_model_1.n1267 [23], input_sha_func_30[23]);
  buf(\xm8051_golden_model_1.n1267 [24], input_sha_func_30[24]);
  buf(\xm8051_golden_model_1.n1267 [25], input_sha_func_30[25]);
  buf(\xm8051_golden_model_1.n1267 [26], input_sha_func_30[26]);
  buf(\xm8051_golden_model_1.n1267 [27], input_sha_func_30[27]);
  buf(\xm8051_golden_model_1.n1267 [28], input_sha_func_30[28]);
  buf(\xm8051_golden_model_1.n1267 [29], input_sha_func_30[29]);
  buf(\xm8051_golden_model_1.n1267 [30], input_sha_func_30[30]);
  buf(\xm8051_golden_model_1.n1267 [31], input_sha_func_30[31]);
  buf(\xm8051_golden_model_1.n1267 [32], input_sha_func_29[0]);
  buf(\xm8051_golden_model_1.n1267 [33], input_sha_func_29[1]);
  buf(\xm8051_golden_model_1.n1267 [34], input_sha_func_29[2]);
  buf(\xm8051_golden_model_1.n1267 [35], input_sha_func_29[3]);
  buf(\xm8051_golden_model_1.n1267 [36], input_sha_func_29[4]);
  buf(\xm8051_golden_model_1.n1267 [37], input_sha_func_29[5]);
  buf(\xm8051_golden_model_1.n1267 [38], input_sha_func_29[6]);
  buf(\xm8051_golden_model_1.n1267 [39], input_sha_func_29[7]);
  buf(\xm8051_golden_model_1.n1267 [40], input_sha_func_29[8]);
  buf(\xm8051_golden_model_1.n1267 [41], input_sha_func_29[9]);
  buf(\xm8051_golden_model_1.n1267 [42], input_sha_func_29[10]);
  buf(\xm8051_golden_model_1.n1267 [43], input_sha_func_29[11]);
  buf(\xm8051_golden_model_1.n1267 [44], input_sha_func_29[12]);
  buf(\xm8051_golden_model_1.n1267 [45], input_sha_func_29[13]);
  buf(\xm8051_golden_model_1.n1267 [46], input_sha_func_29[14]);
  buf(\xm8051_golden_model_1.n1267 [47], input_sha_func_29[15]);
  buf(\xm8051_golden_model_1.n1267 [48], input_sha_func_29[16]);
  buf(\xm8051_golden_model_1.n1267 [49], input_sha_func_29[17]);
  buf(\xm8051_golden_model_1.n1267 [50], input_sha_func_29[18]);
  buf(\xm8051_golden_model_1.n1267 [51], input_sha_func_29[19]);
  buf(\xm8051_golden_model_1.n1267 [52], input_sha_func_29[20]);
  buf(\xm8051_golden_model_1.n1267 [53], input_sha_func_29[21]);
  buf(\xm8051_golden_model_1.n1267 [54], input_sha_func_29[22]);
  buf(\xm8051_golden_model_1.n1267 [55], input_sha_func_29[23]);
  buf(\xm8051_golden_model_1.n1267 [56], input_sha_func_29[24]);
  buf(\xm8051_golden_model_1.n1267 [57], input_sha_func_29[25]);
  buf(\xm8051_golden_model_1.n1267 [58], input_sha_func_29[26]);
  buf(\xm8051_golden_model_1.n1267 [59], input_sha_func_29[27]);
  buf(\xm8051_golden_model_1.n1267 [60], input_sha_func_29[28]);
  buf(\xm8051_golden_model_1.n1267 [61], input_sha_func_29[29]);
  buf(\xm8051_golden_model_1.n1267 [62], input_sha_func_29[30]);
  buf(\xm8051_golden_model_1.n1267 [63], input_sha_func_29[31]);
  buf(\xm8051_golden_model_1.n1267 [64], input_sha_func_29[32]);
  buf(\xm8051_golden_model_1.n1267 [65], input_sha_func_29[33]);
  buf(\xm8051_golden_model_1.n1267 [66], input_sha_func_29[34]);
  buf(\xm8051_golden_model_1.n1267 [67], input_sha_func_29[35]);
  buf(\xm8051_golden_model_1.n1267 [68], input_sha_func_29[36]);
  buf(\xm8051_golden_model_1.n1267 [69], input_sha_func_29[37]);
  buf(\xm8051_golden_model_1.n1267 [70], input_sha_func_29[38]);
  buf(\xm8051_golden_model_1.n1267 [71], input_sha_func_29[39]);
  buf(\xm8051_golden_model_1.n1267 [72], input_sha_func_29[40]);
  buf(\xm8051_golden_model_1.n1267 [73], input_sha_func_29[41]);
  buf(\xm8051_golden_model_1.n1267 [74], input_sha_func_29[42]);
  buf(\xm8051_golden_model_1.n1267 [75], input_sha_func_29[43]);
  buf(\xm8051_golden_model_1.n1267 [76], input_sha_func_29[44]);
  buf(\xm8051_golden_model_1.n1267 [77], input_sha_func_29[45]);
  buf(\xm8051_golden_model_1.n1267 [78], input_sha_func_29[46]);
  buf(\xm8051_golden_model_1.n1267 [79], input_sha_func_29[47]);
  buf(\xm8051_golden_model_1.n1267 [80], input_sha_func_29[48]);
  buf(\xm8051_golden_model_1.n1267 [81], input_sha_func_29[49]);
  buf(\xm8051_golden_model_1.n1267 [82], input_sha_func_29[50]);
  buf(\xm8051_golden_model_1.n1267 [83], input_sha_func_29[51]);
  buf(\xm8051_golden_model_1.n1267 [84], input_sha_func_29[52]);
  buf(\xm8051_golden_model_1.n1267 [85], input_sha_func_29[53]);
  buf(\xm8051_golden_model_1.n1267 [86], input_sha_func_29[54]);
  buf(\xm8051_golden_model_1.n1267 [87], input_sha_func_29[55]);
  buf(\xm8051_golden_model_1.n1267 [88], input_sha_func_29[56]);
  buf(\xm8051_golden_model_1.n1267 [89], input_sha_func_29[57]);
  buf(\xm8051_golden_model_1.n1267 [90], input_sha_func_29[58]);
  buf(\xm8051_golden_model_1.n1267 [91], input_sha_func_29[59]);
  buf(\xm8051_golden_model_1.n1267 [92], input_sha_func_29[60]);
  buf(\xm8051_golden_model_1.n1267 [93], input_sha_func_29[61]);
  buf(\xm8051_golden_model_1.n1267 [94], input_sha_func_29[62]);
  buf(\xm8051_golden_model_1.n1267 [95], input_sha_func_29[63]);
  buf(\xm8051_golden_model_1.n1267 [96], input_sha_func_28[0]);
  buf(\xm8051_golden_model_1.n1267 [97], input_sha_func_28[1]);
  buf(\xm8051_golden_model_1.n1267 [98], input_sha_func_28[2]);
  buf(\xm8051_golden_model_1.n1267 [99], input_sha_func_28[3]);
  buf(\xm8051_golden_model_1.n1267 [100], input_sha_func_28[4]);
  buf(\xm8051_golden_model_1.n1267 [101], input_sha_func_28[5]);
  buf(\xm8051_golden_model_1.n1267 [102], input_sha_func_28[6]);
  buf(\xm8051_golden_model_1.n1267 [103], input_sha_func_28[7]);
  buf(\xm8051_golden_model_1.n1267 [104], input_sha_func_28[8]);
  buf(\xm8051_golden_model_1.n1267 [105], input_sha_func_28[9]);
  buf(\xm8051_golden_model_1.n1267 [106], input_sha_func_28[10]);
  buf(\xm8051_golden_model_1.n1267 [107], input_sha_func_28[11]);
  buf(\xm8051_golden_model_1.n1267 [108], input_sha_func_28[12]);
  buf(\xm8051_golden_model_1.n1267 [109], input_sha_func_28[13]);
  buf(\xm8051_golden_model_1.n1267 [110], input_sha_func_28[14]);
  buf(\xm8051_golden_model_1.n1267 [111], input_sha_func_28[15]);
  buf(\xm8051_golden_model_1.n1267 [112], input_sha_func_28[16]);
  buf(\xm8051_golden_model_1.n1267 [113], input_sha_func_28[17]);
  buf(\xm8051_golden_model_1.n1267 [114], input_sha_func_28[18]);
  buf(\xm8051_golden_model_1.n1267 [115], input_sha_func_28[19]);
  buf(\xm8051_golden_model_1.n1267 [116], input_sha_func_28[20]);
  buf(\xm8051_golden_model_1.n1267 [117], input_sha_func_28[21]);
  buf(\xm8051_golden_model_1.n1267 [118], input_sha_func_28[22]);
  buf(\xm8051_golden_model_1.n1267 [119], input_sha_func_28[23]);
  buf(\xm8051_golden_model_1.n1267 [120], input_sha_func_28[24]);
  buf(\xm8051_golden_model_1.n1267 [121], input_sha_func_28[25]);
  buf(\xm8051_golden_model_1.n1267 [122], input_sha_func_28[26]);
  buf(\xm8051_golden_model_1.n1267 [123], input_sha_func_28[27]);
  buf(\xm8051_golden_model_1.n1267 [124], input_sha_func_28[28]);
  buf(\xm8051_golden_model_1.n1267 [125], input_sha_func_28[29]);
  buf(\xm8051_golden_model_1.n1267 [126], input_sha_func_28[30]);
  buf(\xm8051_golden_model_1.n1267 [127], input_sha_func_28[31]);
  buf(\xm8051_golden_model_1.n1267 [128], input_sha_func_28[32]);
  buf(\xm8051_golden_model_1.n1267 [129], input_sha_func_28[33]);
  buf(\xm8051_golden_model_1.n1267 [130], input_sha_func_28[34]);
  buf(\xm8051_golden_model_1.n1267 [131], input_sha_func_28[35]);
  buf(\xm8051_golden_model_1.n1267 [132], input_sha_func_28[36]);
  buf(\xm8051_golden_model_1.n1267 [133], input_sha_func_28[37]);
  buf(\xm8051_golden_model_1.n1267 [134], input_sha_func_28[38]);
  buf(\xm8051_golden_model_1.n1267 [135], input_sha_func_28[39]);
  buf(\xm8051_golden_model_1.n1267 [136], input_sha_func_28[40]);
  buf(\xm8051_golden_model_1.n1267 [137], input_sha_func_28[41]);
  buf(\xm8051_golden_model_1.n1267 [138], input_sha_func_28[42]);
  buf(\xm8051_golden_model_1.n1267 [139], input_sha_func_28[43]);
  buf(\xm8051_golden_model_1.n1267 [140], input_sha_func_28[44]);
  buf(\xm8051_golden_model_1.n1267 [141], input_sha_func_28[45]);
  buf(\xm8051_golden_model_1.n1267 [142], input_sha_func_28[46]);
  buf(\xm8051_golden_model_1.n1267 [143], input_sha_func_28[47]);
  buf(\xm8051_golden_model_1.n1267 [144], input_sha_func_28[48]);
  buf(\xm8051_golden_model_1.n1267 [145], input_sha_func_28[49]);
  buf(\xm8051_golden_model_1.n1267 [146], input_sha_func_28[50]);
  buf(\xm8051_golden_model_1.n1267 [147], input_sha_func_28[51]);
  buf(\xm8051_golden_model_1.n1267 [148], input_sha_func_28[52]);
  buf(\xm8051_golden_model_1.n1267 [149], input_sha_func_28[53]);
  buf(\xm8051_golden_model_1.n1267 [150], input_sha_func_28[54]);
  buf(\xm8051_golden_model_1.n1267 [151], input_sha_func_28[55]);
  buf(\xm8051_golden_model_1.n1267 [152], input_sha_func_28[56]);
  buf(\xm8051_golden_model_1.n1267 [153], input_sha_func_28[57]);
  buf(\xm8051_golden_model_1.n1267 [154], input_sha_func_28[58]);
  buf(\xm8051_golden_model_1.n1267 [155], input_sha_func_28[59]);
  buf(\xm8051_golden_model_1.n1267 [156], input_sha_func_28[60]);
  buf(\xm8051_golden_model_1.n1267 [157], input_sha_func_28[61]);
  buf(\xm8051_golden_model_1.n1267 [158], input_sha_func_28[62]);
  buf(\xm8051_golden_model_1.n1267 [159], input_sha_func_28[63]);
  buf(\xm8051_golden_model_1.n1263 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n1263 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n1263 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n1263 [3], \xm8051_golden_model_1.sha_bytes_processed [3]);
  buf(\xm8051_golden_model_1.n1263 [4], \xm8051_golden_model_1.sha_bytes_processed [4]);
  buf(\xm8051_golden_model_1.n1263 [5], \xm8051_golden_model_1.sha_bytes_processed [5]);
  buf(\xm8051_golden_model_1.n1263 [6], \xm8051_golden_model_1.sha_bytes_processed_0b [6]);
  buf(\xm8051_golden_model_1.n1263 [7], \xm8051_golden_model_1.sha_bytes_processed_0b [7]);
  buf(\xm8051_golden_model_1.n1263 [8], \xm8051_golden_model_1.sha_bytes_processed_0b [8]);
  buf(\xm8051_golden_model_1.n1263 [9], \xm8051_golden_model_1.sha_bytes_processed_0b [9]);
  buf(\xm8051_golden_model_1.n1263 [10], \xm8051_golden_model_1.sha_bytes_processed_0b [10]);
  buf(\xm8051_golden_model_1.n1263 [11], \xm8051_golden_model_1.sha_bytes_processed_0b [11]);
  buf(\xm8051_golden_model_1.n1263 [12], \xm8051_golden_model_1.sha_bytes_processed_0b [12]);
  buf(\xm8051_golden_model_1.n1263 [13], \xm8051_golden_model_1.sha_bytes_processed_0b [13]);
  buf(\xm8051_golden_model_1.n1263 [14], \xm8051_golden_model_1.sha_bytes_processed_0b [14]);
  buf(\xm8051_golden_model_1.n1263 [15], \xm8051_golden_model_1.sha_bytes_processed_0b [15]);
  buf(\xm8051_golden_model_1.n1262 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n1262 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n1262 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n1262 [3], \xm8051_golden_model_1.sha_bytes_processed [3]);
  buf(\xm8051_golden_model_1.n1262 [4], \xm8051_golden_model_1.sha_bytes_processed [4]);
  buf(\xm8051_golden_model_1.n1262 [5], \xm8051_golden_model_1.sha_bytes_processed [5]);
  buf(\xm8051_golden_model_1.n0233 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0233 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0233 [2], \xm8051_golden_model_1.n0463 [2]);
  buf(\xm8051_golden_model_1.n0233 [3], \xm8051_golden_model_1.n0423 [3]);
  buf(\xm8051_golden_model_1.n0233 [4], \xm8051_golden_model_1.n0423 [4]);
  buf(\xm8051_golden_model_1.n0691 [0], \xm8051_golden_model_1.sha_len [8]);
  buf(\xm8051_golden_model_1.n0691 [1], \xm8051_golden_model_1.sha_len [9]);
  buf(\xm8051_golden_model_1.n0691 [2], \xm8051_golden_model_1.sha_len [10]);
  buf(\xm8051_golden_model_1.n0691 [3], \xm8051_golden_model_1.sha_len [11]);
  buf(\xm8051_golden_model_1.n0691 [4], \xm8051_golden_model_1.sha_len [12]);
  buf(\xm8051_golden_model_1.n0691 [5], \xm8051_golden_model_1.sha_len [13]);
  buf(\xm8051_golden_model_1.n0691 [6], \xm8051_golden_model_1.sha_len [14]);
  buf(\xm8051_golden_model_1.n0691 [7], \xm8051_golden_model_1.sha_len [15]);
  buf(\xm8051_golden_model_1.n0690 [0], \xm8051_golden_model_1.sha_len [0]);
  buf(\xm8051_golden_model_1.n0690 [1], \xm8051_golden_model_1.sha_len [1]);
  buf(\xm8051_golden_model_1.n0690 [2], \xm8051_golden_model_1.sha_len [2]);
  buf(\xm8051_golden_model_1.n0690 [3], \xm8051_golden_model_1.sha_len [3]);
  buf(\xm8051_golden_model_1.n0690 [4], \xm8051_golden_model_1.sha_len [4]);
  buf(\xm8051_golden_model_1.n0690 [5], \xm8051_golden_model_1.sha_len [5]);
  buf(\xm8051_golden_model_1.n0690 [6], \xm8051_golden_model_1.sha_len [6]);
  buf(\xm8051_golden_model_1.n0690 [7], \xm8051_golden_model_1.sha_len [7]);
  buf(\xm8051_golden_model_1.n1256 [0], input_sha_func_27[0]);
  buf(\xm8051_golden_model_1.n1256 [1], input_sha_func_27[1]);
  buf(\xm8051_golden_model_1.n1256 [2], input_sha_func_27[2]);
  buf(\xm8051_golden_model_1.n1256 [3], input_sha_func_27[3]);
  buf(\xm8051_golden_model_1.n1256 [4], input_sha_func_27[4]);
  buf(\xm8051_golden_model_1.n1256 [5], input_sha_func_27[5]);
  buf(\xm8051_golden_model_1.n1256 [6], input_sha_func_27[6]);
  buf(\xm8051_golden_model_1.n1256 [7], input_sha_func_27[7]);
  buf(\xm8051_golden_model_1.n1256 [8], input_sha_func_27[8]);
  buf(\xm8051_golden_model_1.n1256 [9], input_sha_func_27[9]);
  buf(\xm8051_golden_model_1.n1256 [10], input_sha_func_27[10]);
  buf(\xm8051_golden_model_1.n1256 [11], input_sha_func_27[11]);
  buf(\xm8051_golden_model_1.n1256 [12], input_sha_func_27[12]);
  buf(\xm8051_golden_model_1.n1256 [13], input_sha_func_27[13]);
  buf(\xm8051_golden_model_1.n1256 [14], input_sha_func_27[14]);
  buf(\xm8051_golden_model_1.n1256 [15], input_sha_func_27[15]);
  buf(\xm8051_golden_model_1.n1256 [16], input_sha_func_27[16]);
  buf(\xm8051_golden_model_1.n1256 [17], input_sha_func_27[17]);
  buf(\xm8051_golden_model_1.n1256 [18], input_sha_func_27[18]);
  buf(\xm8051_golden_model_1.n1256 [19], input_sha_func_27[19]);
  buf(\xm8051_golden_model_1.n1256 [20], input_sha_func_27[20]);
  buf(\xm8051_golden_model_1.n1256 [21], input_sha_func_27[21]);
  buf(\xm8051_golden_model_1.n1256 [22], input_sha_func_27[22]);
  buf(\xm8051_golden_model_1.n1256 [23], input_sha_func_27[23]);
  buf(\xm8051_golden_model_1.n1256 [24], input_sha_func_27[24]);
  buf(\xm8051_golden_model_1.n1256 [25], input_sha_func_27[25]);
  buf(\xm8051_golden_model_1.n1256 [26], input_sha_func_27[26]);
  buf(\xm8051_golden_model_1.n1256 [27], input_sha_func_27[27]);
  buf(\xm8051_golden_model_1.n1256 [28], input_sha_func_27[28]);
  buf(\xm8051_golden_model_1.n1256 [29], input_sha_func_27[29]);
  buf(\xm8051_golden_model_1.n1256 [30], input_sha_func_27[30]);
  buf(\xm8051_golden_model_1.n1256 [31], input_sha_func_27[31]);
  buf(\xm8051_golden_model_1.n1256 [32], input_sha_func_26[0]);
  buf(\xm8051_golden_model_1.n1256 [33], input_sha_func_26[1]);
  buf(\xm8051_golden_model_1.n1256 [34], input_sha_func_26[2]);
  buf(\xm8051_golden_model_1.n1256 [35], input_sha_func_26[3]);
  buf(\xm8051_golden_model_1.n1256 [36], input_sha_func_26[4]);
  buf(\xm8051_golden_model_1.n1256 [37], input_sha_func_26[5]);
  buf(\xm8051_golden_model_1.n1256 [38], input_sha_func_26[6]);
  buf(\xm8051_golden_model_1.n1256 [39], input_sha_func_26[7]);
  buf(\xm8051_golden_model_1.n1256 [40], input_sha_func_26[8]);
  buf(\xm8051_golden_model_1.n1256 [41], input_sha_func_26[9]);
  buf(\xm8051_golden_model_1.n1256 [42], input_sha_func_26[10]);
  buf(\xm8051_golden_model_1.n1256 [43], input_sha_func_26[11]);
  buf(\xm8051_golden_model_1.n1256 [44], input_sha_func_26[12]);
  buf(\xm8051_golden_model_1.n1256 [45], input_sha_func_26[13]);
  buf(\xm8051_golden_model_1.n1256 [46], input_sha_func_26[14]);
  buf(\xm8051_golden_model_1.n1256 [47], input_sha_func_26[15]);
  buf(\xm8051_golden_model_1.n1256 [48], input_sha_func_26[16]);
  buf(\xm8051_golden_model_1.n1256 [49], input_sha_func_26[17]);
  buf(\xm8051_golden_model_1.n1256 [50], input_sha_func_26[18]);
  buf(\xm8051_golden_model_1.n1256 [51], input_sha_func_26[19]);
  buf(\xm8051_golden_model_1.n1256 [52], input_sha_func_26[20]);
  buf(\xm8051_golden_model_1.n1256 [53], input_sha_func_26[21]);
  buf(\xm8051_golden_model_1.n1256 [54], input_sha_func_26[22]);
  buf(\xm8051_golden_model_1.n1256 [55], input_sha_func_26[23]);
  buf(\xm8051_golden_model_1.n1256 [56], input_sha_func_26[24]);
  buf(\xm8051_golden_model_1.n1256 [57], input_sha_func_26[25]);
  buf(\xm8051_golden_model_1.n1256 [58], input_sha_func_26[26]);
  buf(\xm8051_golden_model_1.n1256 [59], input_sha_func_26[27]);
  buf(\xm8051_golden_model_1.n1256 [60], input_sha_func_26[28]);
  buf(\xm8051_golden_model_1.n1256 [61], input_sha_func_26[29]);
  buf(\xm8051_golden_model_1.n1256 [62], input_sha_func_26[30]);
  buf(\xm8051_golden_model_1.n1256 [63], input_sha_func_26[31]);
  buf(\xm8051_golden_model_1.n1256 [64], input_sha_func_26[32]);
  buf(\xm8051_golden_model_1.n1256 [65], input_sha_func_26[33]);
  buf(\xm8051_golden_model_1.n1256 [66], input_sha_func_26[34]);
  buf(\xm8051_golden_model_1.n1256 [67], input_sha_func_26[35]);
  buf(\xm8051_golden_model_1.n1256 [68], input_sha_func_26[36]);
  buf(\xm8051_golden_model_1.n1256 [69], input_sha_func_26[37]);
  buf(\xm8051_golden_model_1.n1256 [70], input_sha_func_26[38]);
  buf(\xm8051_golden_model_1.n1256 [71], input_sha_func_26[39]);
  buf(\xm8051_golden_model_1.n1256 [72], input_sha_func_26[40]);
  buf(\xm8051_golden_model_1.n1256 [73], input_sha_func_26[41]);
  buf(\xm8051_golden_model_1.n1256 [74], input_sha_func_26[42]);
  buf(\xm8051_golden_model_1.n1256 [75], input_sha_func_26[43]);
  buf(\xm8051_golden_model_1.n1256 [76], input_sha_func_26[44]);
  buf(\xm8051_golden_model_1.n1256 [77], input_sha_func_26[45]);
  buf(\xm8051_golden_model_1.n1256 [78], input_sha_func_26[46]);
  buf(\xm8051_golden_model_1.n1256 [79], input_sha_func_26[47]);
  buf(\xm8051_golden_model_1.n1256 [80], input_sha_func_26[48]);
  buf(\xm8051_golden_model_1.n1256 [81], input_sha_func_26[49]);
  buf(\xm8051_golden_model_1.n1256 [82], input_sha_func_26[50]);
  buf(\xm8051_golden_model_1.n1256 [83], input_sha_func_26[51]);
  buf(\xm8051_golden_model_1.n1256 [84], input_sha_func_26[52]);
  buf(\xm8051_golden_model_1.n1256 [85], input_sha_func_26[53]);
  buf(\xm8051_golden_model_1.n1256 [86], input_sha_func_26[54]);
  buf(\xm8051_golden_model_1.n1256 [87], input_sha_func_26[55]);
  buf(\xm8051_golden_model_1.n1256 [88], input_sha_func_26[56]);
  buf(\xm8051_golden_model_1.n1256 [89], input_sha_func_26[57]);
  buf(\xm8051_golden_model_1.n1256 [90], input_sha_func_26[58]);
  buf(\xm8051_golden_model_1.n1256 [91], input_sha_func_26[59]);
  buf(\xm8051_golden_model_1.n1256 [92], input_sha_func_26[60]);
  buf(\xm8051_golden_model_1.n1256 [93], input_sha_func_26[61]);
  buf(\xm8051_golden_model_1.n1256 [94], input_sha_func_26[62]);
  buf(\xm8051_golden_model_1.n1256 [95], input_sha_func_26[63]);
  buf(\xm8051_golden_model_1.n1256 [96], input_sha_func_25[0]);
  buf(\xm8051_golden_model_1.n1256 [97], input_sha_func_25[1]);
  buf(\xm8051_golden_model_1.n1256 [98], input_sha_func_25[2]);
  buf(\xm8051_golden_model_1.n1256 [99], input_sha_func_25[3]);
  buf(\xm8051_golden_model_1.n1256 [100], input_sha_func_25[4]);
  buf(\xm8051_golden_model_1.n1256 [101], input_sha_func_25[5]);
  buf(\xm8051_golden_model_1.n1256 [102], input_sha_func_25[6]);
  buf(\xm8051_golden_model_1.n1256 [103], input_sha_func_25[7]);
  buf(\xm8051_golden_model_1.n1256 [104], input_sha_func_25[8]);
  buf(\xm8051_golden_model_1.n1256 [105], input_sha_func_25[9]);
  buf(\xm8051_golden_model_1.n1256 [106], input_sha_func_25[10]);
  buf(\xm8051_golden_model_1.n1256 [107], input_sha_func_25[11]);
  buf(\xm8051_golden_model_1.n1256 [108], input_sha_func_25[12]);
  buf(\xm8051_golden_model_1.n1256 [109], input_sha_func_25[13]);
  buf(\xm8051_golden_model_1.n1256 [110], input_sha_func_25[14]);
  buf(\xm8051_golden_model_1.n1256 [111], input_sha_func_25[15]);
  buf(\xm8051_golden_model_1.n1256 [112], input_sha_func_25[16]);
  buf(\xm8051_golden_model_1.n1256 [113], input_sha_func_25[17]);
  buf(\xm8051_golden_model_1.n1256 [114], input_sha_func_25[18]);
  buf(\xm8051_golden_model_1.n1256 [115], input_sha_func_25[19]);
  buf(\xm8051_golden_model_1.n1256 [116], input_sha_func_25[20]);
  buf(\xm8051_golden_model_1.n1256 [117], input_sha_func_25[21]);
  buf(\xm8051_golden_model_1.n1256 [118], input_sha_func_25[22]);
  buf(\xm8051_golden_model_1.n1256 [119], input_sha_func_25[23]);
  buf(\xm8051_golden_model_1.n1256 [120], input_sha_func_25[24]);
  buf(\xm8051_golden_model_1.n1256 [121], input_sha_func_25[25]);
  buf(\xm8051_golden_model_1.n1256 [122], input_sha_func_25[26]);
  buf(\xm8051_golden_model_1.n1256 [123], input_sha_func_25[27]);
  buf(\xm8051_golden_model_1.n1256 [124], input_sha_func_25[28]);
  buf(\xm8051_golden_model_1.n1256 [125], input_sha_func_25[29]);
  buf(\xm8051_golden_model_1.n1256 [126], input_sha_func_25[30]);
  buf(\xm8051_golden_model_1.n1256 [127], input_sha_func_25[31]);
  buf(\xm8051_golden_model_1.n1256 [128], input_sha_func_25[32]);
  buf(\xm8051_golden_model_1.n1256 [129], input_sha_func_25[33]);
  buf(\xm8051_golden_model_1.n1256 [130], input_sha_func_25[34]);
  buf(\xm8051_golden_model_1.n1256 [131], input_sha_func_25[35]);
  buf(\xm8051_golden_model_1.n1256 [132], input_sha_func_25[36]);
  buf(\xm8051_golden_model_1.n1256 [133], input_sha_func_25[37]);
  buf(\xm8051_golden_model_1.n1256 [134], input_sha_func_25[38]);
  buf(\xm8051_golden_model_1.n1256 [135], input_sha_func_25[39]);
  buf(\xm8051_golden_model_1.n1256 [136], input_sha_func_25[40]);
  buf(\xm8051_golden_model_1.n1256 [137], input_sha_func_25[41]);
  buf(\xm8051_golden_model_1.n1256 [138], input_sha_func_25[42]);
  buf(\xm8051_golden_model_1.n1256 [139], input_sha_func_25[43]);
  buf(\xm8051_golden_model_1.n1256 [140], input_sha_func_25[44]);
  buf(\xm8051_golden_model_1.n1256 [141], input_sha_func_25[45]);
  buf(\xm8051_golden_model_1.n1256 [142], input_sha_func_25[46]);
  buf(\xm8051_golden_model_1.n1256 [143], input_sha_func_25[47]);
  buf(\xm8051_golden_model_1.n1256 [144], input_sha_func_25[48]);
  buf(\xm8051_golden_model_1.n1256 [145], input_sha_func_25[49]);
  buf(\xm8051_golden_model_1.n1256 [146], input_sha_func_25[50]);
  buf(\xm8051_golden_model_1.n1256 [147], input_sha_func_25[51]);
  buf(\xm8051_golden_model_1.n1256 [148], input_sha_func_25[52]);
  buf(\xm8051_golden_model_1.n1256 [149], input_sha_func_25[53]);
  buf(\xm8051_golden_model_1.n1256 [150], input_sha_func_25[54]);
  buf(\xm8051_golden_model_1.n1256 [151], input_sha_func_25[55]);
  buf(\xm8051_golden_model_1.n1256 [152], input_sha_func_25[56]);
  buf(\xm8051_golden_model_1.n1256 [153], input_sha_func_25[57]);
  buf(\xm8051_golden_model_1.n1256 [154], input_sha_func_25[58]);
  buf(\xm8051_golden_model_1.n1256 [155], input_sha_func_25[59]);
  buf(\xm8051_golden_model_1.n1256 [156], input_sha_func_25[60]);
  buf(\xm8051_golden_model_1.n1256 [157], input_sha_func_25[61]);
  buf(\xm8051_golden_model_1.n1256 [158], input_sha_func_25[62]);
  buf(\xm8051_golden_model_1.n1256 [159], input_sha_func_25[63]);
  buf(\xm8051_golden_model_1.n1254 [0], input_aes_func_24[0]);
  buf(\xm8051_golden_model_1.n1254 [1], input_aes_func_24[1]);
  buf(\xm8051_golden_model_1.n1254 [2], input_aes_func_24[2]);
  buf(\xm8051_golden_model_1.n1254 [3], input_aes_func_24[3]);
  buf(\xm8051_golden_model_1.n1254 [4], input_aes_func_24[4]);
  buf(\xm8051_golden_model_1.n1254 [5], input_aes_func_24[5]);
  buf(\xm8051_golden_model_1.n1254 [6], input_aes_func_24[6]);
  buf(\xm8051_golden_model_1.n1254 [7], input_aes_func_24[7]);
  buf(\xm8051_golden_model_1.n1254 [8], input_aes_func_24[8]);
  buf(\xm8051_golden_model_1.n1254 [9], input_aes_func_24[9]);
  buf(\xm8051_golden_model_1.n1254 [10], input_aes_func_24[10]);
  buf(\xm8051_golden_model_1.n1254 [11], input_aes_func_24[11]);
  buf(\xm8051_golden_model_1.n1254 [12], input_aes_func_24[12]);
  buf(\xm8051_golden_model_1.n1254 [13], input_aes_func_24[13]);
  buf(\xm8051_golden_model_1.n1254 [14], input_aes_func_24[14]);
  buf(\xm8051_golden_model_1.n1254 [15], input_aes_func_24[15]);
  buf(\xm8051_golden_model_1.n1254 [16], input_aes_func_24[16]);
  buf(\xm8051_golden_model_1.n1254 [17], input_aes_func_24[17]);
  buf(\xm8051_golden_model_1.n1254 [18], input_aes_func_24[18]);
  buf(\xm8051_golden_model_1.n1254 [19], input_aes_func_24[19]);
  buf(\xm8051_golden_model_1.n1254 [20], input_aes_func_24[20]);
  buf(\xm8051_golden_model_1.n1254 [21], input_aes_func_24[21]);
  buf(\xm8051_golden_model_1.n1254 [22], input_aes_func_24[22]);
  buf(\xm8051_golden_model_1.n1254 [23], input_aes_func_24[23]);
  buf(\xm8051_golden_model_1.n1254 [24], input_aes_func_24[24]);
  buf(\xm8051_golden_model_1.n1254 [25], input_aes_func_24[25]);
  buf(\xm8051_golden_model_1.n1254 [26], input_aes_func_24[26]);
  buf(\xm8051_golden_model_1.n1254 [27], input_aes_func_24[27]);
  buf(\xm8051_golden_model_1.n1254 [28], input_aes_func_24[28]);
  buf(\xm8051_golden_model_1.n1254 [29], input_aes_func_24[29]);
  buf(\xm8051_golden_model_1.n1254 [30], input_aes_func_24[30]);
  buf(\xm8051_golden_model_1.n1254 [31], input_aes_func_24[31]);
  buf(\xm8051_golden_model_1.n1254 [32], input_aes_func_24[32]);
  buf(\xm8051_golden_model_1.n1254 [33], input_aes_func_24[33]);
  buf(\xm8051_golden_model_1.n1254 [34], input_aes_func_24[34]);
  buf(\xm8051_golden_model_1.n1254 [35], input_aes_func_24[35]);
  buf(\xm8051_golden_model_1.n1254 [36], input_aes_func_24[36]);
  buf(\xm8051_golden_model_1.n1254 [37], input_aes_func_24[37]);
  buf(\xm8051_golden_model_1.n1254 [38], input_aes_func_24[38]);
  buf(\xm8051_golden_model_1.n1254 [39], input_aes_func_24[39]);
  buf(\xm8051_golden_model_1.n1254 [40], input_aes_func_24[40]);
  buf(\xm8051_golden_model_1.n1254 [41], input_aes_func_24[41]);
  buf(\xm8051_golden_model_1.n1254 [42], input_aes_func_24[42]);
  buf(\xm8051_golden_model_1.n1254 [43], input_aes_func_24[43]);
  buf(\xm8051_golden_model_1.n1254 [44], input_aes_func_24[44]);
  buf(\xm8051_golden_model_1.n1254 [45], input_aes_func_24[45]);
  buf(\xm8051_golden_model_1.n1254 [46], input_aes_func_24[46]);
  buf(\xm8051_golden_model_1.n1254 [47], input_aes_func_24[47]);
  buf(\xm8051_golden_model_1.n1254 [48], input_aes_func_24[48]);
  buf(\xm8051_golden_model_1.n1254 [49], input_aes_func_24[49]);
  buf(\xm8051_golden_model_1.n1254 [50], input_aes_func_24[50]);
  buf(\xm8051_golden_model_1.n1254 [51], input_aes_func_24[51]);
  buf(\xm8051_golden_model_1.n1254 [52], input_aes_func_24[52]);
  buf(\xm8051_golden_model_1.n1254 [53], input_aes_func_24[53]);
  buf(\xm8051_golden_model_1.n1254 [54], input_aes_func_24[54]);
  buf(\xm8051_golden_model_1.n1254 [55], input_aes_func_24[55]);
  buf(\xm8051_golden_model_1.n1254 [56], input_aes_func_24[56]);
  buf(\xm8051_golden_model_1.n1254 [57], input_aes_func_24[57]);
  buf(\xm8051_golden_model_1.n1254 [58], input_aes_func_24[58]);
  buf(\xm8051_golden_model_1.n1254 [59], input_aes_func_24[59]);
  buf(\xm8051_golden_model_1.n1254 [60], input_aes_func_24[60]);
  buf(\xm8051_golden_model_1.n1254 [61], input_aes_func_24[61]);
  buf(\xm8051_golden_model_1.n1254 [62], input_aes_func_24[62]);
  buf(\xm8051_golden_model_1.n1254 [63], input_aes_func_24[63]);
  buf(\xm8051_golden_model_1.n1254 [64], input_aes_func_23[0]);
  buf(\xm8051_golden_model_1.n1254 [65], input_aes_func_23[1]);
  buf(\xm8051_golden_model_1.n1254 [66], input_aes_func_23[2]);
  buf(\xm8051_golden_model_1.n1254 [67], input_aes_func_23[3]);
  buf(\xm8051_golden_model_1.n1254 [68], input_aes_func_23[4]);
  buf(\xm8051_golden_model_1.n1254 [69], input_aes_func_23[5]);
  buf(\xm8051_golden_model_1.n1254 [70], input_aes_func_23[6]);
  buf(\xm8051_golden_model_1.n1254 [71], input_aes_func_23[7]);
  buf(\xm8051_golden_model_1.n1254 [72], input_aes_func_23[8]);
  buf(\xm8051_golden_model_1.n1254 [73], input_aes_func_23[9]);
  buf(\xm8051_golden_model_1.n1254 [74], input_aes_func_23[10]);
  buf(\xm8051_golden_model_1.n1254 [75], input_aes_func_23[11]);
  buf(\xm8051_golden_model_1.n1254 [76], input_aes_func_23[12]);
  buf(\xm8051_golden_model_1.n1254 [77], input_aes_func_23[13]);
  buf(\xm8051_golden_model_1.n1254 [78], input_aes_func_23[14]);
  buf(\xm8051_golden_model_1.n1254 [79], input_aes_func_23[15]);
  buf(\xm8051_golden_model_1.n1254 [80], input_aes_func_23[16]);
  buf(\xm8051_golden_model_1.n1254 [81], input_aes_func_23[17]);
  buf(\xm8051_golden_model_1.n1254 [82], input_aes_func_23[18]);
  buf(\xm8051_golden_model_1.n1254 [83], input_aes_func_23[19]);
  buf(\xm8051_golden_model_1.n1254 [84], input_aes_func_23[20]);
  buf(\xm8051_golden_model_1.n1254 [85], input_aes_func_23[21]);
  buf(\xm8051_golden_model_1.n1254 [86], input_aes_func_23[22]);
  buf(\xm8051_golden_model_1.n1254 [87], input_aes_func_23[23]);
  buf(\xm8051_golden_model_1.n1254 [88], input_aes_func_23[24]);
  buf(\xm8051_golden_model_1.n1254 [89], input_aes_func_23[25]);
  buf(\xm8051_golden_model_1.n1254 [90], input_aes_func_23[26]);
  buf(\xm8051_golden_model_1.n1254 [91], input_aes_func_23[27]);
  buf(\xm8051_golden_model_1.n1254 [92], input_aes_func_23[28]);
  buf(\xm8051_golden_model_1.n1254 [93], input_aes_func_23[29]);
  buf(\xm8051_golden_model_1.n1254 [94], input_aes_func_23[30]);
  buf(\xm8051_golden_model_1.n1254 [95], input_aes_func_23[31]);
  buf(\xm8051_golden_model_1.n1254 [96], input_aes_func_23[32]);
  buf(\xm8051_golden_model_1.n1254 [97], input_aes_func_23[33]);
  buf(\xm8051_golden_model_1.n1254 [98], input_aes_func_23[34]);
  buf(\xm8051_golden_model_1.n1254 [99], input_aes_func_23[35]);
  buf(\xm8051_golden_model_1.n1254 [100], input_aes_func_23[36]);
  buf(\xm8051_golden_model_1.n1254 [101], input_aes_func_23[37]);
  buf(\xm8051_golden_model_1.n1254 [102], input_aes_func_23[38]);
  buf(\xm8051_golden_model_1.n1254 [103], input_aes_func_23[39]);
  buf(\xm8051_golden_model_1.n1254 [104], input_aes_func_23[40]);
  buf(\xm8051_golden_model_1.n1254 [105], input_aes_func_23[41]);
  buf(\xm8051_golden_model_1.n1254 [106], input_aes_func_23[42]);
  buf(\xm8051_golden_model_1.n1254 [107], input_aes_func_23[43]);
  buf(\xm8051_golden_model_1.n1254 [108], input_aes_func_23[44]);
  buf(\xm8051_golden_model_1.n1254 [109], input_aes_func_23[45]);
  buf(\xm8051_golden_model_1.n1254 [110], input_aes_func_23[46]);
  buf(\xm8051_golden_model_1.n1254 [111], input_aes_func_23[47]);
  buf(\xm8051_golden_model_1.n1254 [112], input_aes_func_23[48]);
  buf(\xm8051_golden_model_1.n1254 [113], input_aes_func_23[49]);
  buf(\xm8051_golden_model_1.n1254 [114], input_aes_func_23[50]);
  buf(\xm8051_golden_model_1.n1254 [115], input_aes_func_23[51]);
  buf(\xm8051_golden_model_1.n1254 [116], input_aes_func_23[52]);
  buf(\xm8051_golden_model_1.n1254 [117], input_aes_func_23[53]);
  buf(\xm8051_golden_model_1.n1254 [118], input_aes_func_23[54]);
  buf(\xm8051_golden_model_1.n1254 [119], input_aes_func_23[55]);
  buf(\xm8051_golden_model_1.n1254 [120], input_aes_func_23[56]);
  buf(\xm8051_golden_model_1.n1254 [121], input_aes_func_23[57]);
  buf(\xm8051_golden_model_1.n1254 [122], input_aes_func_23[58]);
  buf(\xm8051_golden_model_1.n1254 [123], input_aes_func_23[59]);
  buf(\xm8051_golden_model_1.n1254 [124], input_aes_func_23[60]);
  buf(\xm8051_golden_model_1.n1254 [125], input_aes_func_23[61]);
  buf(\xm8051_golden_model_1.n1254 [126], input_aes_func_23[62]);
  buf(\xm8051_golden_model_1.n1254 [127], input_aes_func_23[63]);
  buf(\xm8051_golden_model_1.n0218 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0218 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0218 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n0218 [3], \xm8051_golden_model_1.sha_bytes_processed [3]);
  buf(\xm8051_golden_model_1.n0218 [4], \xm8051_golden_model_1.n0413 [4]);
  buf(\xm8051_golden_model_1.n1250 [0], input_sha_func_22[0]);
  buf(\xm8051_golden_model_1.n1250 [1], input_sha_func_22[1]);
  buf(\xm8051_golden_model_1.n1250 [2], input_sha_func_22[2]);
  buf(\xm8051_golden_model_1.n1250 [3], input_sha_func_22[3]);
  buf(\xm8051_golden_model_1.n1250 [4], input_sha_func_22[4]);
  buf(\xm8051_golden_model_1.n1250 [5], input_sha_func_22[5]);
  buf(\xm8051_golden_model_1.n1250 [6], input_sha_func_22[6]);
  buf(\xm8051_golden_model_1.n1250 [7], input_sha_func_22[7]);
  buf(\xm8051_golden_model_1.n1250 [8], input_sha_func_22[8]);
  buf(\xm8051_golden_model_1.n1250 [9], input_sha_func_22[9]);
  buf(\xm8051_golden_model_1.n1250 [10], input_sha_func_22[10]);
  buf(\xm8051_golden_model_1.n1250 [11], input_sha_func_22[11]);
  buf(\xm8051_golden_model_1.n1250 [12], input_sha_func_22[12]);
  buf(\xm8051_golden_model_1.n1250 [13], input_sha_func_22[13]);
  buf(\xm8051_golden_model_1.n1250 [14], input_sha_func_22[14]);
  buf(\xm8051_golden_model_1.n1250 [15], input_sha_func_22[15]);
  buf(\xm8051_golden_model_1.n1250 [16], input_sha_func_22[16]);
  buf(\xm8051_golden_model_1.n1250 [17], input_sha_func_22[17]);
  buf(\xm8051_golden_model_1.n1250 [18], input_sha_func_22[18]);
  buf(\xm8051_golden_model_1.n1250 [19], input_sha_func_22[19]);
  buf(\xm8051_golden_model_1.n1250 [20], input_sha_func_22[20]);
  buf(\xm8051_golden_model_1.n1250 [21], input_sha_func_22[21]);
  buf(\xm8051_golden_model_1.n1250 [22], input_sha_func_22[22]);
  buf(\xm8051_golden_model_1.n1250 [23], input_sha_func_22[23]);
  buf(\xm8051_golden_model_1.n1250 [24], input_sha_func_22[24]);
  buf(\xm8051_golden_model_1.n1250 [25], input_sha_func_22[25]);
  buf(\xm8051_golden_model_1.n1250 [26], input_sha_func_22[26]);
  buf(\xm8051_golden_model_1.n1250 [27], input_sha_func_22[27]);
  buf(\xm8051_golden_model_1.n1250 [28], input_sha_func_22[28]);
  buf(\xm8051_golden_model_1.n1250 [29], input_sha_func_22[29]);
  buf(\xm8051_golden_model_1.n1250 [30], input_sha_func_22[30]);
  buf(\xm8051_golden_model_1.n1250 [31], input_sha_func_22[31]);
  buf(\xm8051_golden_model_1.n1250 [32], input_sha_func_21[0]);
  buf(\xm8051_golden_model_1.n1250 [33], input_sha_func_21[1]);
  buf(\xm8051_golden_model_1.n1250 [34], input_sha_func_21[2]);
  buf(\xm8051_golden_model_1.n1250 [35], input_sha_func_21[3]);
  buf(\xm8051_golden_model_1.n1250 [36], input_sha_func_21[4]);
  buf(\xm8051_golden_model_1.n1250 [37], input_sha_func_21[5]);
  buf(\xm8051_golden_model_1.n1250 [38], input_sha_func_21[6]);
  buf(\xm8051_golden_model_1.n1250 [39], input_sha_func_21[7]);
  buf(\xm8051_golden_model_1.n1250 [40], input_sha_func_21[8]);
  buf(\xm8051_golden_model_1.n1250 [41], input_sha_func_21[9]);
  buf(\xm8051_golden_model_1.n1250 [42], input_sha_func_21[10]);
  buf(\xm8051_golden_model_1.n1250 [43], input_sha_func_21[11]);
  buf(\xm8051_golden_model_1.n1250 [44], input_sha_func_21[12]);
  buf(\xm8051_golden_model_1.n1250 [45], input_sha_func_21[13]);
  buf(\xm8051_golden_model_1.n1250 [46], input_sha_func_21[14]);
  buf(\xm8051_golden_model_1.n1250 [47], input_sha_func_21[15]);
  buf(\xm8051_golden_model_1.n1250 [48], input_sha_func_21[16]);
  buf(\xm8051_golden_model_1.n1250 [49], input_sha_func_21[17]);
  buf(\xm8051_golden_model_1.n1250 [50], input_sha_func_21[18]);
  buf(\xm8051_golden_model_1.n1250 [51], input_sha_func_21[19]);
  buf(\xm8051_golden_model_1.n1250 [52], input_sha_func_21[20]);
  buf(\xm8051_golden_model_1.n1250 [53], input_sha_func_21[21]);
  buf(\xm8051_golden_model_1.n1250 [54], input_sha_func_21[22]);
  buf(\xm8051_golden_model_1.n1250 [55], input_sha_func_21[23]);
  buf(\xm8051_golden_model_1.n1250 [56], input_sha_func_21[24]);
  buf(\xm8051_golden_model_1.n1250 [57], input_sha_func_21[25]);
  buf(\xm8051_golden_model_1.n1250 [58], input_sha_func_21[26]);
  buf(\xm8051_golden_model_1.n1250 [59], input_sha_func_21[27]);
  buf(\xm8051_golden_model_1.n1250 [60], input_sha_func_21[28]);
  buf(\xm8051_golden_model_1.n1250 [61], input_sha_func_21[29]);
  buf(\xm8051_golden_model_1.n1250 [62], input_sha_func_21[30]);
  buf(\xm8051_golden_model_1.n1250 [63], input_sha_func_21[31]);
  buf(\xm8051_golden_model_1.n1250 [64], input_sha_func_21[32]);
  buf(\xm8051_golden_model_1.n1250 [65], input_sha_func_21[33]);
  buf(\xm8051_golden_model_1.n1250 [66], input_sha_func_21[34]);
  buf(\xm8051_golden_model_1.n1250 [67], input_sha_func_21[35]);
  buf(\xm8051_golden_model_1.n1250 [68], input_sha_func_21[36]);
  buf(\xm8051_golden_model_1.n1250 [69], input_sha_func_21[37]);
  buf(\xm8051_golden_model_1.n1250 [70], input_sha_func_21[38]);
  buf(\xm8051_golden_model_1.n1250 [71], input_sha_func_21[39]);
  buf(\xm8051_golden_model_1.n1250 [72], input_sha_func_21[40]);
  buf(\xm8051_golden_model_1.n1250 [73], input_sha_func_21[41]);
  buf(\xm8051_golden_model_1.n1250 [74], input_sha_func_21[42]);
  buf(\xm8051_golden_model_1.n1250 [75], input_sha_func_21[43]);
  buf(\xm8051_golden_model_1.n1250 [76], input_sha_func_21[44]);
  buf(\xm8051_golden_model_1.n1250 [77], input_sha_func_21[45]);
  buf(\xm8051_golden_model_1.n1250 [78], input_sha_func_21[46]);
  buf(\xm8051_golden_model_1.n1250 [79], input_sha_func_21[47]);
  buf(\xm8051_golden_model_1.n1250 [80], input_sha_func_21[48]);
  buf(\xm8051_golden_model_1.n1250 [81], input_sha_func_21[49]);
  buf(\xm8051_golden_model_1.n1250 [82], input_sha_func_21[50]);
  buf(\xm8051_golden_model_1.n1250 [83], input_sha_func_21[51]);
  buf(\xm8051_golden_model_1.n1250 [84], input_sha_func_21[52]);
  buf(\xm8051_golden_model_1.n1250 [85], input_sha_func_21[53]);
  buf(\xm8051_golden_model_1.n1250 [86], input_sha_func_21[54]);
  buf(\xm8051_golden_model_1.n1250 [87], input_sha_func_21[55]);
  buf(\xm8051_golden_model_1.n1250 [88], input_sha_func_21[56]);
  buf(\xm8051_golden_model_1.n1250 [89], input_sha_func_21[57]);
  buf(\xm8051_golden_model_1.n1250 [90], input_sha_func_21[58]);
  buf(\xm8051_golden_model_1.n1250 [91], input_sha_func_21[59]);
  buf(\xm8051_golden_model_1.n1250 [92], input_sha_func_21[60]);
  buf(\xm8051_golden_model_1.n1250 [93], input_sha_func_21[61]);
  buf(\xm8051_golden_model_1.n1250 [94], input_sha_func_21[62]);
  buf(\xm8051_golden_model_1.n1250 [95], input_sha_func_21[63]);
  buf(\xm8051_golden_model_1.n1250 [96], input_sha_func_20[0]);
  buf(\xm8051_golden_model_1.n1250 [97], input_sha_func_20[1]);
  buf(\xm8051_golden_model_1.n1250 [98], input_sha_func_20[2]);
  buf(\xm8051_golden_model_1.n1250 [99], input_sha_func_20[3]);
  buf(\xm8051_golden_model_1.n1250 [100], input_sha_func_20[4]);
  buf(\xm8051_golden_model_1.n1250 [101], input_sha_func_20[5]);
  buf(\xm8051_golden_model_1.n1250 [102], input_sha_func_20[6]);
  buf(\xm8051_golden_model_1.n1250 [103], input_sha_func_20[7]);
  buf(\xm8051_golden_model_1.n1250 [104], input_sha_func_20[8]);
  buf(\xm8051_golden_model_1.n1250 [105], input_sha_func_20[9]);
  buf(\xm8051_golden_model_1.n1250 [106], input_sha_func_20[10]);
  buf(\xm8051_golden_model_1.n1250 [107], input_sha_func_20[11]);
  buf(\xm8051_golden_model_1.n1250 [108], input_sha_func_20[12]);
  buf(\xm8051_golden_model_1.n1250 [109], input_sha_func_20[13]);
  buf(\xm8051_golden_model_1.n1250 [110], input_sha_func_20[14]);
  buf(\xm8051_golden_model_1.n1250 [111], input_sha_func_20[15]);
  buf(\xm8051_golden_model_1.n1250 [112], input_sha_func_20[16]);
  buf(\xm8051_golden_model_1.n1250 [113], input_sha_func_20[17]);
  buf(\xm8051_golden_model_1.n1250 [114], input_sha_func_20[18]);
  buf(\xm8051_golden_model_1.n1250 [115], input_sha_func_20[19]);
  buf(\xm8051_golden_model_1.n1250 [116], input_sha_func_20[20]);
  buf(\xm8051_golden_model_1.n1250 [117], input_sha_func_20[21]);
  buf(\xm8051_golden_model_1.n1250 [118], input_sha_func_20[22]);
  buf(\xm8051_golden_model_1.n1250 [119], input_sha_func_20[23]);
  buf(\xm8051_golden_model_1.n1250 [120], input_sha_func_20[24]);
  buf(\xm8051_golden_model_1.n1250 [121], input_sha_func_20[25]);
  buf(\xm8051_golden_model_1.n1250 [122], input_sha_func_20[26]);
  buf(\xm8051_golden_model_1.n1250 [123], input_sha_func_20[27]);
  buf(\xm8051_golden_model_1.n1250 [124], input_sha_func_20[28]);
  buf(\xm8051_golden_model_1.n1250 [125], input_sha_func_20[29]);
  buf(\xm8051_golden_model_1.n1250 [126], input_sha_func_20[30]);
  buf(\xm8051_golden_model_1.n1250 [127], input_sha_func_20[31]);
  buf(\xm8051_golden_model_1.n1250 [128], input_sha_func_20[32]);
  buf(\xm8051_golden_model_1.n1250 [129], input_sha_func_20[33]);
  buf(\xm8051_golden_model_1.n1250 [130], input_sha_func_20[34]);
  buf(\xm8051_golden_model_1.n1250 [131], input_sha_func_20[35]);
  buf(\xm8051_golden_model_1.n1250 [132], input_sha_func_20[36]);
  buf(\xm8051_golden_model_1.n1250 [133], input_sha_func_20[37]);
  buf(\xm8051_golden_model_1.n1250 [134], input_sha_func_20[38]);
  buf(\xm8051_golden_model_1.n1250 [135], input_sha_func_20[39]);
  buf(\xm8051_golden_model_1.n1250 [136], input_sha_func_20[40]);
  buf(\xm8051_golden_model_1.n1250 [137], input_sha_func_20[41]);
  buf(\xm8051_golden_model_1.n1250 [138], input_sha_func_20[42]);
  buf(\xm8051_golden_model_1.n1250 [139], input_sha_func_20[43]);
  buf(\xm8051_golden_model_1.n1250 [140], input_sha_func_20[44]);
  buf(\xm8051_golden_model_1.n1250 [141], input_sha_func_20[45]);
  buf(\xm8051_golden_model_1.n1250 [142], input_sha_func_20[46]);
  buf(\xm8051_golden_model_1.n1250 [143], input_sha_func_20[47]);
  buf(\xm8051_golden_model_1.n1250 [144], input_sha_func_20[48]);
  buf(\xm8051_golden_model_1.n1250 [145], input_sha_func_20[49]);
  buf(\xm8051_golden_model_1.n1250 [146], input_sha_func_20[50]);
  buf(\xm8051_golden_model_1.n1250 [147], input_sha_func_20[51]);
  buf(\xm8051_golden_model_1.n1250 [148], input_sha_func_20[52]);
  buf(\xm8051_golden_model_1.n1250 [149], input_sha_func_20[53]);
  buf(\xm8051_golden_model_1.n1250 [150], input_sha_func_20[54]);
  buf(\xm8051_golden_model_1.n1250 [151], input_sha_func_20[55]);
  buf(\xm8051_golden_model_1.n1250 [152], input_sha_func_20[56]);
  buf(\xm8051_golden_model_1.n1250 [153], input_sha_func_20[57]);
  buf(\xm8051_golden_model_1.n1250 [154], input_sha_func_20[58]);
  buf(\xm8051_golden_model_1.n1250 [155], input_sha_func_20[59]);
  buf(\xm8051_golden_model_1.n1250 [156], input_sha_func_20[60]);
  buf(\xm8051_golden_model_1.n1250 [157], input_sha_func_20[61]);
  buf(\xm8051_golden_model_1.n1250 [158], input_sha_func_20[62]);
  buf(\xm8051_golden_model_1.n1250 [159], input_sha_func_20[63]);
  buf(\xm8051_golden_model_1.n1248 [0], RD_xram_80[0]);
  buf(\xm8051_golden_model_1.n1248 [1], RD_xram_80[1]);
  buf(\xm8051_golden_model_1.n1248 [2], RD_xram_80[2]);
  buf(\xm8051_golden_model_1.n1248 [3], RD_xram_80[3]);
  buf(\xm8051_golden_model_1.n1248 [4], RD_xram_80[4]);
  buf(\xm8051_golden_model_1.n1248 [5], RD_xram_80[5]);
  buf(\xm8051_golden_model_1.n1248 [6], RD_xram_80[6]);
  buf(\xm8051_golden_model_1.n1248 [7], RD_xram_80[7]);
  buf(\xm8051_golden_model_1.n1248 [8], RD_xram_79[0]);
  buf(\xm8051_golden_model_1.n1248 [9], RD_xram_79[1]);
  buf(\xm8051_golden_model_1.n1248 [10], RD_xram_79[2]);
  buf(\xm8051_golden_model_1.n1248 [11], RD_xram_79[3]);
  buf(\xm8051_golden_model_1.n1248 [12], RD_xram_79[4]);
  buf(\xm8051_golden_model_1.n1248 [13], RD_xram_79[5]);
  buf(\xm8051_golden_model_1.n1248 [14], RD_xram_79[6]);
  buf(\xm8051_golden_model_1.n1248 [15], RD_xram_79[7]);
  buf(\xm8051_golden_model_1.n1248 [16], RD_xram_78[0]);
  buf(\xm8051_golden_model_1.n1248 [17], RD_xram_78[1]);
  buf(\xm8051_golden_model_1.n1248 [18], RD_xram_78[2]);
  buf(\xm8051_golden_model_1.n1248 [19], RD_xram_78[3]);
  buf(\xm8051_golden_model_1.n1248 [20], RD_xram_78[4]);
  buf(\xm8051_golden_model_1.n1248 [21], RD_xram_78[5]);
  buf(\xm8051_golden_model_1.n1248 [22], RD_xram_78[6]);
  buf(\xm8051_golden_model_1.n1248 [23], RD_xram_78[7]);
  buf(\xm8051_golden_model_1.n1248 [24], RD_xram_77[0]);
  buf(\xm8051_golden_model_1.n1248 [25], RD_xram_77[1]);
  buf(\xm8051_golden_model_1.n1248 [26], RD_xram_77[2]);
  buf(\xm8051_golden_model_1.n1248 [27], RD_xram_77[3]);
  buf(\xm8051_golden_model_1.n1248 [28], RD_xram_77[4]);
  buf(\xm8051_golden_model_1.n1248 [29], RD_xram_77[5]);
  buf(\xm8051_golden_model_1.n1248 [30], RD_xram_77[6]);
  buf(\xm8051_golden_model_1.n1248 [31], RD_xram_77[7]);
  buf(\xm8051_golden_model_1.n1248 [32], RD_xram_76[0]);
  buf(\xm8051_golden_model_1.n1248 [33], RD_xram_76[1]);
  buf(\xm8051_golden_model_1.n1248 [34], RD_xram_76[2]);
  buf(\xm8051_golden_model_1.n1248 [35], RD_xram_76[3]);
  buf(\xm8051_golden_model_1.n1248 [36], RD_xram_76[4]);
  buf(\xm8051_golden_model_1.n1248 [37], RD_xram_76[5]);
  buf(\xm8051_golden_model_1.n1248 [38], RD_xram_76[6]);
  buf(\xm8051_golden_model_1.n1248 [39], RD_xram_76[7]);
  buf(\xm8051_golden_model_1.n1248 [40], RD_xram_75[0]);
  buf(\xm8051_golden_model_1.n1248 [41], RD_xram_75[1]);
  buf(\xm8051_golden_model_1.n1248 [42], RD_xram_75[2]);
  buf(\xm8051_golden_model_1.n1248 [43], RD_xram_75[3]);
  buf(\xm8051_golden_model_1.n1248 [44], RD_xram_75[4]);
  buf(\xm8051_golden_model_1.n1248 [45], RD_xram_75[5]);
  buf(\xm8051_golden_model_1.n1248 [46], RD_xram_75[6]);
  buf(\xm8051_golden_model_1.n1248 [47], RD_xram_75[7]);
  buf(\xm8051_golden_model_1.n1248 [48], RD_xram_74[0]);
  buf(\xm8051_golden_model_1.n1248 [49], RD_xram_74[1]);
  buf(\xm8051_golden_model_1.n1248 [50], RD_xram_74[2]);
  buf(\xm8051_golden_model_1.n1248 [51], RD_xram_74[3]);
  buf(\xm8051_golden_model_1.n1248 [52], RD_xram_74[4]);
  buf(\xm8051_golden_model_1.n1248 [53], RD_xram_74[5]);
  buf(\xm8051_golden_model_1.n1248 [54], RD_xram_74[6]);
  buf(\xm8051_golden_model_1.n1248 [55], RD_xram_74[7]);
  buf(\xm8051_golden_model_1.n1248 [56], RD_xram_73[0]);
  buf(\xm8051_golden_model_1.n1248 [57], RD_xram_73[1]);
  buf(\xm8051_golden_model_1.n1248 [58], RD_xram_73[2]);
  buf(\xm8051_golden_model_1.n1248 [59], RD_xram_73[3]);
  buf(\xm8051_golden_model_1.n1248 [60], RD_xram_73[4]);
  buf(\xm8051_golden_model_1.n1248 [61], RD_xram_73[5]);
  buf(\xm8051_golden_model_1.n1248 [62], RD_xram_73[6]);
  buf(\xm8051_golden_model_1.n1248 [63], RD_xram_73[7]);
  buf(\xm8051_golden_model_1.n1248 [64], RD_xram_72[0]);
  buf(\xm8051_golden_model_1.n1248 [65], RD_xram_72[1]);
  buf(\xm8051_golden_model_1.n1248 [66], RD_xram_72[2]);
  buf(\xm8051_golden_model_1.n1248 [67], RD_xram_72[3]);
  buf(\xm8051_golden_model_1.n1248 [68], RD_xram_72[4]);
  buf(\xm8051_golden_model_1.n1248 [69], RD_xram_72[5]);
  buf(\xm8051_golden_model_1.n1248 [70], RD_xram_72[6]);
  buf(\xm8051_golden_model_1.n1248 [71], RD_xram_72[7]);
  buf(\xm8051_golden_model_1.n1248 [72], RD_xram_71[0]);
  buf(\xm8051_golden_model_1.n1248 [73], RD_xram_71[1]);
  buf(\xm8051_golden_model_1.n1248 [74], RD_xram_71[2]);
  buf(\xm8051_golden_model_1.n1248 [75], RD_xram_71[3]);
  buf(\xm8051_golden_model_1.n1248 [76], RD_xram_71[4]);
  buf(\xm8051_golden_model_1.n1248 [77], RD_xram_71[5]);
  buf(\xm8051_golden_model_1.n1248 [78], RD_xram_71[6]);
  buf(\xm8051_golden_model_1.n1248 [79], RD_xram_71[7]);
  buf(\xm8051_golden_model_1.n1248 [80], RD_xram_70[0]);
  buf(\xm8051_golden_model_1.n1248 [81], RD_xram_70[1]);
  buf(\xm8051_golden_model_1.n1248 [82], RD_xram_70[2]);
  buf(\xm8051_golden_model_1.n1248 [83], RD_xram_70[3]);
  buf(\xm8051_golden_model_1.n1248 [84], RD_xram_70[4]);
  buf(\xm8051_golden_model_1.n1248 [85], RD_xram_70[5]);
  buf(\xm8051_golden_model_1.n1248 [86], RD_xram_70[6]);
  buf(\xm8051_golden_model_1.n1248 [87], RD_xram_70[7]);
  buf(\xm8051_golden_model_1.n1248 [88], RD_xram_69[0]);
  buf(\xm8051_golden_model_1.n1248 [89], RD_xram_69[1]);
  buf(\xm8051_golden_model_1.n1248 [90], RD_xram_69[2]);
  buf(\xm8051_golden_model_1.n1248 [91], RD_xram_69[3]);
  buf(\xm8051_golden_model_1.n1248 [92], RD_xram_69[4]);
  buf(\xm8051_golden_model_1.n1248 [93], RD_xram_69[5]);
  buf(\xm8051_golden_model_1.n1248 [94], RD_xram_69[6]);
  buf(\xm8051_golden_model_1.n1248 [95], RD_xram_69[7]);
  buf(\xm8051_golden_model_1.n1248 [96], RD_xram_68[0]);
  buf(\xm8051_golden_model_1.n1248 [97], RD_xram_68[1]);
  buf(\xm8051_golden_model_1.n1248 [98], RD_xram_68[2]);
  buf(\xm8051_golden_model_1.n1248 [99], RD_xram_68[3]);
  buf(\xm8051_golden_model_1.n1248 [100], RD_xram_68[4]);
  buf(\xm8051_golden_model_1.n1248 [101], RD_xram_68[5]);
  buf(\xm8051_golden_model_1.n1248 [102], RD_xram_68[6]);
  buf(\xm8051_golden_model_1.n1248 [103], RD_xram_68[7]);
  buf(\xm8051_golden_model_1.n1248 [104], RD_xram_67[0]);
  buf(\xm8051_golden_model_1.n1248 [105], RD_xram_67[1]);
  buf(\xm8051_golden_model_1.n1248 [106], RD_xram_67[2]);
  buf(\xm8051_golden_model_1.n1248 [107], RD_xram_67[3]);
  buf(\xm8051_golden_model_1.n1248 [108], RD_xram_67[4]);
  buf(\xm8051_golden_model_1.n1248 [109], RD_xram_67[5]);
  buf(\xm8051_golden_model_1.n1248 [110], RD_xram_67[6]);
  buf(\xm8051_golden_model_1.n1248 [111], RD_xram_67[7]);
  buf(\xm8051_golden_model_1.n1248 [112], RD_xram_66[0]);
  buf(\xm8051_golden_model_1.n1248 [113], RD_xram_66[1]);
  buf(\xm8051_golden_model_1.n1248 [114], RD_xram_66[2]);
  buf(\xm8051_golden_model_1.n1248 [115], RD_xram_66[3]);
  buf(\xm8051_golden_model_1.n1248 [116], RD_xram_66[4]);
  buf(\xm8051_golden_model_1.n1248 [117], RD_xram_66[5]);
  buf(\xm8051_golden_model_1.n1248 [118], RD_xram_66[6]);
  buf(\xm8051_golden_model_1.n1248 [119], RD_xram_66[7]);
  buf(\xm8051_golden_model_1.n1248 [120], RD_xram_65[0]);
  buf(\xm8051_golden_model_1.n1248 [121], RD_xram_65[1]);
  buf(\xm8051_golden_model_1.n1248 [122], RD_xram_65[2]);
  buf(\xm8051_golden_model_1.n1248 [123], RD_xram_65[3]);
  buf(\xm8051_golden_model_1.n1248 [124], RD_xram_65[4]);
  buf(\xm8051_golden_model_1.n1248 [125], RD_xram_65[5]);
  buf(\xm8051_golden_model_1.n1248 [126], RD_xram_65[6]);
  buf(\xm8051_golden_model_1.n1248 [127], RD_xram_65[7]);
  buf(\xm8051_golden_model_1.n1248 [128], RD_xram_64[0]);
  buf(\xm8051_golden_model_1.n1248 [129], RD_xram_64[1]);
  buf(\xm8051_golden_model_1.n1248 [130], RD_xram_64[2]);
  buf(\xm8051_golden_model_1.n1248 [131], RD_xram_64[3]);
  buf(\xm8051_golden_model_1.n1248 [132], RD_xram_64[4]);
  buf(\xm8051_golden_model_1.n1248 [133], RD_xram_64[5]);
  buf(\xm8051_golden_model_1.n1248 [134], RD_xram_64[6]);
  buf(\xm8051_golden_model_1.n1248 [135], RD_xram_64[7]);
  buf(\xm8051_golden_model_1.n1248 [136], RD_xram_63[0]);
  buf(\xm8051_golden_model_1.n1248 [137], RD_xram_63[1]);
  buf(\xm8051_golden_model_1.n1248 [138], RD_xram_63[2]);
  buf(\xm8051_golden_model_1.n1248 [139], RD_xram_63[3]);
  buf(\xm8051_golden_model_1.n1248 [140], RD_xram_63[4]);
  buf(\xm8051_golden_model_1.n1248 [141], RD_xram_63[5]);
  buf(\xm8051_golden_model_1.n1248 [142], RD_xram_63[6]);
  buf(\xm8051_golden_model_1.n1248 [143], RD_xram_63[7]);
  buf(\xm8051_golden_model_1.n1248 [144], RD_xram_62[0]);
  buf(\xm8051_golden_model_1.n1248 [145], RD_xram_62[1]);
  buf(\xm8051_golden_model_1.n1248 [146], RD_xram_62[2]);
  buf(\xm8051_golden_model_1.n1248 [147], RD_xram_62[3]);
  buf(\xm8051_golden_model_1.n1248 [148], RD_xram_62[4]);
  buf(\xm8051_golden_model_1.n1248 [149], RD_xram_62[5]);
  buf(\xm8051_golden_model_1.n1248 [150], RD_xram_62[6]);
  buf(\xm8051_golden_model_1.n1248 [151], RD_xram_62[7]);
  buf(\xm8051_golden_model_1.n1248 [152], RD_xram_61[0]);
  buf(\xm8051_golden_model_1.n1248 [153], RD_xram_61[1]);
  buf(\xm8051_golden_model_1.n1248 [154], RD_xram_61[2]);
  buf(\xm8051_golden_model_1.n1248 [155], RD_xram_61[3]);
  buf(\xm8051_golden_model_1.n1248 [156], RD_xram_61[4]);
  buf(\xm8051_golden_model_1.n1248 [157], RD_xram_61[5]);
  buf(\xm8051_golden_model_1.n1248 [158], RD_xram_61[6]);
  buf(\xm8051_golden_model_1.n1248 [159], RD_xram_61[7]);
  buf(\xm8051_golden_model_1.n1248 [160], RD_xram_60[0]);
  buf(\xm8051_golden_model_1.n1248 [161], RD_xram_60[1]);
  buf(\xm8051_golden_model_1.n1248 [162], RD_xram_60[2]);
  buf(\xm8051_golden_model_1.n1248 [163], RD_xram_60[3]);
  buf(\xm8051_golden_model_1.n1248 [164], RD_xram_60[4]);
  buf(\xm8051_golden_model_1.n1248 [165], RD_xram_60[5]);
  buf(\xm8051_golden_model_1.n1248 [166], RD_xram_60[6]);
  buf(\xm8051_golden_model_1.n1248 [167], RD_xram_60[7]);
  buf(\xm8051_golden_model_1.n1248 [168], RD_xram_59[0]);
  buf(\xm8051_golden_model_1.n1248 [169], RD_xram_59[1]);
  buf(\xm8051_golden_model_1.n1248 [170], RD_xram_59[2]);
  buf(\xm8051_golden_model_1.n1248 [171], RD_xram_59[3]);
  buf(\xm8051_golden_model_1.n1248 [172], RD_xram_59[4]);
  buf(\xm8051_golden_model_1.n1248 [173], RD_xram_59[5]);
  buf(\xm8051_golden_model_1.n1248 [174], RD_xram_59[6]);
  buf(\xm8051_golden_model_1.n1248 [175], RD_xram_59[7]);
  buf(\xm8051_golden_model_1.n1248 [176], RD_xram_58[0]);
  buf(\xm8051_golden_model_1.n1248 [177], RD_xram_58[1]);
  buf(\xm8051_golden_model_1.n1248 [178], RD_xram_58[2]);
  buf(\xm8051_golden_model_1.n1248 [179], RD_xram_58[3]);
  buf(\xm8051_golden_model_1.n1248 [180], RD_xram_58[4]);
  buf(\xm8051_golden_model_1.n1248 [181], RD_xram_58[5]);
  buf(\xm8051_golden_model_1.n1248 [182], RD_xram_58[6]);
  buf(\xm8051_golden_model_1.n1248 [183], RD_xram_58[7]);
  buf(\xm8051_golden_model_1.n1248 [184], RD_xram_57[0]);
  buf(\xm8051_golden_model_1.n1248 [185], RD_xram_57[1]);
  buf(\xm8051_golden_model_1.n1248 [186], RD_xram_57[2]);
  buf(\xm8051_golden_model_1.n1248 [187], RD_xram_57[3]);
  buf(\xm8051_golden_model_1.n1248 [188], RD_xram_57[4]);
  buf(\xm8051_golden_model_1.n1248 [189], RD_xram_57[5]);
  buf(\xm8051_golden_model_1.n1248 [190], RD_xram_57[6]);
  buf(\xm8051_golden_model_1.n1248 [191], RD_xram_57[7]);
  buf(\xm8051_golden_model_1.n1248 [192], RD_xram_56[0]);
  buf(\xm8051_golden_model_1.n1248 [193], RD_xram_56[1]);
  buf(\xm8051_golden_model_1.n1248 [194], RD_xram_56[2]);
  buf(\xm8051_golden_model_1.n1248 [195], RD_xram_56[3]);
  buf(\xm8051_golden_model_1.n1248 [196], RD_xram_56[4]);
  buf(\xm8051_golden_model_1.n1248 [197], RD_xram_56[5]);
  buf(\xm8051_golden_model_1.n1248 [198], RD_xram_56[6]);
  buf(\xm8051_golden_model_1.n1248 [199], RD_xram_56[7]);
  buf(\xm8051_golden_model_1.n1248 [200], RD_xram_55[0]);
  buf(\xm8051_golden_model_1.n1248 [201], RD_xram_55[1]);
  buf(\xm8051_golden_model_1.n1248 [202], RD_xram_55[2]);
  buf(\xm8051_golden_model_1.n1248 [203], RD_xram_55[3]);
  buf(\xm8051_golden_model_1.n1248 [204], RD_xram_55[4]);
  buf(\xm8051_golden_model_1.n1248 [205], RD_xram_55[5]);
  buf(\xm8051_golden_model_1.n1248 [206], RD_xram_55[6]);
  buf(\xm8051_golden_model_1.n1248 [207], RD_xram_55[7]);
  buf(\xm8051_golden_model_1.n1248 [208], RD_xram_54[0]);
  buf(\xm8051_golden_model_1.n1248 [209], RD_xram_54[1]);
  buf(\xm8051_golden_model_1.n1248 [210], RD_xram_54[2]);
  buf(\xm8051_golden_model_1.n1248 [211], RD_xram_54[3]);
  buf(\xm8051_golden_model_1.n1248 [212], RD_xram_54[4]);
  buf(\xm8051_golden_model_1.n1248 [213], RD_xram_54[5]);
  buf(\xm8051_golden_model_1.n1248 [214], RD_xram_54[6]);
  buf(\xm8051_golden_model_1.n1248 [215], RD_xram_54[7]);
  buf(\xm8051_golden_model_1.n1248 [216], RD_xram_53[0]);
  buf(\xm8051_golden_model_1.n1248 [217], RD_xram_53[1]);
  buf(\xm8051_golden_model_1.n1248 [218], RD_xram_53[2]);
  buf(\xm8051_golden_model_1.n1248 [219], RD_xram_53[3]);
  buf(\xm8051_golden_model_1.n1248 [220], RD_xram_53[4]);
  buf(\xm8051_golden_model_1.n1248 [221], RD_xram_53[5]);
  buf(\xm8051_golden_model_1.n1248 [222], RD_xram_53[6]);
  buf(\xm8051_golden_model_1.n1248 [223], RD_xram_53[7]);
  buf(\xm8051_golden_model_1.n1248 [224], RD_xram_52[0]);
  buf(\xm8051_golden_model_1.n1248 [225], RD_xram_52[1]);
  buf(\xm8051_golden_model_1.n1248 [226], RD_xram_52[2]);
  buf(\xm8051_golden_model_1.n1248 [227], RD_xram_52[3]);
  buf(\xm8051_golden_model_1.n1248 [228], RD_xram_52[4]);
  buf(\xm8051_golden_model_1.n1248 [229], RD_xram_52[5]);
  buf(\xm8051_golden_model_1.n1248 [230], RD_xram_52[6]);
  buf(\xm8051_golden_model_1.n1248 [231], RD_xram_52[7]);
  buf(\xm8051_golden_model_1.n1248 [232], RD_xram_51[0]);
  buf(\xm8051_golden_model_1.n1248 [233], RD_xram_51[1]);
  buf(\xm8051_golden_model_1.n1248 [234], RD_xram_51[2]);
  buf(\xm8051_golden_model_1.n1248 [235], RD_xram_51[3]);
  buf(\xm8051_golden_model_1.n1248 [236], RD_xram_51[4]);
  buf(\xm8051_golden_model_1.n1248 [237], RD_xram_51[5]);
  buf(\xm8051_golden_model_1.n1248 [238], RD_xram_51[6]);
  buf(\xm8051_golden_model_1.n1248 [239], RD_xram_51[7]);
  buf(\xm8051_golden_model_1.n1248 [240], RD_xram_50[0]);
  buf(\xm8051_golden_model_1.n1248 [241], RD_xram_50[1]);
  buf(\xm8051_golden_model_1.n1248 [242], RD_xram_50[2]);
  buf(\xm8051_golden_model_1.n1248 [243], RD_xram_50[3]);
  buf(\xm8051_golden_model_1.n1248 [244], RD_xram_50[4]);
  buf(\xm8051_golden_model_1.n1248 [245], RD_xram_50[5]);
  buf(\xm8051_golden_model_1.n1248 [246], RD_xram_50[6]);
  buf(\xm8051_golden_model_1.n1248 [247], RD_xram_50[7]);
  buf(\xm8051_golden_model_1.n1248 [248], RD_xram_49[0]);
  buf(\xm8051_golden_model_1.n1248 [249], RD_xram_49[1]);
  buf(\xm8051_golden_model_1.n1248 [250], RD_xram_49[2]);
  buf(\xm8051_golden_model_1.n1248 [251], RD_xram_49[3]);
  buf(\xm8051_golden_model_1.n1248 [252], RD_xram_49[4]);
  buf(\xm8051_golden_model_1.n1248 [253], RD_xram_49[5]);
  buf(\xm8051_golden_model_1.n1248 [254], RD_xram_49[6]);
  buf(\xm8051_golden_model_1.n1248 [255], RD_xram_49[7]);
  buf(\xm8051_golden_model_1.n1248 [256], RD_xram_48[0]);
  buf(\xm8051_golden_model_1.n1248 [257], RD_xram_48[1]);
  buf(\xm8051_golden_model_1.n1248 [258], RD_xram_48[2]);
  buf(\xm8051_golden_model_1.n1248 [259], RD_xram_48[3]);
  buf(\xm8051_golden_model_1.n1248 [260], RD_xram_48[4]);
  buf(\xm8051_golden_model_1.n1248 [261], RD_xram_48[5]);
  buf(\xm8051_golden_model_1.n1248 [262], RD_xram_48[6]);
  buf(\xm8051_golden_model_1.n1248 [263], RD_xram_48[7]);
  buf(\xm8051_golden_model_1.n1248 [264], RD_xram_47[0]);
  buf(\xm8051_golden_model_1.n1248 [265], RD_xram_47[1]);
  buf(\xm8051_golden_model_1.n1248 [266], RD_xram_47[2]);
  buf(\xm8051_golden_model_1.n1248 [267], RD_xram_47[3]);
  buf(\xm8051_golden_model_1.n1248 [268], RD_xram_47[4]);
  buf(\xm8051_golden_model_1.n1248 [269], RD_xram_47[5]);
  buf(\xm8051_golden_model_1.n1248 [270], RD_xram_47[6]);
  buf(\xm8051_golden_model_1.n1248 [271], RD_xram_47[7]);
  buf(\xm8051_golden_model_1.n1248 [272], RD_xram_46[0]);
  buf(\xm8051_golden_model_1.n1248 [273], RD_xram_46[1]);
  buf(\xm8051_golden_model_1.n1248 [274], RD_xram_46[2]);
  buf(\xm8051_golden_model_1.n1248 [275], RD_xram_46[3]);
  buf(\xm8051_golden_model_1.n1248 [276], RD_xram_46[4]);
  buf(\xm8051_golden_model_1.n1248 [277], RD_xram_46[5]);
  buf(\xm8051_golden_model_1.n1248 [278], RD_xram_46[6]);
  buf(\xm8051_golden_model_1.n1248 [279], RD_xram_46[7]);
  buf(\xm8051_golden_model_1.n1248 [280], RD_xram_45[0]);
  buf(\xm8051_golden_model_1.n1248 [281], RD_xram_45[1]);
  buf(\xm8051_golden_model_1.n1248 [282], RD_xram_45[2]);
  buf(\xm8051_golden_model_1.n1248 [283], RD_xram_45[3]);
  buf(\xm8051_golden_model_1.n1248 [284], RD_xram_45[4]);
  buf(\xm8051_golden_model_1.n1248 [285], RD_xram_45[5]);
  buf(\xm8051_golden_model_1.n1248 [286], RD_xram_45[6]);
  buf(\xm8051_golden_model_1.n1248 [287], RD_xram_45[7]);
  buf(\xm8051_golden_model_1.n1248 [288], RD_xram_44[0]);
  buf(\xm8051_golden_model_1.n1248 [289], RD_xram_44[1]);
  buf(\xm8051_golden_model_1.n1248 [290], RD_xram_44[2]);
  buf(\xm8051_golden_model_1.n1248 [291], RD_xram_44[3]);
  buf(\xm8051_golden_model_1.n1248 [292], RD_xram_44[4]);
  buf(\xm8051_golden_model_1.n1248 [293], RD_xram_44[5]);
  buf(\xm8051_golden_model_1.n1248 [294], RD_xram_44[6]);
  buf(\xm8051_golden_model_1.n1248 [295], RD_xram_44[7]);
  buf(\xm8051_golden_model_1.n1248 [296], RD_xram_43[0]);
  buf(\xm8051_golden_model_1.n1248 [297], RD_xram_43[1]);
  buf(\xm8051_golden_model_1.n1248 [298], RD_xram_43[2]);
  buf(\xm8051_golden_model_1.n1248 [299], RD_xram_43[3]);
  buf(\xm8051_golden_model_1.n1248 [300], RD_xram_43[4]);
  buf(\xm8051_golden_model_1.n1248 [301], RD_xram_43[5]);
  buf(\xm8051_golden_model_1.n1248 [302], RD_xram_43[6]);
  buf(\xm8051_golden_model_1.n1248 [303], RD_xram_43[7]);
  buf(\xm8051_golden_model_1.n1248 [304], RD_xram_42[0]);
  buf(\xm8051_golden_model_1.n1248 [305], RD_xram_42[1]);
  buf(\xm8051_golden_model_1.n1248 [306], RD_xram_42[2]);
  buf(\xm8051_golden_model_1.n1248 [307], RD_xram_42[3]);
  buf(\xm8051_golden_model_1.n1248 [308], RD_xram_42[4]);
  buf(\xm8051_golden_model_1.n1248 [309], RD_xram_42[5]);
  buf(\xm8051_golden_model_1.n1248 [310], RD_xram_42[6]);
  buf(\xm8051_golden_model_1.n1248 [311], RD_xram_42[7]);
  buf(\xm8051_golden_model_1.n1248 [312], RD_xram_41[0]);
  buf(\xm8051_golden_model_1.n1248 [313], RD_xram_41[1]);
  buf(\xm8051_golden_model_1.n1248 [314], RD_xram_41[2]);
  buf(\xm8051_golden_model_1.n1248 [315], RD_xram_41[3]);
  buf(\xm8051_golden_model_1.n1248 [316], RD_xram_41[4]);
  buf(\xm8051_golden_model_1.n1248 [317], RD_xram_41[5]);
  buf(\xm8051_golden_model_1.n1248 [318], RD_xram_41[6]);
  buf(\xm8051_golden_model_1.n1248 [319], RD_xram_41[7]);
  buf(\xm8051_golden_model_1.n1248 [320], RD_xram_40[0]);
  buf(\xm8051_golden_model_1.n1248 [321], RD_xram_40[1]);
  buf(\xm8051_golden_model_1.n1248 [322], RD_xram_40[2]);
  buf(\xm8051_golden_model_1.n1248 [323], RD_xram_40[3]);
  buf(\xm8051_golden_model_1.n1248 [324], RD_xram_40[4]);
  buf(\xm8051_golden_model_1.n1248 [325], RD_xram_40[5]);
  buf(\xm8051_golden_model_1.n1248 [326], RD_xram_40[6]);
  buf(\xm8051_golden_model_1.n1248 [327], RD_xram_40[7]);
  buf(\xm8051_golden_model_1.n1248 [328], RD_xram_39[0]);
  buf(\xm8051_golden_model_1.n1248 [329], RD_xram_39[1]);
  buf(\xm8051_golden_model_1.n1248 [330], RD_xram_39[2]);
  buf(\xm8051_golden_model_1.n1248 [331], RD_xram_39[3]);
  buf(\xm8051_golden_model_1.n1248 [332], RD_xram_39[4]);
  buf(\xm8051_golden_model_1.n1248 [333], RD_xram_39[5]);
  buf(\xm8051_golden_model_1.n1248 [334], RD_xram_39[6]);
  buf(\xm8051_golden_model_1.n1248 [335], RD_xram_39[7]);
  buf(\xm8051_golden_model_1.n1248 [336], RD_xram_38[0]);
  buf(\xm8051_golden_model_1.n1248 [337], RD_xram_38[1]);
  buf(\xm8051_golden_model_1.n1248 [338], RD_xram_38[2]);
  buf(\xm8051_golden_model_1.n1248 [339], RD_xram_38[3]);
  buf(\xm8051_golden_model_1.n1248 [340], RD_xram_38[4]);
  buf(\xm8051_golden_model_1.n1248 [341], RD_xram_38[5]);
  buf(\xm8051_golden_model_1.n1248 [342], RD_xram_38[6]);
  buf(\xm8051_golden_model_1.n1248 [343], RD_xram_38[7]);
  buf(\xm8051_golden_model_1.n1248 [344], RD_xram_37[0]);
  buf(\xm8051_golden_model_1.n1248 [345], RD_xram_37[1]);
  buf(\xm8051_golden_model_1.n1248 [346], RD_xram_37[2]);
  buf(\xm8051_golden_model_1.n1248 [347], RD_xram_37[3]);
  buf(\xm8051_golden_model_1.n1248 [348], RD_xram_37[4]);
  buf(\xm8051_golden_model_1.n1248 [349], RD_xram_37[5]);
  buf(\xm8051_golden_model_1.n1248 [350], RD_xram_37[6]);
  buf(\xm8051_golden_model_1.n1248 [351], RD_xram_37[7]);
  buf(\xm8051_golden_model_1.n1248 [352], RD_xram_36[0]);
  buf(\xm8051_golden_model_1.n1248 [353], RD_xram_36[1]);
  buf(\xm8051_golden_model_1.n1248 [354], RD_xram_36[2]);
  buf(\xm8051_golden_model_1.n1248 [355], RD_xram_36[3]);
  buf(\xm8051_golden_model_1.n1248 [356], RD_xram_36[4]);
  buf(\xm8051_golden_model_1.n1248 [357], RD_xram_36[5]);
  buf(\xm8051_golden_model_1.n1248 [358], RD_xram_36[6]);
  buf(\xm8051_golden_model_1.n1248 [359], RD_xram_36[7]);
  buf(\xm8051_golden_model_1.n1248 [360], RD_xram_35[0]);
  buf(\xm8051_golden_model_1.n1248 [361], RD_xram_35[1]);
  buf(\xm8051_golden_model_1.n1248 [362], RD_xram_35[2]);
  buf(\xm8051_golden_model_1.n1248 [363], RD_xram_35[3]);
  buf(\xm8051_golden_model_1.n1248 [364], RD_xram_35[4]);
  buf(\xm8051_golden_model_1.n1248 [365], RD_xram_35[5]);
  buf(\xm8051_golden_model_1.n1248 [366], RD_xram_35[6]);
  buf(\xm8051_golden_model_1.n1248 [367], RD_xram_35[7]);
  buf(\xm8051_golden_model_1.n1248 [368], RD_xram_34[0]);
  buf(\xm8051_golden_model_1.n1248 [369], RD_xram_34[1]);
  buf(\xm8051_golden_model_1.n1248 [370], RD_xram_34[2]);
  buf(\xm8051_golden_model_1.n1248 [371], RD_xram_34[3]);
  buf(\xm8051_golden_model_1.n1248 [372], RD_xram_34[4]);
  buf(\xm8051_golden_model_1.n1248 [373], RD_xram_34[5]);
  buf(\xm8051_golden_model_1.n1248 [374], RD_xram_34[6]);
  buf(\xm8051_golden_model_1.n1248 [375], RD_xram_34[7]);
  buf(\xm8051_golden_model_1.n1248 [376], RD_xram_33[0]);
  buf(\xm8051_golden_model_1.n1248 [377], RD_xram_33[1]);
  buf(\xm8051_golden_model_1.n1248 [378], RD_xram_33[2]);
  buf(\xm8051_golden_model_1.n1248 [379], RD_xram_33[3]);
  buf(\xm8051_golden_model_1.n1248 [380], RD_xram_33[4]);
  buf(\xm8051_golden_model_1.n1248 [381], RD_xram_33[5]);
  buf(\xm8051_golden_model_1.n1248 [382], RD_xram_33[6]);
  buf(\xm8051_golden_model_1.n1248 [383], RD_xram_33[7]);
  buf(\xm8051_golden_model_1.n1248 [384], RD_xram_32[0]);
  buf(\xm8051_golden_model_1.n1248 [385], RD_xram_32[1]);
  buf(\xm8051_golden_model_1.n1248 [386], RD_xram_32[2]);
  buf(\xm8051_golden_model_1.n1248 [387], RD_xram_32[3]);
  buf(\xm8051_golden_model_1.n1248 [388], RD_xram_32[4]);
  buf(\xm8051_golden_model_1.n1248 [389], RD_xram_32[5]);
  buf(\xm8051_golden_model_1.n1248 [390], RD_xram_32[6]);
  buf(\xm8051_golden_model_1.n1248 [391], RD_xram_32[7]);
  buf(\xm8051_golden_model_1.n1248 [392], RD_xram_31[0]);
  buf(\xm8051_golden_model_1.n1248 [393], RD_xram_31[1]);
  buf(\xm8051_golden_model_1.n1248 [394], RD_xram_31[2]);
  buf(\xm8051_golden_model_1.n1248 [395], RD_xram_31[3]);
  buf(\xm8051_golden_model_1.n1248 [396], RD_xram_31[4]);
  buf(\xm8051_golden_model_1.n1248 [397], RD_xram_31[5]);
  buf(\xm8051_golden_model_1.n1248 [398], RD_xram_31[6]);
  buf(\xm8051_golden_model_1.n1248 [399], RD_xram_31[7]);
  buf(\xm8051_golden_model_1.n1248 [400], RD_xram_30[0]);
  buf(\xm8051_golden_model_1.n1248 [401], RD_xram_30[1]);
  buf(\xm8051_golden_model_1.n1248 [402], RD_xram_30[2]);
  buf(\xm8051_golden_model_1.n1248 [403], RD_xram_30[3]);
  buf(\xm8051_golden_model_1.n1248 [404], RD_xram_30[4]);
  buf(\xm8051_golden_model_1.n1248 [405], RD_xram_30[5]);
  buf(\xm8051_golden_model_1.n1248 [406], RD_xram_30[6]);
  buf(\xm8051_golden_model_1.n1248 [407], RD_xram_30[7]);
  buf(\xm8051_golden_model_1.n1248 [408], RD_xram_29[0]);
  buf(\xm8051_golden_model_1.n1248 [409], RD_xram_29[1]);
  buf(\xm8051_golden_model_1.n1248 [410], RD_xram_29[2]);
  buf(\xm8051_golden_model_1.n1248 [411], RD_xram_29[3]);
  buf(\xm8051_golden_model_1.n1248 [412], RD_xram_29[4]);
  buf(\xm8051_golden_model_1.n1248 [413], RD_xram_29[5]);
  buf(\xm8051_golden_model_1.n1248 [414], RD_xram_29[6]);
  buf(\xm8051_golden_model_1.n1248 [415], RD_xram_29[7]);
  buf(\xm8051_golden_model_1.n1248 [416], RD_xram_28[0]);
  buf(\xm8051_golden_model_1.n1248 [417], RD_xram_28[1]);
  buf(\xm8051_golden_model_1.n1248 [418], RD_xram_28[2]);
  buf(\xm8051_golden_model_1.n1248 [419], RD_xram_28[3]);
  buf(\xm8051_golden_model_1.n1248 [420], RD_xram_28[4]);
  buf(\xm8051_golden_model_1.n1248 [421], RD_xram_28[5]);
  buf(\xm8051_golden_model_1.n1248 [422], RD_xram_28[6]);
  buf(\xm8051_golden_model_1.n1248 [423], RD_xram_28[7]);
  buf(\xm8051_golden_model_1.n1248 [424], RD_xram_27[0]);
  buf(\xm8051_golden_model_1.n1248 [425], RD_xram_27[1]);
  buf(\xm8051_golden_model_1.n1248 [426], RD_xram_27[2]);
  buf(\xm8051_golden_model_1.n1248 [427], RD_xram_27[3]);
  buf(\xm8051_golden_model_1.n1248 [428], RD_xram_27[4]);
  buf(\xm8051_golden_model_1.n1248 [429], RD_xram_27[5]);
  buf(\xm8051_golden_model_1.n1248 [430], RD_xram_27[6]);
  buf(\xm8051_golden_model_1.n1248 [431], RD_xram_27[7]);
  buf(\xm8051_golden_model_1.n1248 [432], RD_xram_26[0]);
  buf(\xm8051_golden_model_1.n1248 [433], RD_xram_26[1]);
  buf(\xm8051_golden_model_1.n1248 [434], RD_xram_26[2]);
  buf(\xm8051_golden_model_1.n1248 [435], RD_xram_26[3]);
  buf(\xm8051_golden_model_1.n1248 [436], RD_xram_26[4]);
  buf(\xm8051_golden_model_1.n1248 [437], RD_xram_26[5]);
  buf(\xm8051_golden_model_1.n1248 [438], RD_xram_26[6]);
  buf(\xm8051_golden_model_1.n1248 [439], RD_xram_26[7]);
  buf(\xm8051_golden_model_1.n1248 [440], RD_xram_25[0]);
  buf(\xm8051_golden_model_1.n1248 [441], RD_xram_25[1]);
  buf(\xm8051_golden_model_1.n1248 [442], RD_xram_25[2]);
  buf(\xm8051_golden_model_1.n1248 [443], RD_xram_25[3]);
  buf(\xm8051_golden_model_1.n1248 [444], RD_xram_25[4]);
  buf(\xm8051_golden_model_1.n1248 [445], RD_xram_25[5]);
  buf(\xm8051_golden_model_1.n1248 [446], RD_xram_25[6]);
  buf(\xm8051_golden_model_1.n1248 [447], RD_xram_25[7]);
  buf(\xm8051_golden_model_1.n1248 [448], RD_xram_24[0]);
  buf(\xm8051_golden_model_1.n1248 [449], RD_xram_24[1]);
  buf(\xm8051_golden_model_1.n1248 [450], RD_xram_24[2]);
  buf(\xm8051_golden_model_1.n1248 [451], RD_xram_24[3]);
  buf(\xm8051_golden_model_1.n1248 [452], RD_xram_24[4]);
  buf(\xm8051_golden_model_1.n1248 [453], RD_xram_24[5]);
  buf(\xm8051_golden_model_1.n1248 [454], RD_xram_24[6]);
  buf(\xm8051_golden_model_1.n1248 [455], RD_xram_24[7]);
  buf(\xm8051_golden_model_1.n1248 [456], RD_xram_23[0]);
  buf(\xm8051_golden_model_1.n1248 [457], RD_xram_23[1]);
  buf(\xm8051_golden_model_1.n1248 [458], RD_xram_23[2]);
  buf(\xm8051_golden_model_1.n1248 [459], RD_xram_23[3]);
  buf(\xm8051_golden_model_1.n1248 [460], RD_xram_23[4]);
  buf(\xm8051_golden_model_1.n1248 [461], RD_xram_23[5]);
  buf(\xm8051_golden_model_1.n1248 [462], RD_xram_23[6]);
  buf(\xm8051_golden_model_1.n1248 [463], RD_xram_23[7]);
  buf(\xm8051_golden_model_1.n1248 [464], RD_xram_22[0]);
  buf(\xm8051_golden_model_1.n1248 [465], RD_xram_22[1]);
  buf(\xm8051_golden_model_1.n1248 [466], RD_xram_22[2]);
  buf(\xm8051_golden_model_1.n1248 [467], RD_xram_22[3]);
  buf(\xm8051_golden_model_1.n1248 [468], RD_xram_22[4]);
  buf(\xm8051_golden_model_1.n1248 [469], RD_xram_22[5]);
  buf(\xm8051_golden_model_1.n1248 [470], RD_xram_22[6]);
  buf(\xm8051_golden_model_1.n1248 [471], RD_xram_22[7]);
  buf(\xm8051_golden_model_1.n1248 [472], RD_xram_21[0]);
  buf(\xm8051_golden_model_1.n1248 [473], RD_xram_21[1]);
  buf(\xm8051_golden_model_1.n1248 [474], RD_xram_21[2]);
  buf(\xm8051_golden_model_1.n1248 [475], RD_xram_21[3]);
  buf(\xm8051_golden_model_1.n1248 [476], RD_xram_21[4]);
  buf(\xm8051_golden_model_1.n1248 [477], RD_xram_21[5]);
  buf(\xm8051_golden_model_1.n1248 [478], RD_xram_21[6]);
  buf(\xm8051_golden_model_1.n1248 [479], RD_xram_21[7]);
  buf(\xm8051_golden_model_1.n1248 [480], RD_xram_20[0]);
  buf(\xm8051_golden_model_1.n1248 [481], RD_xram_20[1]);
  buf(\xm8051_golden_model_1.n1248 [482], RD_xram_20[2]);
  buf(\xm8051_golden_model_1.n1248 [483], RD_xram_20[3]);
  buf(\xm8051_golden_model_1.n1248 [484], RD_xram_20[4]);
  buf(\xm8051_golden_model_1.n1248 [485], RD_xram_20[5]);
  buf(\xm8051_golden_model_1.n1248 [486], RD_xram_20[6]);
  buf(\xm8051_golden_model_1.n1248 [487], RD_xram_20[7]);
  buf(\xm8051_golden_model_1.n1248 [488], RD_xram_19[0]);
  buf(\xm8051_golden_model_1.n1248 [489], RD_xram_19[1]);
  buf(\xm8051_golden_model_1.n1248 [490], RD_xram_19[2]);
  buf(\xm8051_golden_model_1.n1248 [491], RD_xram_19[3]);
  buf(\xm8051_golden_model_1.n1248 [492], RD_xram_19[4]);
  buf(\xm8051_golden_model_1.n1248 [493], RD_xram_19[5]);
  buf(\xm8051_golden_model_1.n1248 [494], RD_xram_19[6]);
  buf(\xm8051_golden_model_1.n1248 [495], RD_xram_19[7]);
  buf(\xm8051_golden_model_1.n1248 [496], RD_xram_18[0]);
  buf(\xm8051_golden_model_1.n1248 [497], RD_xram_18[1]);
  buf(\xm8051_golden_model_1.n1248 [498], RD_xram_18[2]);
  buf(\xm8051_golden_model_1.n1248 [499], RD_xram_18[3]);
  buf(\xm8051_golden_model_1.n1248 [500], RD_xram_18[4]);
  buf(\xm8051_golden_model_1.n1248 [501], RD_xram_18[5]);
  buf(\xm8051_golden_model_1.n1248 [502], RD_xram_18[6]);
  buf(\xm8051_golden_model_1.n1248 [503], RD_xram_18[7]);
  buf(\xm8051_golden_model_1.n1248 [504], RD_xram_17[0]);
  buf(\xm8051_golden_model_1.n1248 [505], RD_xram_17[1]);
  buf(\xm8051_golden_model_1.n1248 [506], RD_xram_17[2]);
  buf(\xm8051_golden_model_1.n1248 [507], RD_xram_17[3]);
  buf(\xm8051_golden_model_1.n1248 [508], RD_xram_17[4]);
  buf(\xm8051_golden_model_1.n1248 [509], RD_xram_17[5]);
  buf(\xm8051_golden_model_1.n1248 [510], RD_xram_17[6]);
  buf(\xm8051_golden_model_1.n1248 [511], RD_xram_17[7]);
  buf(\xm8051_golden_model_1.n0209 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0209 [1], \xm8051_golden_model_1.aes_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0209 [2], \xm8051_golden_model_1.aes_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n0209 [3], \xm8051_golden_model_1.aes_bytes_processed [3]);
  buf(\xm8051_golden_model_1.n0209 [4], \xm8051_golden_model_1.aes_bytes_processed [4]);
  buf(\xm8051_golden_model_1.n0209 [5], \xm8051_golden_model_1.aes_bytes_processed [5]);
  buf(\xm8051_golden_model_1.n0209 [6], \xm8051_golden_model_1.aes_bytes_processed [6]);
  buf(\xm8051_golden_model_1.n0209 [7], \xm8051_golden_model_1.aes_bytes_processed [7]);
  buf(\xm8051_golden_model_1.n0209 [8], \xm8051_golden_model_1.aes_bytes_processed [8]);
  buf(\xm8051_golden_model_1.n0209 [9], \xm8051_golden_model_1.aes_bytes_processed [9]);
  buf(\xm8051_golden_model_1.n0209 [10], \xm8051_golden_model_1.aes_bytes_processed [10]);
  buf(\xm8051_golden_model_1.n0209 [11], \xm8051_golden_model_1.aes_bytes_processed [11]);
  buf(\xm8051_golden_model_1.n0209 [12], \xm8051_golden_model_1.aes_bytes_processed [12]);
  buf(\xm8051_golden_model_1.n0209 [13], \xm8051_golden_model_1.aes_bytes_processed [13]);
  buf(\xm8051_golden_model_1.n0209 [14], \xm8051_golden_model_1.aes_bytes_processed [14]);
  buf(\xm8051_golden_model_1.n0209 [15], \xm8051_golden_model_1.aes_bytes_processed [15]);
  buf(\xm8051_golden_model_1.n1244 [0], input_sha_func_19[0]);
  buf(\xm8051_golden_model_1.n1244 [1], input_sha_func_19[1]);
  buf(\xm8051_golden_model_1.n1244 [2], input_sha_func_19[2]);
  buf(\xm8051_golden_model_1.n1244 [3], input_sha_func_19[3]);
  buf(\xm8051_golden_model_1.n1244 [4], input_sha_func_19[4]);
  buf(\xm8051_golden_model_1.n1244 [5], input_sha_func_19[5]);
  buf(\xm8051_golden_model_1.n1244 [6], input_sha_func_19[6]);
  buf(\xm8051_golden_model_1.n1244 [7], input_sha_func_19[7]);
  buf(\xm8051_golden_model_1.n1244 [8], input_sha_func_19[8]);
  buf(\xm8051_golden_model_1.n1244 [9], input_sha_func_19[9]);
  buf(\xm8051_golden_model_1.n1244 [10], input_sha_func_19[10]);
  buf(\xm8051_golden_model_1.n1244 [11], input_sha_func_19[11]);
  buf(\xm8051_golden_model_1.n1244 [12], input_sha_func_19[12]);
  buf(\xm8051_golden_model_1.n1244 [13], input_sha_func_19[13]);
  buf(\xm8051_golden_model_1.n1244 [14], input_sha_func_19[14]);
  buf(\xm8051_golden_model_1.n1244 [15], input_sha_func_19[15]);
  buf(\xm8051_golden_model_1.n1244 [16], input_sha_func_19[16]);
  buf(\xm8051_golden_model_1.n1244 [17], input_sha_func_19[17]);
  buf(\xm8051_golden_model_1.n1244 [18], input_sha_func_19[18]);
  buf(\xm8051_golden_model_1.n1244 [19], input_sha_func_19[19]);
  buf(\xm8051_golden_model_1.n1244 [20], input_sha_func_19[20]);
  buf(\xm8051_golden_model_1.n1244 [21], input_sha_func_19[21]);
  buf(\xm8051_golden_model_1.n1244 [22], input_sha_func_19[22]);
  buf(\xm8051_golden_model_1.n1244 [23], input_sha_func_19[23]);
  buf(\xm8051_golden_model_1.n1244 [24], input_sha_func_19[24]);
  buf(\xm8051_golden_model_1.n1244 [25], input_sha_func_19[25]);
  buf(\xm8051_golden_model_1.n1244 [26], input_sha_func_19[26]);
  buf(\xm8051_golden_model_1.n1244 [27], input_sha_func_19[27]);
  buf(\xm8051_golden_model_1.n1244 [28], input_sha_func_19[28]);
  buf(\xm8051_golden_model_1.n1244 [29], input_sha_func_19[29]);
  buf(\xm8051_golden_model_1.n1244 [30], input_sha_func_19[30]);
  buf(\xm8051_golden_model_1.n1244 [31], input_sha_func_19[31]);
  buf(\xm8051_golden_model_1.n1244 [32], input_sha_func_18[0]);
  buf(\xm8051_golden_model_1.n1244 [33], input_sha_func_18[1]);
  buf(\xm8051_golden_model_1.n1244 [34], input_sha_func_18[2]);
  buf(\xm8051_golden_model_1.n1244 [35], input_sha_func_18[3]);
  buf(\xm8051_golden_model_1.n1244 [36], input_sha_func_18[4]);
  buf(\xm8051_golden_model_1.n1244 [37], input_sha_func_18[5]);
  buf(\xm8051_golden_model_1.n1244 [38], input_sha_func_18[6]);
  buf(\xm8051_golden_model_1.n1244 [39], input_sha_func_18[7]);
  buf(\xm8051_golden_model_1.n1244 [40], input_sha_func_18[8]);
  buf(\xm8051_golden_model_1.n1244 [41], input_sha_func_18[9]);
  buf(\xm8051_golden_model_1.n1244 [42], input_sha_func_18[10]);
  buf(\xm8051_golden_model_1.n1244 [43], input_sha_func_18[11]);
  buf(\xm8051_golden_model_1.n1244 [44], input_sha_func_18[12]);
  buf(\xm8051_golden_model_1.n1244 [45], input_sha_func_18[13]);
  buf(\xm8051_golden_model_1.n1244 [46], input_sha_func_18[14]);
  buf(\xm8051_golden_model_1.n1244 [47], input_sha_func_18[15]);
  buf(\xm8051_golden_model_1.n1244 [48], input_sha_func_18[16]);
  buf(\xm8051_golden_model_1.n1244 [49], input_sha_func_18[17]);
  buf(\xm8051_golden_model_1.n1244 [50], input_sha_func_18[18]);
  buf(\xm8051_golden_model_1.n1244 [51], input_sha_func_18[19]);
  buf(\xm8051_golden_model_1.n1244 [52], input_sha_func_18[20]);
  buf(\xm8051_golden_model_1.n1244 [53], input_sha_func_18[21]);
  buf(\xm8051_golden_model_1.n1244 [54], input_sha_func_18[22]);
  buf(\xm8051_golden_model_1.n1244 [55], input_sha_func_18[23]);
  buf(\xm8051_golden_model_1.n1244 [56], input_sha_func_18[24]);
  buf(\xm8051_golden_model_1.n1244 [57], input_sha_func_18[25]);
  buf(\xm8051_golden_model_1.n1244 [58], input_sha_func_18[26]);
  buf(\xm8051_golden_model_1.n1244 [59], input_sha_func_18[27]);
  buf(\xm8051_golden_model_1.n1244 [60], input_sha_func_18[28]);
  buf(\xm8051_golden_model_1.n1244 [61], input_sha_func_18[29]);
  buf(\xm8051_golden_model_1.n1244 [62], input_sha_func_18[30]);
  buf(\xm8051_golden_model_1.n1244 [63], input_sha_func_18[31]);
  buf(\xm8051_golden_model_1.n1244 [64], input_sha_func_18[32]);
  buf(\xm8051_golden_model_1.n1244 [65], input_sha_func_18[33]);
  buf(\xm8051_golden_model_1.n1244 [66], input_sha_func_18[34]);
  buf(\xm8051_golden_model_1.n1244 [67], input_sha_func_18[35]);
  buf(\xm8051_golden_model_1.n1244 [68], input_sha_func_18[36]);
  buf(\xm8051_golden_model_1.n1244 [69], input_sha_func_18[37]);
  buf(\xm8051_golden_model_1.n1244 [70], input_sha_func_18[38]);
  buf(\xm8051_golden_model_1.n1244 [71], input_sha_func_18[39]);
  buf(\xm8051_golden_model_1.n1244 [72], input_sha_func_18[40]);
  buf(\xm8051_golden_model_1.n1244 [73], input_sha_func_18[41]);
  buf(\xm8051_golden_model_1.n1244 [74], input_sha_func_18[42]);
  buf(\xm8051_golden_model_1.n1244 [75], input_sha_func_18[43]);
  buf(\xm8051_golden_model_1.n1244 [76], input_sha_func_18[44]);
  buf(\xm8051_golden_model_1.n1244 [77], input_sha_func_18[45]);
  buf(\xm8051_golden_model_1.n1244 [78], input_sha_func_18[46]);
  buf(\xm8051_golden_model_1.n1244 [79], input_sha_func_18[47]);
  buf(\xm8051_golden_model_1.n1244 [80], input_sha_func_18[48]);
  buf(\xm8051_golden_model_1.n1244 [81], input_sha_func_18[49]);
  buf(\xm8051_golden_model_1.n1244 [82], input_sha_func_18[50]);
  buf(\xm8051_golden_model_1.n1244 [83], input_sha_func_18[51]);
  buf(\xm8051_golden_model_1.n1244 [84], input_sha_func_18[52]);
  buf(\xm8051_golden_model_1.n1244 [85], input_sha_func_18[53]);
  buf(\xm8051_golden_model_1.n1244 [86], input_sha_func_18[54]);
  buf(\xm8051_golden_model_1.n1244 [87], input_sha_func_18[55]);
  buf(\xm8051_golden_model_1.n1244 [88], input_sha_func_18[56]);
  buf(\xm8051_golden_model_1.n1244 [89], input_sha_func_18[57]);
  buf(\xm8051_golden_model_1.n1244 [90], input_sha_func_18[58]);
  buf(\xm8051_golden_model_1.n1244 [91], input_sha_func_18[59]);
  buf(\xm8051_golden_model_1.n1244 [92], input_sha_func_18[60]);
  buf(\xm8051_golden_model_1.n1244 [93], input_sha_func_18[61]);
  buf(\xm8051_golden_model_1.n1244 [94], input_sha_func_18[62]);
  buf(\xm8051_golden_model_1.n1244 [95], input_sha_func_18[63]);
  buf(\xm8051_golden_model_1.n1244 [96], input_sha_func_17[0]);
  buf(\xm8051_golden_model_1.n1244 [97], input_sha_func_17[1]);
  buf(\xm8051_golden_model_1.n1244 [98], input_sha_func_17[2]);
  buf(\xm8051_golden_model_1.n1244 [99], input_sha_func_17[3]);
  buf(\xm8051_golden_model_1.n1244 [100], input_sha_func_17[4]);
  buf(\xm8051_golden_model_1.n1244 [101], input_sha_func_17[5]);
  buf(\xm8051_golden_model_1.n1244 [102], input_sha_func_17[6]);
  buf(\xm8051_golden_model_1.n1244 [103], input_sha_func_17[7]);
  buf(\xm8051_golden_model_1.n1244 [104], input_sha_func_17[8]);
  buf(\xm8051_golden_model_1.n1244 [105], input_sha_func_17[9]);
  buf(\xm8051_golden_model_1.n1244 [106], input_sha_func_17[10]);
  buf(\xm8051_golden_model_1.n1244 [107], input_sha_func_17[11]);
  buf(\xm8051_golden_model_1.n1244 [108], input_sha_func_17[12]);
  buf(\xm8051_golden_model_1.n1244 [109], input_sha_func_17[13]);
  buf(\xm8051_golden_model_1.n1244 [110], input_sha_func_17[14]);
  buf(\xm8051_golden_model_1.n1244 [111], input_sha_func_17[15]);
  buf(\xm8051_golden_model_1.n1244 [112], input_sha_func_17[16]);
  buf(\xm8051_golden_model_1.n1244 [113], input_sha_func_17[17]);
  buf(\xm8051_golden_model_1.n1244 [114], input_sha_func_17[18]);
  buf(\xm8051_golden_model_1.n1244 [115], input_sha_func_17[19]);
  buf(\xm8051_golden_model_1.n1244 [116], input_sha_func_17[20]);
  buf(\xm8051_golden_model_1.n1244 [117], input_sha_func_17[21]);
  buf(\xm8051_golden_model_1.n1244 [118], input_sha_func_17[22]);
  buf(\xm8051_golden_model_1.n1244 [119], input_sha_func_17[23]);
  buf(\xm8051_golden_model_1.n1244 [120], input_sha_func_17[24]);
  buf(\xm8051_golden_model_1.n1244 [121], input_sha_func_17[25]);
  buf(\xm8051_golden_model_1.n1244 [122], input_sha_func_17[26]);
  buf(\xm8051_golden_model_1.n1244 [123], input_sha_func_17[27]);
  buf(\xm8051_golden_model_1.n1244 [124], input_sha_func_17[28]);
  buf(\xm8051_golden_model_1.n1244 [125], input_sha_func_17[29]);
  buf(\xm8051_golden_model_1.n1244 [126], input_sha_func_17[30]);
  buf(\xm8051_golden_model_1.n1244 [127], input_sha_func_17[31]);
  buf(\xm8051_golden_model_1.n1244 [128], input_sha_func_17[32]);
  buf(\xm8051_golden_model_1.n1244 [129], input_sha_func_17[33]);
  buf(\xm8051_golden_model_1.n1244 [130], input_sha_func_17[34]);
  buf(\xm8051_golden_model_1.n1244 [131], input_sha_func_17[35]);
  buf(\xm8051_golden_model_1.n1244 [132], input_sha_func_17[36]);
  buf(\xm8051_golden_model_1.n1244 [133], input_sha_func_17[37]);
  buf(\xm8051_golden_model_1.n1244 [134], input_sha_func_17[38]);
  buf(\xm8051_golden_model_1.n1244 [135], input_sha_func_17[39]);
  buf(\xm8051_golden_model_1.n1244 [136], input_sha_func_17[40]);
  buf(\xm8051_golden_model_1.n1244 [137], input_sha_func_17[41]);
  buf(\xm8051_golden_model_1.n1244 [138], input_sha_func_17[42]);
  buf(\xm8051_golden_model_1.n1244 [139], input_sha_func_17[43]);
  buf(\xm8051_golden_model_1.n1244 [140], input_sha_func_17[44]);
  buf(\xm8051_golden_model_1.n1244 [141], input_sha_func_17[45]);
  buf(\xm8051_golden_model_1.n1244 [142], input_sha_func_17[46]);
  buf(\xm8051_golden_model_1.n1244 [143], input_sha_func_17[47]);
  buf(\xm8051_golden_model_1.n1244 [144], input_sha_func_17[48]);
  buf(\xm8051_golden_model_1.n1244 [145], input_sha_func_17[49]);
  buf(\xm8051_golden_model_1.n1244 [146], input_sha_func_17[50]);
  buf(\xm8051_golden_model_1.n1244 [147], input_sha_func_17[51]);
  buf(\xm8051_golden_model_1.n1244 [148], input_sha_func_17[52]);
  buf(\xm8051_golden_model_1.n1244 [149], input_sha_func_17[53]);
  buf(\xm8051_golden_model_1.n1244 [150], input_sha_func_17[54]);
  buf(\xm8051_golden_model_1.n1244 [151], input_sha_func_17[55]);
  buf(\xm8051_golden_model_1.n1244 [152], input_sha_func_17[56]);
  buf(\xm8051_golden_model_1.n1244 [153], input_sha_func_17[57]);
  buf(\xm8051_golden_model_1.n1244 [154], input_sha_func_17[58]);
  buf(\xm8051_golden_model_1.n1244 [155], input_sha_func_17[59]);
  buf(\xm8051_golden_model_1.n1244 [156], input_sha_func_17[60]);
  buf(\xm8051_golden_model_1.n1244 [157], input_sha_func_17[61]);
  buf(\xm8051_golden_model_1.n1244 [158], input_sha_func_17[62]);
  buf(\xm8051_golden_model_1.n1244 [159], input_sha_func_17[63]);
  buf(\xm8051_golden_model_1.n1240 [0], RD_xram_64[0]);
  buf(\xm8051_golden_model_1.n1240 [1], RD_xram_64[1]);
  buf(\xm8051_golden_model_1.n1240 [2], RD_xram_64[2]);
  buf(\xm8051_golden_model_1.n1240 [3], RD_xram_64[3]);
  buf(\xm8051_golden_model_1.n1240 [4], RD_xram_64[4]);
  buf(\xm8051_golden_model_1.n1240 [5], RD_xram_64[5]);
  buf(\xm8051_golden_model_1.n1240 [6], RD_xram_64[6]);
  buf(\xm8051_golden_model_1.n1240 [7], RD_xram_64[7]);
  buf(\xm8051_golden_model_1.n1240 [8], RD_xram_63[0]);
  buf(\xm8051_golden_model_1.n1240 [9], RD_xram_63[1]);
  buf(\xm8051_golden_model_1.n1240 [10], RD_xram_63[2]);
  buf(\xm8051_golden_model_1.n1240 [11], RD_xram_63[3]);
  buf(\xm8051_golden_model_1.n1240 [12], RD_xram_63[4]);
  buf(\xm8051_golden_model_1.n1240 [13], RD_xram_63[5]);
  buf(\xm8051_golden_model_1.n1240 [14], RD_xram_63[6]);
  buf(\xm8051_golden_model_1.n1240 [15], RD_xram_63[7]);
  buf(\xm8051_golden_model_1.n1240 [16], RD_xram_62[0]);
  buf(\xm8051_golden_model_1.n1240 [17], RD_xram_62[1]);
  buf(\xm8051_golden_model_1.n1240 [18], RD_xram_62[2]);
  buf(\xm8051_golden_model_1.n1240 [19], RD_xram_62[3]);
  buf(\xm8051_golden_model_1.n1240 [20], RD_xram_62[4]);
  buf(\xm8051_golden_model_1.n1240 [21], RD_xram_62[5]);
  buf(\xm8051_golden_model_1.n1240 [22], RD_xram_62[6]);
  buf(\xm8051_golden_model_1.n1240 [23], RD_xram_62[7]);
  buf(\xm8051_golden_model_1.n1240 [24], RD_xram_61[0]);
  buf(\xm8051_golden_model_1.n1240 [25], RD_xram_61[1]);
  buf(\xm8051_golden_model_1.n1240 [26], RD_xram_61[2]);
  buf(\xm8051_golden_model_1.n1240 [27], RD_xram_61[3]);
  buf(\xm8051_golden_model_1.n1240 [28], RD_xram_61[4]);
  buf(\xm8051_golden_model_1.n1240 [29], RD_xram_61[5]);
  buf(\xm8051_golden_model_1.n1240 [30], RD_xram_61[6]);
  buf(\xm8051_golden_model_1.n1240 [31], RD_xram_61[7]);
  buf(\xm8051_golden_model_1.n1240 [32], RD_xram_60[0]);
  buf(\xm8051_golden_model_1.n1240 [33], RD_xram_60[1]);
  buf(\xm8051_golden_model_1.n1240 [34], RD_xram_60[2]);
  buf(\xm8051_golden_model_1.n1240 [35], RD_xram_60[3]);
  buf(\xm8051_golden_model_1.n1240 [36], RD_xram_60[4]);
  buf(\xm8051_golden_model_1.n1240 [37], RD_xram_60[5]);
  buf(\xm8051_golden_model_1.n1240 [38], RD_xram_60[6]);
  buf(\xm8051_golden_model_1.n1240 [39], RD_xram_60[7]);
  buf(\xm8051_golden_model_1.n1240 [40], RD_xram_59[0]);
  buf(\xm8051_golden_model_1.n1240 [41], RD_xram_59[1]);
  buf(\xm8051_golden_model_1.n1240 [42], RD_xram_59[2]);
  buf(\xm8051_golden_model_1.n1240 [43], RD_xram_59[3]);
  buf(\xm8051_golden_model_1.n1240 [44], RD_xram_59[4]);
  buf(\xm8051_golden_model_1.n1240 [45], RD_xram_59[5]);
  buf(\xm8051_golden_model_1.n1240 [46], RD_xram_59[6]);
  buf(\xm8051_golden_model_1.n1240 [47], RD_xram_59[7]);
  buf(\xm8051_golden_model_1.n1240 [48], RD_xram_58[0]);
  buf(\xm8051_golden_model_1.n1240 [49], RD_xram_58[1]);
  buf(\xm8051_golden_model_1.n1240 [50], RD_xram_58[2]);
  buf(\xm8051_golden_model_1.n1240 [51], RD_xram_58[3]);
  buf(\xm8051_golden_model_1.n1240 [52], RD_xram_58[4]);
  buf(\xm8051_golden_model_1.n1240 [53], RD_xram_58[5]);
  buf(\xm8051_golden_model_1.n1240 [54], RD_xram_58[6]);
  buf(\xm8051_golden_model_1.n1240 [55], RD_xram_58[7]);
  buf(\xm8051_golden_model_1.n1240 [56], RD_xram_57[0]);
  buf(\xm8051_golden_model_1.n1240 [57], RD_xram_57[1]);
  buf(\xm8051_golden_model_1.n1240 [58], RD_xram_57[2]);
  buf(\xm8051_golden_model_1.n1240 [59], RD_xram_57[3]);
  buf(\xm8051_golden_model_1.n1240 [60], RD_xram_57[4]);
  buf(\xm8051_golden_model_1.n1240 [61], RD_xram_57[5]);
  buf(\xm8051_golden_model_1.n1240 [62], RD_xram_57[6]);
  buf(\xm8051_golden_model_1.n1240 [63], RD_xram_57[7]);
  buf(\xm8051_golden_model_1.n1240 [64], RD_xram_56[0]);
  buf(\xm8051_golden_model_1.n1240 [65], RD_xram_56[1]);
  buf(\xm8051_golden_model_1.n1240 [66], RD_xram_56[2]);
  buf(\xm8051_golden_model_1.n1240 [67], RD_xram_56[3]);
  buf(\xm8051_golden_model_1.n1240 [68], RD_xram_56[4]);
  buf(\xm8051_golden_model_1.n1240 [69], RD_xram_56[5]);
  buf(\xm8051_golden_model_1.n1240 [70], RD_xram_56[6]);
  buf(\xm8051_golden_model_1.n1240 [71], RD_xram_56[7]);
  buf(\xm8051_golden_model_1.n1240 [72], RD_xram_55[0]);
  buf(\xm8051_golden_model_1.n1240 [73], RD_xram_55[1]);
  buf(\xm8051_golden_model_1.n1240 [74], RD_xram_55[2]);
  buf(\xm8051_golden_model_1.n1240 [75], RD_xram_55[3]);
  buf(\xm8051_golden_model_1.n1240 [76], RD_xram_55[4]);
  buf(\xm8051_golden_model_1.n1240 [77], RD_xram_55[5]);
  buf(\xm8051_golden_model_1.n1240 [78], RD_xram_55[6]);
  buf(\xm8051_golden_model_1.n1240 [79], RD_xram_55[7]);
  buf(\xm8051_golden_model_1.n1240 [80], RD_xram_54[0]);
  buf(\xm8051_golden_model_1.n1240 [81], RD_xram_54[1]);
  buf(\xm8051_golden_model_1.n1240 [82], RD_xram_54[2]);
  buf(\xm8051_golden_model_1.n1240 [83], RD_xram_54[3]);
  buf(\xm8051_golden_model_1.n1240 [84], RD_xram_54[4]);
  buf(\xm8051_golden_model_1.n1240 [85], RD_xram_54[5]);
  buf(\xm8051_golden_model_1.n1240 [86], RD_xram_54[6]);
  buf(\xm8051_golden_model_1.n1240 [87], RD_xram_54[7]);
  buf(\xm8051_golden_model_1.n1240 [88], RD_xram_53[0]);
  buf(\xm8051_golden_model_1.n1240 [89], RD_xram_53[1]);
  buf(\xm8051_golden_model_1.n1240 [90], RD_xram_53[2]);
  buf(\xm8051_golden_model_1.n1240 [91], RD_xram_53[3]);
  buf(\xm8051_golden_model_1.n1240 [92], RD_xram_53[4]);
  buf(\xm8051_golden_model_1.n1240 [93], RD_xram_53[5]);
  buf(\xm8051_golden_model_1.n1240 [94], RD_xram_53[6]);
  buf(\xm8051_golden_model_1.n1240 [95], RD_xram_53[7]);
  buf(\xm8051_golden_model_1.n1240 [96], RD_xram_52[0]);
  buf(\xm8051_golden_model_1.n1240 [97], RD_xram_52[1]);
  buf(\xm8051_golden_model_1.n1240 [98], RD_xram_52[2]);
  buf(\xm8051_golden_model_1.n1240 [99], RD_xram_52[3]);
  buf(\xm8051_golden_model_1.n1240 [100], RD_xram_52[4]);
  buf(\xm8051_golden_model_1.n1240 [101], RD_xram_52[5]);
  buf(\xm8051_golden_model_1.n1240 [102], RD_xram_52[6]);
  buf(\xm8051_golden_model_1.n1240 [103], RD_xram_52[7]);
  buf(\xm8051_golden_model_1.n1240 [104], RD_xram_51[0]);
  buf(\xm8051_golden_model_1.n1240 [105], RD_xram_51[1]);
  buf(\xm8051_golden_model_1.n1240 [106], RD_xram_51[2]);
  buf(\xm8051_golden_model_1.n1240 [107], RD_xram_51[3]);
  buf(\xm8051_golden_model_1.n1240 [108], RD_xram_51[4]);
  buf(\xm8051_golden_model_1.n1240 [109], RD_xram_51[5]);
  buf(\xm8051_golden_model_1.n1240 [110], RD_xram_51[6]);
  buf(\xm8051_golden_model_1.n1240 [111], RD_xram_51[7]);
  buf(\xm8051_golden_model_1.n1240 [112], RD_xram_50[0]);
  buf(\xm8051_golden_model_1.n1240 [113], RD_xram_50[1]);
  buf(\xm8051_golden_model_1.n1240 [114], RD_xram_50[2]);
  buf(\xm8051_golden_model_1.n1240 [115], RD_xram_50[3]);
  buf(\xm8051_golden_model_1.n1240 [116], RD_xram_50[4]);
  buf(\xm8051_golden_model_1.n1240 [117], RD_xram_50[5]);
  buf(\xm8051_golden_model_1.n1240 [118], RD_xram_50[6]);
  buf(\xm8051_golden_model_1.n1240 [119], RD_xram_50[7]);
  buf(\xm8051_golden_model_1.n1240 [120], RD_xram_49[0]);
  buf(\xm8051_golden_model_1.n1240 [121], RD_xram_49[1]);
  buf(\xm8051_golden_model_1.n1240 [122], RD_xram_49[2]);
  buf(\xm8051_golden_model_1.n1240 [123], RD_xram_49[3]);
  buf(\xm8051_golden_model_1.n1240 [124], RD_xram_49[4]);
  buf(\xm8051_golden_model_1.n1240 [125], RD_xram_49[5]);
  buf(\xm8051_golden_model_1.n1240 [126], RD_xram_49[6]);
  buf(\xm8051_golden_model_1.n1240 [127], RD_xram_49[7]);
  buf(\xm8051_golden_model_1.n1240 [128], RD_xram_48[0]);
  buf(\xm8051_golden_model_1.n1240 [129], RD_xram_48[1]);
  buf(\xm8051_golden_model_1.n1240 [130], RD_xram_48[2]);
  buf(\xm8051_golden_model_1.n1240 [131], RD_xram_48[3]);
  buf(\xm8051_golden_model_1.n1240 [132], RD_xram_48[4]);
  buf(\xm8051_golden_model_1.n1240 [133], RD_xram_48[5]);
  buf(\xm8051_golden_model_1.n1240 [134], RD_xram_48[6]);
  buf(\xm8051_golden_model_1.n1240 [135], RD_xram_48[7]);
  buf(\xm8051_golden_model_1.n1240 [136], RD_xram_47[0]);
  buf(\xm8051_golden_model_1.n1240 [137], RD_xram_47[1]);
  buf(\xm8051_golden_model_1.n1240 [138], RD_xram_47[2]);
  buf(\xm8051_golden_model_1.n1240 [139], RD_xram_47[3]);
  buf(\xm8051_golden_model_1.n1240 [140], RD_xram_47[4]);
  buf(\xm8051_golden_model_1.n1240 [141], RD_xram_47[5]);
  buf(\xm8051_golden_model_1.n1240 [142], RD_xram_47[6]);
  buf(\xm8051_golden_model_1.n1240 [143], RD_xram_47[7]);
  buf(\xm8051_golden_model_1.n1240 [144], RD_xram_46[0]);
  buf(\xm8051_golden_model_1.n1240 [145], RD_xram_46[1]);
  buf(\xm8051_golden_model_1.n1240 [146], RD_xram_46[2]);
  buf(\xm8051_golden_model_1.n1240 [147], RD_xram_46[3]);
  buf(\xm8051_golden_model_1.n1240 [148], RD_xram_46[4]);
  buf(\xm8051_golden_model_1.n1240 [149], RD_xram_46[5]);
  buf(\xm8051_golden_model_1.n1240 [150], RD_xram_46[6]);
  buf(\xm8051_golden_model_1.n1240 [151], RD_xram_46[7]);
  buf(\xm8051_golden_model_1.n1240 [152], RD_xram_45[0]);
  buf(\xm8051_golden_model_1.n1240 [153], RD_xram_45[1]);
  buf(\xm8051_golden_model_1.n1240 [154], RD_xram_45[2]);
  buf(\xm8051_golden_model_1.n1240 [155], RD_xram_45[3]);
  buf(\xm8051_golden_model_1.n1240 [156], RD_xram_45[4]);
  buf(\xm8051_golden_model_1.n1240 [157], RD_xram_45[5]);
  buf(\xm8051_golden_model_1.n1240 [158], RD_xram_45[6]);
  buf(\xm8051_golden_model_1.n1240 [159], RD_xram_45[7]);
  buf(\xm8051_golden_model_1.n1240 [160], RD_xram_44[0]);
  buf(\xm8051_golden_model_1.n1240 [161], RD_xram_44[1]);
  buf(\xm8051_golden_model_1.n1240 [162], RD_xram_44[2]);
  buf(\xm8051_golden_model_1.n1240 [163], RD_xram_44[3]);
  buf(\xm8051_golden_model_1.n1240 [164], RD_xram_44[4]);
  buf(\xm8051_golden_model_1.n1240 [165], RD_xram_44[5]);
  buf(\xm8051_golden_model_1.n1240 [166], RD_xram_44[6]);
  buf(\xm8051_golden_model_1.n1240 [167], RD_xram_44[7]);
  buf(\xm8051_golden_model_1.n1240 [168], RD_xram_43[0]);
  buf(\xm8051_golden_model_1.n1240 [169], RD_xram_43[1]);
  buf(\xm8051_golden_model_1.n1240 [170], RD_xram_43[2]);
  buf(\xm8051_golden_model_1.n1240 [171], RD_xram_43[3]);
  buf(\xm8051_golden_model_1.n1240 [172], RD_xram_43[4]);
  buf(\xm8051_golden_model_1.n1240 [173], RD_xram_43[5]);
  buf(\xm8051_golden_model_1.n1240 [174], RD_xram_43[6]);
  buf(\xm8051_golden_model_1.n1240 [175], RD_xram_43[7]);
  buf(\xm8051_golden_model_1.n1240 [176], RD_xram_42[0]);
  buf(\xm8051_golden_model_1.n1240 [177], RD_xram_42[1]);
  buf(\xm8051_golden_model_1.n1240 [178], RD_xram_42[2]);
  buf(\xm8051_golden_model_1.n1240 [179], RD_xram_42[3]);
  buf(\xm8051_golden_model_1.n1240 [180], RD_xram_42[4]);
  buf(\xm8051_golden_model_1.n1240 [181], RD_xram_42[5]);
  buf(\xm8051_golden_model_1.n1240 [182], RD_xram_42[6]);
  buf(\xm8051_golden_model_1.n1240 [183], RD_xram_42[7]);
  buf(\xm8051_golden_model_1.n1240 [184], RD_xram_41[0]);
  buf(\xm8051_golden_model_1.n1240 [185], RD_xram_41[1]);
  buf(\xm8051_golden_model_1.n1240 [186], RD_xram_41[2]);
  buf(\xm8051_golden_model_1.n1240 [187], RD_xram_41[3]);
  buf(\xm8051_golden_model_1.n1240 [188], RD_xram_41[4]);
  buf(\xm8051_golden_model_1.n1240 [189], RD_xram_41[5]);
  buf(\xm8051_golden_model_1.n1240 [190], RD_xram_41[6]);
  buf(\xm8051_golden_model_1.n1240 [191], RD_xram_41[7]);
  buf(\xm8051_golden_model_1.n1240 [192], RD_xram_40[0]);
  buf(\xm8051_golden_model_1.n1240 [193], RD_xram_40[1]);
  buf(\xm8051_golden_model_1.n1240 [194], RD_xram_40[2]);
  buf(\xm8051_golden_model_1.n1240 [195], RD_xram_40[3]);
  buf(\xm8051_golden_model_1.n1240 [196], RD_xram_40[4]);
  buf(\xm8051_golden_model_1.n1240 [197], RD_xram_40[5]);
  buf(\xm8051_golden_model_1.n1240 [198], RD_xram_40[6]);
  buf(\xm8051_golden_model_1.n1240 [199], RD_xram_40[7]);
  buf(\xm8051_golden_model_1.n1240 [200], RD_xram_39[0]);
  buf(\xm8051_golden_model_1.n1240 [201], RD_xram_39[1]);
  buf(\xm8051_golden_model_1.n1240 [202], RD_xram_39[2]);
  buf(\xm8051_golden_model_1.n1240 [203], RD_xram_39[3]);
  buf(\xm8051_golden_model_1.n1240 [204], RD_xram_39[4]);
  buf(\xm8051_golden_model_1.n1240 [205], RD_xram_39[5]);
  buf(\xm8051_golden_model_1.n1240 [206], RD_xram_39[6]);
  buf(\xm8051_golden_model_1.n1240 [207], RD_xram_39[7]);
  buf(\xm8051_golden_model_1.n1240 [208], RD_xram_38[0]);
  buf(\xm8051_golden_model_1.n1240 [209], RD_xram_38[1]);
  buf(\xm8051_golden_model_1.n1240 [210], RD_xram_38[2]);
  buf(\xm8051_golden_model_1.n1240 [211], RD_xram_38[3]);
  buf(\xm8051_golden_model_1.n1240 [212], RD_xram_38[4]);
  buf(\xm8051_golden_model_1.n1240 [213], RD_xram_38[5]);
  buf(\xm8051_golden_model_1.n1240 [214], RD_xram_38[6]);
  buf(\xm8051_golden_model_1.n1240 [215], RD_xram_38[7]);
  buf(\xm8051_golden_model_1.n1240 [216], RD_xram_37[0]);
  buf(\xm8051_golden_model_1.n1240 [217], RD_xram_37[1]);
  buf(\xm8051_golden_model_1.n1240 [218], RD_xram_37[2]);
  buf(\xm8051_golden_model_1.n1240 [219], RD_xram_37[3]);
  buf(\xm8051_golden_model_1.n1240 [220], RD_xram_37[4]);
  buf(\xm8051_golden_model_1.n1240 [221], RD_xram_37[5]);
  buf(\xm8051_golden_model_1.n1240 [222], RD_xram_37[6]);
  buf(\xm8051_golden_model_1.n1240 [223], RD_xram_37[7]);
  buf(\xm8051_golden_model_1.n1240 [224], RD_xram_36[0]);
  buf(\xm8051_golden_model_1.n1240 [225], RD_xram_36[1]);
  buf(\xm8051_golden_model_1.n1240 [226], RD_xram_36[2]);
  buf(\xm8051_golden_model_1.n1240 [227], RD_xram_36[3]);
  buf(\xm8051_golden_model_1.n1240 [228], RD_xram_36[4]);
  buf(\xm8051_golden_model_1.n1240 [229], RD_xram_36[5]);
  buf(\xm8051_golden_model_1.n1240 [230], RD_xram_36[6]);
  buf(\xm8051_golden_model_1.n1240 [231], RD_xram_36[7]);
  buf(\xm8051_golden_model_1.n1240 [232], RD_xram_35[0]);
  buf(\xm8051_golden_model_1.n1240 [233], RD_xram_35[1]);
  buf(\xm8051_golden_model_1.n1240 [234], RD_xram_35[2]);
  buf(\xm8051_golden_model_1.n1240 [235], RD_xram_35[3]);
  buf(\xm8051_golden_model_1.n1240 [236], RD_xram_35[4]);
  buf(\xm8051_golden_model_1.n1240 [237], RD_xram_35[5]);
  buf(\xm8051_golden_model_1.n1240 [238], RD_xram_35[6]);
  buf(\xm8051_golden_model_1.n1240 [239], RD_xram_35[7]);
  buf(\xm8051_golden_model_1.n1240 [240], RD_xram_34[0]);
  buf(\xm8051_golden_model_1.n1240 [241], RD_xram_34[1]);
  buf(\xm8051_golden_model_1.n1240 [242], RD_xram_34[2]);
  buf(\xm8051_golden_model_1.n1240 [243], RD_xram_34[3]);
  buf(\xm8051_golden_model_1.n1240 [244], RD_xram_34[4]);
  buf(\xm8051_golden_model_1.n1240 [245], RD_xram_34[5]);
  buf(\xm8051_golden_model_1.n1240 [246], RD_xram_34[6]);
  buf(\xm8051_golden_model_1.n1240 [247], RD_xram_34[7]);
  buf(\xm8051_golden_model_1.n1240 [248], RD_xram_33[0]);
  buf(\xm8051_golden_model_1.n1240 [249], RD_xram_33[1]);
  buf(\xm8051_golden_model_1.n1240 [250], RD_xram_33[2]);
  buf(\xm8051_golden_model_1.n1240 [251], RD_xram_33[3]);
  buf(\xm8051_golden_model_1.n1240 [252], RD_xram_33[4]);
  buf(\xm8051_golden_model_1.n1240 [253], RD_xram_33[5]);
  buf(\xm8051_golden_model_1.n1240 [254], RD_xram_33[6]);
  buf(\xm8051_golden_model_1.n1240 [255], RD_xram_33[7]);
  buf(\xm8051_golden_model_1.n1240 [256], RD_xram_32[0]);
  buf(\xm8051_golden_model_1.n1240 [257], RD_xram_32[1]);
  buf(\xm8051_golden_model_1.n1240 [258], RD_xram_32[2]);
  buf(\xm8051_golden_model_1.n1240 [259], RD_xram_32[3]);
  buf(\xm8051_golden_model_1.n1240 [260], RD_xram_32[4]);
  buf(\xm8051_golden_model_1.n1240 [261], RD_xram_32[5]);
  buf(\xm8051_golden_model_1.n1240 [262], RD_xram_32[6]);
  buf(\xm8051_golden_model_1.n1240 [263], RD_xram_32[7]);
  buf(\xm8051_golden_model_1.n1240 [264], RD_xram_31[0]);
  buf(\xm8051_golden_model_1.n1240 [265], RD_xram_31[1]);
  buf(\xm8051_golden_model_1.n1240 [266], RD_xram_31[2]);
  buf(\xm8051_golden_model_1.n1240 [267], RD_xram_31[3]);
  buf(\xm8051_golden_model_1.n1240 [268], RD_xram_31[4]);
  buf(\xm8051_golden_model_1.n1240 [269], RD_xram_31[5]);
  buf(\xm8051_golden_model_1.n1240 [270], RD_xram_31[6]);
  buf(\xm8051_golden_model_1.n1240 [271], RD_xram_31[7]);
  buf(\xm8051_golden_model_1.n1240 [272], RD_xram_30[0]);
  buf(\xm8051_golden_model_1.n1240 [273], RD_xram_30[1]);
  buf(\xm8051_golden_model_1.n1240 [274], RD_xram_30[2]);
  buf(\xm8051_golden_model_1.n1240 [275], RD_xram_30[3]);
  buf(\xm8051_golden_model_1.n1240 [276], RD_xram_30[4]);
  buf(\xm8051_golden_model_1.n1240 [277], RD_xram_30[5]);
  buf(\xm8051_golden_model_1.n1240 [278], RD_xram_30[6]);
  buf(\xm8051_golden_model_1.n1240 [279], RD_xram_30[7]);
  buf(\xm8051_golden_model_1.n1240 [280], RD_xram_29[0]);
  buf(\xm8051_golden_model_1.n1240 [281], RD_xram_29[1]);
  buf(\xm8051_golden_model_1.n1240 [282], RD_xram_29[2]);
  buf(\xm8051_golden_model_1.n1240 [283], RD_xram_29[3]);
  buf(\xm8051_golden_model_1.n1240 [284], RD_xram_29[4]);
  buf(\xm8051_golden_model_1.n1240 [285], RD_xram_29[5]);
  buf(\xm8051_golden_model_1.n1240 [286], RD_xram_29[6]);
  buf(\xm8051_golden_model_1.n1240 [287], RD_xram_29[7]);
  buf(\xm8051_golden_model_1.n1240 [288], RD_xram_28[0]);
  buf(\xm8051_golden_model_1.n1240 [289], RD_xram_28[1]);
  buf(\xm8051_golden_model_1.n1240 [290], RD_xram_28[2]);
  buf(\xm8051_golden_model_1.n1240 [291], RD_xram_28[3]);
  buf(\xm8051_golden_model_1.n1240 [292], RD_xram_28[4]);
  buf(\xm8051_golden_model_1.n1240 [293], RD_xram_28[5]);
  buf(\xm8051_golden_model_1.n1240 [294], RD_xram_28[6]);
  buf(\xm8051_golden_model_1.n1240 [295], RD_xram_28[7]);
  buf(\xm8051_golden_model_1.n1240 [296], RD_xram_27[0]);
  buf(\xm8051_golden_model_1.n1240 [297], RD_xram_27[1]);
  buf(\xm8051_golden_model_1.n1240 [298], RD_xram_27[2]);
  buf(\xm8051_golden_model_1.n1240 [299], RD_xram_27[3]);
  buf(\xm8051_golden_model_1.n1240 [300], RD_xram_27[4]);
  buf(\xm8051_golden_model_1.n1240 [301], RD_xram_27[5]);
  buf(\xm8051_golden_model_1.n1240 [302], RD_xram_27[6]);
  buf(\xm8051_golden_model_1.n1240 [303], RD_xram_27[7]);
  buf(\xm8051_golden_model_1.n1240 [304], RD_xram_26[0]);
  buf(\xm8051_golden_model_1.n1240 [305], RD_xram_26[1]);
  buf(\xm8051_golden_model_1.n1240 [306], RD_xram_26[2]);
  buf(\xm8051_golden_model_1.n1240 [307], RD_xram_26[3]);
  buf(\xm8051_golden_model_1.n1240 [308], RD_xram_26[4]);
  buf(\xm8051_golden_model_1.n1240 [309], RD_xram_26[5]);
  buf(\xm8051_golden_model_1.n1240 [310], RD_xram_26[6]);
  buf(\xm8051_golden_model_1.n1240 [311], RD_xram_26[7]);
  buf(\xm8051_golden_model_1.n1240 [312], RD_xram_25[0]);
  buf(\xm8051_golden_model_1.n1240 [313], RD_xram_25[1]);
  buf(\xm8051_golden_model_1.n1240 [314], RD_xram_25[2]);
  buf(\xm8051_golden_model_1.n1240 [315], RD_xram_25[3]);
  buf(\xm8051_golden_model_1.n1240 [316], RD_xram_25[4]);
  buf(\xm8051_golden_model_1.n1240 [317], RD_xram_25[5]);
  buf(\xm8051_golden_model_1.n1240 [318], RD_xram_25[6]);
  buf(\xm8051_golden_model_1.n1240 [319], RD_xram_25[7]);
  buf(\xm8051_golden_model_1.n1240 [320], RD_xram_24[0]);
  buf(\xm8051_golden_model_1.n1240 [321], RD_xram_24[1]);
  buf(\xm8051_golden_model_1.n1240 [322], RD_xram_24[2]);
  buf(\xm8051_golden_model_1.n1240 [323], RD_xram_24[3]);
  buf(\xm8051_golden_model_1.n1240 [324], RD_xram_24[4]);
  buf(\xm8051_golden_model_1.n1240 [325], RD_xram_24[5]);
  buf(\xm8051_golden_model_1.n1240 [326], RD_xram_24[6]);
  buf(\xm8051_golden_model_1.n1240 [327], RD_xram_24[7]);
  buf(\xm8051_golden_model_1.n1240 [328], RD_xram_23[0]);
  buf(\xm8051_golden_model_1.n1240 [329], RD_xram_23[1]);
  buf(\xm8051_golden_model_1.n1240 [330], RD_xram_23[2]);
  buf(\xm8051_golden_model_1.n1240 [331], RD_xram_23[3]);
  buf(\xm8051_golden_model_1.n1240 [332], RD_xram_23[4]);
  buf(\xm8051_golden_model_1.n1240 [333], RD_xram_23[5]);
  buf(\xm8051_golden_model_1.n1240 [334], RD_xram_23[6]);
  buf(\xm8051_golden_model_1.n1240 [335], RD_xram_23[7]);
  buf(\xm8051_golden_model_1.n1240 [336], RD_xram_22[0]);
  buf(\xm8051_golden_model_1.n1240 [337], RD_xram_22[1]);
  buf(\xm8051_golden_model_1.n1240 [338], RD_xram_22[2]);
  buf(\xm8051_golden_model_1.n1240 [339], RD_xram_22[3]);
  buf(\xm8051_golden_model_1.n1240 [340], RD_xram_22[4]);
  buf(\xm8051_golden_model_1.n1240 [341], RD_xram_22[5]);
  buf(\xm8051_golden_model_1.n1240 [342], RD_xram_22[6]);
  buf(\xm8051_golden_model_1.n1240 [343], RD_xram_22[7]);
  buf(\xm8051_golden_model_1.n1240 [344], RD_xram_21[0]);
  buf(\xm8051_golden_model_1.n1240 [345], RD_xram_21[1]);
  buf(\xm8051_golden_model_1.n1240 [346], RD_xram_21[2]);
  buf(\xm8051_golden_model_1.n1240 [347], RD_xram_21[3]);
  buf(\xm8051_golden_model_1.n1240 [348], RD_xram_21[4]);
  buf(\xm8051_golden_model_1.n1240 [349], RD_xram_21[5]);
  buf(\xm8051_golden_model_1.n1240 [350], RD_xram_21[6]);
  buf(\xm8051_golden_model_1.n1240 [351], RD_xram_21[7]);
  buf(\xm8051_golden_model_1.n1240 [352], RD_xram_20[0]);
  buf(\xm8051_golden_model_1.n1240 [353], RD_xram_20[1]);
  buf(\xm8051_golden_model_1.n1240 [354], RD_xram_20[2]);
  buf(\xm8051_golden_model_1.n1240 [355], RD_xram_20[3]);
  buf(\xm8051_golden_model_1.n1240 [356], RD_xram_20[4]);
  buf(\xm8051_golden_model_1.n1240 [357], RD_xram_20[5]);
  buf(\xm8051_golden_model_1.n1240 [358], RD_xram_20[6]);
  buf(\xm8051_golden_model_1.n1240 [359], RD_xram_20[7]);
  buf(\xm8051_golden_model_1.n1240 [360], RD_xram_19[0]);
  buf(\xm8051_golden_model_1.n1240 [361], RD_xram_19[1]);
  buf(\xm8051_golden_model_1.n1240 [362], RD_xram_19[2]);
  buf(\xm8051_golden_model_1.n1240 [363], RD_xram_19[3]);
  buf(\xm8051_golden_model_1.n1240 [364], RD_xram_19[4]);
  buf(\xm8051_golden_model_1.n1240 [365], RD_xram_19[5]);
  buf(\xm8051_golden_model_1.n1240 [366], RD_xram_19[6]);
  buf(\xm8051_golden_model_1.n1240 [367], RD_xram_19[7]);
  buf(\xm8051_golden_model_1.n1240 [368], RD_xram_18[0]);
  buf(\xm8051_golden_model_1.n1240 [369], RD_xram_18[1]);
  buf(\xm8051_golden_model_1.n1240 [370], RD_xram_18[2]);
  buf(\xm8051_golden_model_1.n1240 [371], RD_xram_18[3]);
  buf(\xm8051_golden_model_1.n1240 [372], RD_xram_18[4]);
  buf(\xm8051_golden_model_1.n1240 [373], RD_xram_18[5]);
  buf(\xm8051_golden_model_1.n1240 [374], RD_xram_18[6]);
  buf(\xm8051_golden_model_1.n1240 [375], RD_xram_18[7]);
  buf(\xm8051_golden_model_1.n1240 [376], RD_xram_17[0]);
  buf(\xm8051_golden_model_1.n1240 [377], RD_xram_17[1]);
  buf(\xm8051_golden_model_1.n1240 [378], RD_xram_17[2]);
  buf(\xm8051_golden_model_1.n1240 [379], RD_xram_17[3]);
  buf(\xm8051_golden_model_1.n1240 [380], RD_xram_17[4]);
  buf(\xm8051_golden_model_1.n1240 [381], RD_xram_17[5]);
  buf(\xm8051_golden_model_1.n1240 [382], RD_xram_17[6]);
  buf(\xm8051_golden_model_1.n1240 [383], RD_xram_17[7]);
  buf(\xm8051_golden_model_1.n1240 [384], RD_xram_16[0]);
  buf(\xm8051_golden_model_1.n1240 [385], RD_xram_16[1]);
  buf(\xm8051_golden_model_1.n1240 [386], RD_xram_16[2]);
  buf(\xm8051_golden_model_1.n1240 [387], RD_xram_16[3]);
  buf(\xm8051_golden_model_1.n1240 [388], RD_xram_16[4]);
  buf(\xm8051_golden_model_1.n1240 [389], RD_xram_16[5]);
  buf(\xm8051_golden_model_1.n1240 [390], RD_xram_16[6]);
  buf(\xm8051_golden_model_1.n1240 [391], RD_xram_16[7]);
  buf(\xm8051_golden_model_1.n1240 [392], RD_xram_15[0]);
  buf(\xm8051_golden_model_1.n1240 [393], RD_xram_15[1]);
  buf(\xm8051_golden_model_1.n1240 [394], RD_xram_15[2]);
  buf(\xm8051_golden_model_1.n1240 [395], RD_xram_15[3]);
  buf(\xm8051_golden_model_1.n1240 [396], RD_xram_15[4]);
  buf(\xm8051_golden_model_1.n1240 [397], RD_xram_15[5]);
  buf(\xm8051_golden_model_1.n1240 [398], RD_xram_15[6]);
  buf(\xm8051_golden_model_1.n1240 [399], RD_xram_15[7]);
  buf(\xm8051_golden_model_1.n1240 [400], RD_xram_14[0]);
  buf(\xm8051_golden_model_1.n1240 [401], RD_xram_14[1]);
  buf(\xm8051_golden_model_1.n1240 [402], RD_xram_14[2]);
  buf(\xm8051_golden_model_1.n1240 [403], RD_xram_14[3]);
  buf(\xm8051_golden_model_1.n1240 [404], RD_xram_14[4]);
  buf(\xm8051_golden_model_1.n1240 [405], RD_xram_14[5]);
  buf(\xm8051_golden_model_1.n1240 [406], RD_xram_14[6]);
  buf(\xm8051_golden_model_1.n1240 [407], RD_xram_14[7]);
  buf(\xm8051_golden_model_1.n1240 [408], RD_xram_13[0]);
  buf(\xm8051_golden_model_1.n1240 [409], RD_xram_13[1]);
  buf(\xm8051_golden_model_1.n1240 [410], RD_xram_13[2]);
  buf(\xm8051_golden_model_1.n1240 [411], RD_xram_13[3]);
  buf(\xm8051_golden_model_1.n1240 [412], RD_xram_13[4]);
  buf(\xm8051_golden_model_1.n1240 [413], RD_xram_13[5]);
  buf(\xm8051_golden_model_1.n1240 [414], RD_xram_13[6]);
  buf(\xm8051_golden_model_1.n1240 [415], RD_xram_13[7]);
  buf(\xm8051_golden_model_1.n1240 [416], RD_xram_12[0]);
  buf(\xm8051_golden_model_1.n1240 [417], RD_xram_12[1]);
  buf(\xm8051_golden_model_1.n1240 [418], RD_xram_12[2]);
  buf(\xm8051_golden_model_1.n1240 [419], RD_xram_12[3]);
  buf(\xm8051_golden_model_1.n1240 [420], RD_xram_12[4]);
  buf(\xm8051_golden_model_1.n1240 [421], RD_xram_12[5]);
  buf(\xm8051_golden_model_1.n1240 [422], RD_xram_12[6]);
  buf(\xm8051_golden_model_1.n1240 [423], RD_xram_12[7]);
  buf(\xm8051_golden_model_1.n1240 [424], RD_xram_11[0]);
  buf(\xm8051_golden_model_1.n1240 [425], RD_xram_11[1]);
  buf(\xm8051_golden_model_1.n1240 [426], RD_xram_11[2]);
  buf(\xm8051_golden_model_1.n1240 [427], RD_xram_11[3]);
  buf(\xm8051_golden_model_1.n1240 [428], RD_xram_11[4]);
  buf(\xm8051_golden_model_1.n1240 [429], RD_xram_11[5]);
  buf(\xm8051_golden_model_1.n1240 [430], RD_xram_11[6]);
  buf(\xm8051_golden_model_1.n1240 [431], RD_xram_11[7]);
  buf(\xm8051_golden_model_1.n1240 [432], RD_xram_10[0]);
  buf(\xm8051_golden_model_1.n1240 [433], RD_xram_10[1]);
  buf(\xm8051_golden_model_1.n1240 [434], RD_xram_10[2]);
  buf(\xm8051_golden_model_1.n1240 [435], RD_xram_10[3]);
  buf(\xm8051_golden_model_1.n1240 [436], RD_xram_10[4]);
  buf(\xm8051_golden_model_1.n1240 [437], RD_xram_10[5]);
  buf(\xm8051_golden_model_1.n1240 [438], RD_xram_10[6]);
  buf(\xm8051_golden_model_1.n1240 [439], RD_xram_10[7]);
  buf(\xm8051_golden_model_1.n1240 [440], RD_xram_9[0]);
  buf(\xm8051_golden_model_1.n1240 [441], RD_xram_9[1]);
  buf(\xm8051_golden_model_1.n1240 [442], RD_xram_9[2]);
  buf(\xm8051_golden_model_1.n1240 [443], RD_xram_9[3]);
  buf(\xm8051_golden_model_1.n1240 [444], RD_xram_9[4]);
  buf(\xm8051_golden_model_1.n1240 [445], RD_xram_9[5]);
  buf(\xm8051_golden_model_1.n1240 [446], RD_xram_9[6]);
  buf(\xm8051_golden_model_1.n1240 [447], RD_xram_9[7]);
  buf(\xm8051_golden_model_1.n1240 [448], RD_xram_8[0]);
  buf(\xm8051_golden_model_1.n1240 [449], RD_xram_8[1]);
  buf(\xm8051_golden_model_1.n1240 [450], RD_xram_8[2]);
  buf(\xm8051_golden_model_1.n1240 [451], RD_xram_8[3]);
  buf(\xm8051_golden_model_1.n1240 [452], RD_xram_8[4]);
  buf(\xm8051_golden_model_1.n1240 [453], RD_xram_8[5]);
  buf(\xm8051_golden_model_1.n1240 [454], RD_xram_8[6]);
  buf(\xm8051_golden_model_1.n1240 [455], RD_xram_8[7]);
  buf(\xm8051_golden_model_1.n1240 [456], RD_xram_7[0]);
  buf(\xm8051_golden_model_1.n1240 [457], RD_xram_7[1]);
  buf(\xm8051_golden_model_1.n1240 [458], RD_xram_7[2]);
  buf(\xm8051_golden_model_1.n1240 [459], RD_xram_7[3]);
  buf(\xm8051_golden_model_1.n1240 [460], RD_xram_7[4]);
  buf(\xm8051_golden_model_1.n1240 [461], RD_xram_7[5]);
  buf(\xm8051_golden_model_1.n1240 [462], RD_xram_7[6]);
  buf(\xm8051_golden_model_1.n1240 [463], RD_xram_7[7]);
  buf(\xm8051_golden_model_1.n1240 [464], RD_xram_6[0]);
  buf(\xm8051_golden_model_1.n1240 [465], RD_xram_6[1]);
  buf(\xm8051_golden_model_1.n1240 [466], RD_xram_6[2]);
  buf(\xm8051_golden_model_1.n1240 [467], RD_xram_6[3]);
  buf(\xm8051_golden_model_1.n1240 [468], RD_xram_6[4]);
  buf(\xm8051_golden_model_1.n1240 [469], RD_xram_6[5]);
  buf(\xm8051_golden_model_1.n1240 [470], RD_xram_6[6]);
  buf(\xm8051_golden_model_1.n1240 [471], RD_xram_6[7]);
  buf(\xm8051_golden_model_1.n1240 [472], RD_xram_5[0]);
  buf(\xm8051_golden_model_1.n1240 [473], RD_xram_5[1]);
  buf(\xm8051_golden_model_1.n1240 [474], RD_xram_5[2]);
  buf(\xm8051_golden_model_1.n1240 [475], RD_xram_5[3]);
  buf(\xm8051_golden_model_1.n1240 [476], RD_xram_5[4]);
  buf(\xm8051_golden_model_1.n1240 [477], RD_xram_5[5]);
  buf(\xm8051_golden_model_1.n1240 [478], RD_xram_5[6]);
  buf(\xm8051_golden_model_1.n1240 [479], RD_xram_5[7]);
  buf(\xm8051_golden_model_1.n1240 [480], RD_xram_4[0]);
  buf(\xm8051_golden_model_1.n1240 [481], RD_xram_4[1]);
  buf(\xm8051_golden_model_1.n1240 [482], RD_xram_4[2]);
  buf(\xm8051_golden_model_1.n1240 [483], RD_xram_4[3]);
  buf(\xm8051_golden_model_1.n1240 [484], RD_xram_4[4]);
  buf(\xm8051_golden_model_1.n1240 [485], RD_xram_4[5]);
  buf(\xm8051_golden_model_1.n1240 [486], RD_xram_4[6]);
  buf(\xm8051_golden_model_1.n1240 [487], RD_xram_4[7]);
  buf(\xm8051_golden_model_1.n1240 [488], RD_xram_3[0]);
  buf(\xm8051_golden_model_1.n1240 [489], RD_xram_3[1]);
  buf(\xm8051_golden_model_1.n1240 [490], RD_xram_3[2]);
  buf(\xm8051_golden_model_1.n1240 [491], RD_xram_3[3]);
  buf(\xm8051_golden_model_1.n1240 [492], RD_xram_3[4]);
  buf(\xm8051_golden_model_1.n1240 [493], RD_xram_3[5]);
  buf(\xm8051_golden_model_1.n1240 [494], RD_xram_3[6]);
  buf(\xm8051_golden_model_1.n1240 [495], RD_xram_3[7]);
  buf(\xm8051_golden_model_1.n1240 [496], RD_xram_2[0]);
  buf(\xm8051_golden_model_1.n1240 [497], RD_xram_2[1]);
  buf(\xm8051_golden_model_1.n1240 [498], RD_xram_2[2]);
  buf(\xm8051_golden_model_1.n1240 [499], RD_xram_2[3]);
  buf(\xm8051_golden_model_1.n1240 [500], RD_xram_2[4]);
  buf(\xm8051_golden_model_1.n1240 [501], RD_xram_2[5]);
  buf(\xm8051_golden_model_1.n1240 [502], RD_xram_2[6]);
  buf(\xm8051_golden_model_1.n1240 [503], RD_xram_2[7]);
  buf(\xm8051_golden_model_1.n1240 [504], RD_xram_1[0]);
  buf(\xm8051_golden_model_1.n1240 [505], RD_xram_1[1]);
  buf(\xm8051_golden_model_1.n1240 [506], RD_xram_1[2]);
  buf(\xm8051_golden_model_1.n1240 [507], RD_xram_1[3]);
  buf(\xm8051_golden_model_1.n1240 [508], RD_xram_1[4]);
  buf(\xm8051_golden_model_1.n1240 [509], RD_xram_1[5]);
  buf(\xm8051_golden_model_1.n1240 [510], RD_xram_1[6]);
  buf(\xm8051_golden_model_1.n1240 [511], RD_xram_1[7]);
  buf(\xm8051_golden_model_1.n1236 [0], input_sha_func_16[0]);
  buf(\xm8051_golden_model_1.n1236 [1], input_sha_func_16[1]);
  buf(\xm8051_golden_model_1.n1236 [2], input_sha_func_16[2]);
  buf(\xm8051_golden_model_1.n1236 [3], input_sha_func_16[3]);
  buf(\xm8051_golden_model_1.n1236 [4], input_sha_func_16[4]);
  buf(\xm8051_golden_model_1.n1236 [5], input_sha_func_16[5]);
  buf(\xm8051_golden_model_1.n1236 [6], input_sha_func_16[6]);
  buf(\xm8051_golden_model_1.n1236 [7], input_sha_func_16[7]);
  buf(\xm8051_golden_model_1.n1236 [8], input_sha_func_16[8]);
  buf(\xm8051_golden_model_1.n1236 [9], input_sha_func_16[9]);
  buf(\xm8051_golden_model_1.n1236 [10], input_sha_func_16[10]);
  buf(\xm8051_golden_model_1.n1236 [11], input_sha_func_16[11]);
  buf(\xm8051_golden_model_1.n1236 [12], input_sha_func_16[12]);
  buf(\xm8051_golden_model_1.n1236 [13], input_sha_func_16[13]);
  buf(\xm8051_golden_model_1.n1236 [14], input_sha_func_16[14]);
  buf(\xm8051_golden_model_1.n1236 [15], input_sha_func_16[15]);
  buf(\xm8051_golden_model_1.n1236 [16], input_sha_func_16[16]);
  buf(\xm8051_golden_model_1.n1236 [17], input_sha_func_16[17]);
  buf(\xm8051_golden_model_1.n1236 [18], input_sha_func_16[18]);
  buf(\xm8051_golden_model_1.n1236 [19], input_sha_func_16[19]);
  buf(\xm8051_golden_model_1.n1236 [20], input_sha_func_16[20]);
  buf(\xm8051_golden_model_1.n1236 [21], input_sha_func_16[21]);
  buf(\xm8051_golden_model_1.n1236 [22], input_sha_func_16[22]);
  buf(\xm8051_golden_model_1.n1236 [23], input_sha_func_16[23]);
  buf(\xm8051_golden_model_1.n1236 [24], input_sha_func_16[24]);
  buf(\xm8051_golden_model_1.n1236 [25], input_sha_func_16[25]);
  buf(\xm8051_golden_model_1.n1236 [26], input_sha_func_16[26]);
  buf(\xm8051_golden_model_1.n1236 [27], input_sha_func_16[27]);
  buf(\xm8051_golden_model_1.n1236 [28], input_sha_func_16[28]);
  buf(\xm8051_golden_model_1.n1236 [29], input_sha_func_16[29]);
  buf(\xm8051_golden_model_1.n1236 [30], input_sha_func_16[30]);
  buf(\xm8051_golden_model_1.n1236 [31], input_sha_func_16[31]);
  buf(\xm8051_golden_model_1.n1236 [32], input_sha_func_15[0]);
  buf(\xm8051_golden_model_1.n1236 [33], input_sha_func_15[1]);
  buf(\xm8051_golden_model_1.n1236 [34], input_sha_func_15[2]);
  buf(\xm8051_golden_model_1.n1236 [35], input_sha_func_15[3]);
  buf(\xm8051_golden_model_1.n1236 [36], input_sha_func_15[4]);
  buf(\xm8051_golden_model_1.n1236 [37], input_sha_func_15[5]);
  buf(\xm8051_golden_model_1.n1236 [38], input_sha_func_15[6]);
  buf(\xm8051_golden_model_1.n1236 [39], input_sha_func_15[7]);
  buf(\xm8051_golden_model_1.n1236 [40], input_sha_func_15[8]);
  buf(\xm8051_golden_model_1.n1236 [41], input_sha_func_15[9]);
  buf(\xm8051_golden_model_1.n1236 [42], input_sha_func_15[10]);
  buf(\xm8051_golden_model_1.n1236 [43], input_sha_func_15[11]);
  buf(\xm8051_golden_model_1.n1236 [44], input_sha_func_15[12]);
  buf(\xm8051_golden_model_1.n1236 [45], input_sha_func_15[13]);
  buf(\xm8051_golden_model_1.n1236 [46], input_sha_func_15[14]);
  buf(\xm8051_golden_model_1.n1236 [47], input_sha_func_15[15]);
  buf(\xm8051_golden_model_1.n1236 [48], input_sha_func_15[16]);
  buf(\xm8051_golden_model_1.n1236 [49], input_sha_func_15[17]);
  buf(\xm8051_golden_model_1.n1236 [50], input_sha_func_15[18]);
  buf(\xm8051_golden_model_1.n1236 [51], input_sha_func_15[19]);
  buf(\xm8051_golden_model_1.n1236 [52], input_sha_func_15[20]);
  buf(\xm8051_golden_model_1.n1236 [53], input_sha_func_15[21]);
  buf(\xm8051_golden_model_1.n1236 [54], input_sha_func_15[22]);
  buf(\xm8051_golden_model_1.n1236 [55], input_sha_func_15[23]);
  buf(\xm8051_golden_model_1.n1236 [56], input_sha_func_15[24]);
  buf(\xm8051_golden_model_1.n1236 [57], input_sha_func_15[25]);
  buf(\xm8051_golden_model_1.n1236 [58], input_sha_func_15[26]);
  buf(\xm8051_golden_model_1.n1236 [59], input_sha_func_15[27]);
  buf(\xm8051_golden_model_1.n1236 [60], input_sha_func_15[28]);
  buf(\xm8051_golden_model_1.n1236 [61], input_sha_func_15[29]);
  buf(\xm8051_golden_model_1.n1236 [62], input_sha_func_15[30]);
  buf(\xm8051_golden_model_1.n1236 [63], input_sha_func_15[31]);
  buf(\xm8051_golden_model_1.n1236 [64], input_sha_func_15[32]);
  buf(\xm8051_golden_model_1.n1236 [65], input_sha_func_15[33]);
  buf(\xm8051_golden_model_1.n1236 [66], input_sha_func_15[34]);
  buf(\xm8051_golden_model_1.n1236 [67], input_sha_func_15[35]);
  buf(\xm8051_golden_model_1.n1236 [68], input_sha_func_15[36]);
  buf(\xm8051_golden_model_1.n1236 [69], input_sha_func_15[37]);
  buf(\xm8051_golden_model_1.n1236 [70], input_sha_func_15[38]);
  buf(\xm8051_golden_model_1.n1236 [71], input_sha_func_15[39]);
  buf(\xm8051_golden_model_1.n1236 [72], input_sha_func_15[40]);
  buf(\xm8051_golden_model_1.n1236 [73], input_sha_func_15[41]);
  buf(\xm8051_golden_model_1.n1236 [74], input_sha_func_15[42]);
  buf(\xm8051_golden_model_1.n1236 [75], input_sha_func_15[43]);
  buf(\xm8051_golden_model_1.n1236 [76], input_sha_func_15[44]);
  buf(\xm8051_golden_model_1.n1236 [77], input_sha_func_15[45]);
  buf(\xm8051_golden_model_1.n1236 [78], input_sha_func_15[46]);
  buf(\xm8051_golden_model_1.n1236 [79], input_sha_func_15[47]);
  buf(\xm8051_golden_model_1.n1236 [80], input_sha_func_15[48]);
  buf(\xm8051_golden_model_1.n1236 [81], input_sha_func_15[49]);
  buf(\xm8051_golden_model_1.n1236 [82], input_sha_func_15[50]);
  buf(\xm8051_golden_model_1.n1236 [83], input_sha_func_15[51]);
  buf(\xm8051_golden_model_1.n1236 [84], input_sha_func_15[52]);
  buf(\xm8051_golden_model_1.n1236 [85], input_sha_func_15[53]);
  buf(\xm8051_golden_model_1.n1236 [86], input_sha_func_15[54]);
  buf(\xm8051_golden_model_1.n1236 [87], input_sha_func_15[55]);
  buf(\xm8051_golden_model_1.n1236 [88], input_sha_func_15[56]);
  buf(\xm8051_golden_model_1.n1236 [89], input_sha_func_15[57]);
  buf(\xm8051_golden_model_1.n1236 [90], input_sha_func_15[58]);
  buf(\xm8051_golden_model_1.n1236 [91], input_sha_func_15[59]);
  buf(\xm8051_golden_model_1.n1236 [92], input_sha_func_15[60]);
  buf(\xm8051_golden_model_1.n1236 [93], input_sha_func_15[61]);
  buf(\xm8051_golden_model_1.n1236 [94], input_sha_func_15[62]);
  buf(\xm8051_golden_model_1.n1236 [95], input_sha_func_15[63]);
  buf(\xm8051_golden_model_1.n1236 [96], input_sha_func_14[0]);
  buf(\xm8051_golden_model_1.n1236 [97], input_sha_func_14[1]);
  buf(\xm8051_golden_model_1.n1236 [98], input_sha_func_14[2]);
  buf(\xm8051_golden_model_1.n1236 [99], input_sha_func_14[3]);
  buf(\xm8051_golden_model_1.n1236 [100], input_sha_func_14[4]);
  buf(\xm8051_golden_model_1.n1236 [101], input_sha_func_14[5]);
  buf(\xm8051_golden_model_1.n1236 [102], input_sha_func_14[6]);
  buf(\xm8051_golden_model_1.n1236 [103], input_sha_func_14[7]);
  buf(\xm8051_golden_model_1.n1236 [104], input_sha_func_14[8]);
  buf(\xm8051_golden_model_1.n1236 [105], input_sha_func_14[9]);
  buf(\xm8051_golden_model_1.n1236 [106], input_sha_func_14[10]);
  buf(\xm8051_golden_model_1.n1236 [107], input_sha_func_14[11]);
  buf(\xm8051_golden_model_1.n1236 [108], input_sha_func_14[12]);
  buf(\xm8051_golden_model_1.n1236 [109], input_sha_func_14[13]);
  buf(\xm8051_golden_model_1.n1236 [110], input_sha_func_14[14]);
  buf(\xm8051_golden_model_1.n1236 [111], input_sha_func_14[15]);
  buf(\xm8051_golden_model_1.n1236 [112], input_sha_func_14[16]);
  buf(\xm8051_golden_model_1.n1236 [113], input_sha_func_14[17]);
  buf(\xm8051_golden_model_1.n1236 [114], input_sha_func_14[18]);
  buf(\xm8051_golden_model_1.n1236 [115], input_sha_func_14[19]);
  buf(\xm8051_golden_model_1.n1236 [116], input_sha_func_14[20]);
  buf(\xm8051_golden_model_1.n1236 [117], input_sha_func_14[21]);
  buf(\xm8051_golden_model_1.n1236 [118], input_sha_func_14[22]);
  buf(\xm8051_golden_model_1.n1236 [119], input_sha_func_14[23]);
  buf(\xm8051_golden_model_1.n1236 [120], input_sha_func_14[24]);
  buf(\xm8051_golden_model_1.n1236 [121], input_sha_func_14[25]);
  buf(\xm8051_golden_model_1.n1236 [122], input_sha_func_14[26]);
  buf(\xm8051_golden_model_1.n1236 [123], input_sha_func_14[27]);
  buf(\xm8051_golden_model_1.n1236 [124], input_sha_func_14[28]);
  buf(\xm8051_golden_model_1.n1236 [125], input_sha_func_14[29]);
  buf(\xm8051_golden_model_1.n1236 [126], input_sha_func_14[30]);
  buf(\xm8051_golden_model_1.n1236 [127], input_sha_func_14[31]);
  buf(\xm8051_golden_model_1.n1236 [128], input_sha_func_14[32]);
  buf(\xm8051_golden_model_1.n1236 [129], input_sha_func_14[33]);
  buf(\xm8051_golden_model_1.n1236 [130], input_sha_func_14[34]);
  buf(\xm8051_golden_model_1.n1236 [131], input_sha_func_14[35]);
  buf(\xm8051_golden_model_1.n1236 [132], input_sha_func_14[36]);
  buf(\xm8051_golden_model_1.n1236 [133], input_sha_func_14[37]);
  buf(\xm8051_golden_model_1.n1236 [134], input_sha_func_14[38]);
  buf(\xm8051_golden_model_1.n1236 [135], input_sha_func_14[39]);
  buf(\xm8051_golden_model_1.n1236 [136], input_sha_func_14[40]);
  buf(\xm8051_golden_model_1.n1236 [137], input_sha_func_14[41]);
  buf(\xm8051_golden_model_1.n1236 [138], input_sha_func_14[42]);
  buf(\xm8051_golden_model_1.n1236 [139], input_sha_func_14[43]);
  buf(\xm8051_golden_model_1.n1236 [140], input_sha_func_14[44]);
  buf(\xm8051_golden_model_1.n1236 [141], input_sha_func_14[45]);
  buf(\xm8051_golden_model_1.n1236 [142], input_sha_func_14[46]);
  buf(\xm8051_golden_model_1.n1236 [143], input_sha_func_14[47]);
  buf(\xm8051_golden_model_1.n1236 [144], input_sha_func_14[48]);
  buf(\xm8051_golden_model_1.n1236 [145], input_sha_func_14[49]);
  buf(\xm8051_golden_model_1.n1236 [146], input_sha_func_14[50]);
  buf(\xm8051_golden_model_1.n1236 [147], input_sha_func_14[51]);
  buf(\xm8051_golden_model_1.n1236 [148], input_sha_func_14[52]);
  buf(\xm8051_golden_model_1.n1236 [149], input_sha_func_14[53]);
  buf(\xm8051_golden_model_1.n1236 [150], input_sha_func_14[54]);
  buf(\xm8051_golden_model_1.n1236 [151], input_sha_func_14[55]);
  buf(\xm8051_golden_model_1.n1236 [152], input_sha_func_14[56]);
  buf(\xm8051_golden_model_1.n1236 [153], input_sha_func_14[57]);
  buf(\xm8051_golden_model_1.n1236 [154], input_sha_func_14[58]);
  buf(\xm8051_golden_model_1.n1236 [155], input_sha_func_14[59]);
  buf(\xm8051_golden_model_1.n1236 [156], input_sha_func_14[60]);
  buf(\xm8051_golden_model_1.n1236 [157], input_sha_func_14[61]);
  buf(\xm8051_golden_model_1.n1236 [158], input_sha_func_14[62]);
  buf(\xm8051_golden_model_1.n1236 [159], input_sha_func_14[63]);
  buf(\xm8051_golden_model_1.n0196 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0196 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0196 [2], \xm8051_golden_model_1.n0483 [2]);
  buf(\xm8051_golden_model_1.n0196 [3], \xm8051_golden_model_1.n0483 [3]);
  buf(\xm8051_golden_model_1.n0196 [4], \xm8051_golden_model_1.n0401 [4]);
  buf(\xm8051_golden_model_1.n0187 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0174 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0174 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0174 [2], \xm8051_golden_model_1.n0473 [2]);
  buf(\xm8051_golden_model_1.n0174 [3], \xm8051_golden_model_1.n0473 [3]);
  buf(\xm8051_golden_model_1.n0174 [4], \xm8051_golden_model_1.n0389 [4]);
  buf(\xm8051_golden_model_1.n0165 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0165 [1], \xm8051_golden_model_1.aes_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0152 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0152 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0152 [2], \xm8051_golden_model_1.n0463 [2]);
  buf(\xm8051_golden_model_1.n0152 [3], \xm8051_golden_model_1.n0463 [3]);
  buf(\xm8051_golden_model_1.n0152 [4], \xm8051_golden_model_1.n0377 [4]);
  buf(\xm8051_golden_model_1.n0143 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0143 [1], \xm8051_golden_model_1.n0187 [1]);
  buf(\xm8051_golden_model_1.n0130 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0130 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0130 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n0130 [3], \xm8051_golden_model_1.n0453 [3]);
  buf(\xm8051_golden_model_1.n0130 [4], \xm8051_golden_model_1.n0365 [4]);
  buf(\xm8051_golden_model_1.n0121 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0121 [1], \xm8051_golden_model_1.aes_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0121 [2], \xm8051_golden_model_1.aes_bytes_processed [2]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0b [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0b [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0b [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0b [3], \xm8051_golden_model_1.sha_bytes_processed [3]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0b [4], \xm8051_golden_model_1.sha_bytes_processed [4]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0b [5], \xm8051_golden_model_1.sha_bytes_processed [5]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [3], \xm8051_golden_model_1.sha_bytes_processed [3]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [4], \xm8051_golden_model_1.sha_bytes_processed [4]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [5], \xm8051_golden_model_1.sha_bytes_processed [5]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [6], \xm8051_golden_model_1.sha_bytes_processed_0b [6]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [7], \xm8051_golden_model_1.sha_bytes_processed_0b [7]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [8], \xm8051_golden_model_1.sha_bytes_processed_0b [8]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [9], \xm8051_golden_model_1.sha_bytes_processed_0b [9]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [10], \xm8051_golden_model_1.sha_bytes_processed_0b [10]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [11], \xm8051_golden_model_1.sha_bytes_processed_0b [11]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [12], \xm8051_golden_model_1.sha_bytes_processed_0b [12]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [13], \xm8051_golden_model_1.sha_bytes_processed_0b [13]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [14], \xm8051_golden_model_1.sha_bytes_processed_0b [14]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_0a [15], \xm8051_golden_model_1.sha_bytes_processed_0b [15]);
  buf(\xm8051_golden_model_1.n0108 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0108 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0108 [2], \xm8051_golden_model_1.n0483 [2]);
  buf(\xm8051_golden_model_1.n0108 [3], \xm8051_golden_model_1.n0443 [3]);
  buf(\xm8051_golden_model_1.n0108 [4], \xm8051_golden_model_1.n0353 [4]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [3], \xm8051_golden_model_1.sha_bytes_processed [3]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [4], \xm8051_golden_model_1.sha_bytes_processed [4]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [5], \xm8051_golden_model_1.sha_bytes_processed [5]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [6], \xm8051_golden_model_1.sha_bytes_processed_0b [6]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [7], \xm8051_golden_model_1.sha_bytes_processed_0b [7]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [8], \xm8051_golden_model_1.sha_bytes_processed_0b [8]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [9], \xm8051_golden_model_1.sha_bytes_processed_0b [9]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [10], \xm8051_golden_model_1.sha_bytes_processed_0b [10]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [11], \xm8051_golden_model_1.sha_bytes_processed_0b [11]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [12], \xm8051_golden_model_1.sha_bytes_processed_0b [12]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [13], \xm8051_golden_model_1.sha_bytes_processed_0b [13]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [14], \xm8051_golden_model_1.sha_bytes_processed_0b [14]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_09 [15], \xm8051_golden_model_1.sha_bytes_processed_0b [15]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [3], \xm8051_golden_model_1.sha_bytes_processed [3]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [4], \xm8051_golden_model_1.sha_bytes_processed [4]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [5], \xm8051_golden_model_1.sha_bytes_processed [5]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [6], \xm8051_golden_model_1.sha_bytes_processed_0b [6]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [7], \xm8051_golden_model_1.sha_bytes_processed_0b [7]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [8], \xm8051_golden_model_1.sha_bytes_processed_0b [8]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [9], \xm8051_golden_model_1.sha_bytes_processed_0b [9]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [10], \xm8051_golden_model_1.sha_bytes_processed_0b [10]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [11], \xm8051_golden_model_1.sha_bytes_processed_0b [11]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [12], \xm8051_golden_model_1.sha_bytes_processed_0b [12]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [13], \xm8051_golden_model_1.sha_bytes_processed_0b [13]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [14], \xm8051_golden_model_1.sha_bytes_processed_0b [14]);
  buf(\xm8051_golden_model_1.sha_bytes_processed_08 [15], \xm8051_golden_model_1.sha_bytes_processed_0b [15]);
  buf(\xm8051_golden_model_1.n0983 [0], input_sha_func_13[0]);
  buf(\xm8051_golden_model_1.n0983 [1], input_sha_func_13[1]);
  buf(\xm8051_golden_model_1.n0983 [2], input_sha_func_13[2]);
  buf(\xm8051_golden_model_1.n0983 [3], input_sha_func_13[3]);
  buf(\xm8051_golden_model_1.n0983 [4], input_sha_func_13[4]);
  buf(\xm8051_golden_model_1.n0983 [5], input_sha_func_13[5]);
  buf(\xm8051_golden_model_1.n0983 [6], input_sha_func_13[6]);
  buf(\xm8051_golden_model_1.n0983 [7], input_sha_func_13[7]);
  buf(\xm8051_golden_model_1.n0983 [8], input_sha_func_13[8]);
  buf(\xm8051_golden_model_1.n0983 [9], input_sha_func_13[9]);
  buf(\xm8051_golden_model_1.n0983 [10], input_sha_func_13[10]);
  buf(\xm8051_golden_model_1.n0983 [11], input_sha_func_13[11]);
  buf(\xm8051_golden_model_1.n0983 [12], input_sha_func_13[12]);
  buf(\xm8051_golden_model_1.n0983 [13], input_sha_func_13[13]);
  buf(\xm8051_golden_model_1.n0983 [14], input_sha_func_13[14]);
  buf(\xm8051_golden_model_1.n0983 [15], input_sha_func_13[15]);
  buf(\xm8051_golden_model_1.n0983 [16], input_sha_func_13[16]);
  buf(\xm8051_golden_model_1.n0983 [17], input_sha_func_13[17]);
  buf(\xm8051_golden_model_1.n0983 [18], input_sha_func_13[18]);
  buf(\xm8051_golden_model_1.n0983 [19], input_sha_func_13[19]);
  buf(\xm8051_golden_model_1.n0983 [20], input_sha_func_13[20]);
  buf(\xm8051_golden_model_1.n0983 [21], input_sha_func_13[21]);
  buf(\xm8051_golden_model_1.n0983 [22], input_sha_func_13[22]);
  buf(\xm8051_golden_model_1.n0983 [23], input_sha_func_13[23]);
  buf(\xm8051_golden_model_1.n0983 [24], input_sha_func_13[24]);
  buf(\xm8051_golden_model_1.n0983 [25], input_sha_func_13[25]);
  buf(\xm8051_golden_model_1.n0983 [26], input_sha_func_13[26]);
  buf(\xm8051_golden_model_1.n0983 [27], input_sha_func_13[27]);
  buf(\xm8051_golden_model_1.n0983 [28], input_sha_func_13[28]);
  buf(\xm8051_golden_model_1.n0983 [29], input_sha_func_13[29]);
  buf(\xm8051_golden_model_1.n0983 [30], input_sha_func_13[30]);
  buf(\xm8051_golden_model_1.n0983 [31], input_sha_func_13[31]);
  buf(\xm8051_golden_model_1.n0983 [32], input_sha_func_12[0]);
  buf(\xm8051_golden_model_1.n0983 [33], input_sha_func_12[1]);
  buf(\xm8051_golden_model_1.n0983 [34], input_sha_func_12[2]);
  buf(\xm8051_golden_model_1.n0983 [35], input_sha_func_12[3]);
  buf(\xm8051_golden_model_1.n0983 [36], input_sha_func_12[4]);
  buf(\xm8051_golden_model_1.n0983 [37], input_sha_func_12[5]);
  buf(\xm8051_golden_model_1.n0983 [38], input_sha_func_12[6]);
  buf(\xm8051_golden_model_1.n0983 [39], input_sha_func_12[7]);
  buf(\xm8051_golden_model_1.n0983 [40], input_sha_func_12[8]);
  buf(\xm8051_golden_model_1.n0983 [41], input_sha_func_12[9]);
  buf(\xm8051_golden_model_1.n0983 [42], input_sha_func_12[10]);
  buf(\xm8051_golden_model_1.n0983 [43], input_sha_func_12[11]);
  buf(\xm8051_golden_model_1.n0983 [44], input_sha_func_12[12]);
  buf(\xm8051_golden_model_1.n0983 [45], input_sha_func_12[13]);
  buf(\xm8051_golden_model_1.n0983 [46], input_sha_func_12[14]);
  buf(\xm8051_golden_model_1.n0983 [47], input_sha_func_12[15]);
  buf(\xm8051_golden_model_1.n0983 [48], input_sha_func_12[16]);
  buf(\xm8051_golden_model_1.n0983 [49], input_sha_func_12[17]);
  buf(\xm8051_golden_model_1.n0983 [50], input_sha_func_12[18]);
  buf(\xm8051_golden_model_1.n0983 [51], input_sha_func_12[19]);
  buf(\xm8051_golden_model_1.n0983 [52], input_sha_func_12[20]);
  buf(\xm8051_golden_model_1.n0983 [53], input_sha_func_12[21]);
  buf(\xm8051_golden_model_1.n0983 [54], input_sha_func_12[22]);
  buf(\xm8051_golden_model_1.n0983 [55], input_sha_func_12[23]);
  buf(\xm8051_golden_model_1.n0983 [56], input_sha_func_12[24]);
  buf(\xm8051_golden_model_1.n0983 [57], input_sha_func_12[25]);
  buf(\xm8051_golden_model_1.n0983 [58], input_sha_func_12[26]);
  buf(\xm8051_golden_model_1.n0983 [59], input_sha_func_12[27]);
  buf(\xm8051_golden_model_1.n0983 [60], input_sha_func_12[28]);
  buf(\xm8051_golden_model_1.n0983 [61], input_sha_func_12[29]);
  buf(\xm8051_golden_model_1.n0983 [62], input_sha_func_12[30]);
  buf(\xm8051_golden_model_1.n0983 [63], input_sha_func_12[31]);
  buf(\xm8051_golden_model_1.n0983 [64], input_sha_func_12[32]);
  buf(\xm8051_golden_model_1.n0983 [65], input_sha_func_12[33]);
  buf(\xm8051_golden_model_1.n0983 [66], input_sha_func_12[34]);
  buf(\xm8051_golden_model_1.n0983 [67], input_sha_func_12[35]);
  buf(\xm8051_golden_model_1.n0983 [68], input_sha_func_12[36]);
  buf(\xm8051_golden_model_1.n0983 [69], input_sha_func_12[37]);
  buf(\xm8051_golden_model_1.n0983 [70], input_sha_func_12[38]);
  buf(\xm8051_golden_model_1.n0983 [71], input_sha_func_12[39]);
  buf(\xm8051_golden_model_1.n0983 [72], input_sha_func_12[40]);
  buf(\xm8051_golden_model_1.n0983 [73], input_sha_func_12[41]);
  buf(\xm8051_golden_model_1.n0983 [74], input_sha_func_12[42]);
  buf(\xm8051_golden_model_1.n0983 [75], input_sha_func_12[43]);
  buf(\xm8051_golden_model_1.n0983 [76], input_sha_func_12[44]);
  buf(\xm8051_golden_model_1.n0983 [77], input_sha_func_12[45]);
  buf(\xm8051_golden_model_1.n0983 [78], input_sha_func_12[46]);
  buf(\xm8051_golden_model_1.n0983 [79], input_sha_func_12[47]);
  buf(\xm8051_golden_model_1.n0983 [80], input_sha_func_12[48]);
  buf(\xm8051_golden_model_1.n0983 [81], input_sha_func_12[49]);
  buf(\xm8051_golden_model_1.n0983 [82], input_sha_func_12[50]);
  buf(\xm8051_golden_model_1.n0983 [83], input_sha_func_12[51]);
  buf(\xm8051_golden_model_1.n0983 [84], input_sha_func_12[52]);
  buf(\xm8051_golden_model_1.n0983 [85], input_sha_func_12[53]);
  buf(\xm8051_golden_model_1.n0983 [86], input_sha_func_12[54]);
  buf(\xm8051_golden_model_1.n0983 [87], input_sha_func_12[55]);
  buf(\xm8051_golden_model_1.n0983 [88], input_sha_func_12[56]);
  buf(\xm8051_golden_model_1.n0983 [89], input_sha_func_12[57]);
  buf(\xm8051_golden_model_1.n0983 [90], input_sha_func_12[58]);
  buf(\xm8051_golden_model_1.n0983 [91], input_sha_func_12[59]);
  buf(\xm8051_golden_model_1.n0983 [92], input_sha_func_12[60]);
  buf(\xm8051_golden_model_1.n0983 [93], input_sha_func_12[61]);
  buf(\xm8051_golden_model_1.n0983 [94], input_sha_func_12[62]);
  buf(\xm8051_golden_model_1.n0983 [95], input_sha_func_12[63]);
  buf(\xm8051_golden_model_1.n0983 [96], input_sha_func_11[0]);
  buf(\xm8051_golden_model_1.n0983 [97], input_sha_func_11[1]);
  buf(\xm8051_golden_model_1.n0983 [98], input_sha_func_11[2]);
  buf(\xm8051_golden_model_1.n0983 [99], input_sha_func_11[3]);
  buf(\xm8051_golden_model_1.n0983 [100], input_sha_func_11[4]);
  buf(\xm8051_golden_model_1.n0983 [101], input_sha_func_11[5]);
  buf(\xm8051_golden_model_1.n0983 [102], input_sha_func_11[6]);
  buf(\xm8051_golden_model_1.n0983 [103], input_sha_func_11[7]);
  buf(\xm8051_golden_model_1.n0983 [104], input_sha_func_11[8]);
  buf(\xm8051_golden_model_1.n0983 [105], input_sha_func_11[9]);
  buf(\xm8051_golden_model_1.n0983 [106], input_sha_func_11[10]);
  buf(\xm8051_golden_model_1.n0983 [107], input_sha_func_11[11]);
  buf(\xm8051_golden_model_1.n0983 [108], input_sha_func_11[12]);
  buf(\xm8051_golden_model_1.n0983 [109], input_sha_func_11[13]);
  buf(\xm8051_golden_model_1.n0983 [110], input_sha_func_11[14]);
  buf(\xm8051_golden_model_1.n0983 [111], input_sha_func_11[15]);
  buf(\xm8051_golden_model_1.n0983 [112], input_sha_func_11[16]);
  buf(\xm8051_golden_model_1.n0983 [113], input_sha_func_11[17]);
  buf(\xm8051_golden_model_1.n0983 [114], input_sha_func_11[18]);
  buf(\xm8051_golden_model_1.n0983 [115], input_sha_func_11[19]);
  buf(\xm8051_golden_model_1.n0983 [116], input_sha_func_11[20]);
  buf(\xm8051_golden_model_1.n0983 [117], input_sha_func_11[21]);
  buf(\xm8051_golden_model_1.n0983 [118], input_sha_func_11[22]);
  buf(\xm8051_golden_model_1.n0983 [119], input_sha_func_11[23]);
  buf(\xm8051_golden_model_1.n0983 [120], input_sha_func_11[24]);
  buf(\xm8051_golden_model_1.n0983 [121], input_sha_func_11[25]);
  buf(\xm8051_golden_model_1.n0983 [122], input_sha_func_11[26]);
  buf(\xm8051_golden_model_1.n0983 [123], input_sha_func_11[27]);
  buf(\xm8051_golden_model_1.n0983 [124], input_sha_func_11[28]);
  buf(\xm8051_golden_model_1.n0983 [125], input_sha_func_11[29]);
  buf(\xm8051_golden_model_1.n0983 [126], input_sha_func_11[30]);
  buf(\xm8051_golden_model_1.n0983 [127], input_sha_func_11[31]);
  buf(\xm8051_golden_model_1.n0983 [128], input_sha_func_11[32]);
  buf(\xm8051_golden_model_1.n0983 [129], input_sha_func_11[33]);
  buf(\xm8051_golden_model_1.n0983 [130], input_sha_func_11[34]);
  buf(\xm8051_golden_model_1.n0983 [131], input_sha_func_11[35]);
  buf(\xm8051_golden_model_1.n0983 [132], input_sha_func_11[36]);
  buf(\xm8051_golden_model_1.n0983 [133], input_sha_func_11[37]);
  buf(\xm8051_golden_model_1.n0983 [134], input_sha_func_11[38]);
  buf(\xm8051_golden_model_1.n0983 [135], input_sha_func_11[39]);
  buf(\xm8051_golden_model_1.n0983 [136], input_sha_func_11[40]);
  buf(\xm8051_golden_model_1.n0983 [137], input_sha_func_11[41]);
  buf(\xm8051_golden_model_1.n0983 [138], input_sha_func_11[42]);
  buf(\xm8051_golden_model_1.n0983 [139], input_sha_func_11[43]);
  buf(\xm8051_golden_model_1.n0983 [140], input_sha_func_11[44]);
  buf(\xm8051_golden_model_1.n0983 [141], input_sha_func_11[45]);
  buf(\xm8051_golden_model_1.n0983 [142], input_sha_func_11[46]);
  buf(\xm8051_golden_model_1.n0983 [143], input_sha_func_11[47]);
  buf(\xm8051_golden_model_1.n0983 [144], input_sha_func_11[48]);
  buf(\xm8051_golden_model_1.n0983 [145], input_sha_func_11[49]);
  buf(\xm8051_golden_model_1.n0983 [146], input_sha_func_11[50]);
  buf(\xm8051_golden_model_1.n0983 [147], input_sha_func_11[51]);
  buf(\xm8051_golden_model_1.n0983 [148], input_sha_func_11[52]);
  buf(\xm8051_golden_model_1.n0983 [149], input_sha_func_11[53]);
  buf(\xm8051_golden_model_1.n0983 [150], input_sha_func_11[54]);
  buf(\xm8051_golden_model_1.n0983 [151], input_sha_func_11[55]);
  buf(\xm8051_golden_model_1.n0983 [152], input_sha_func_11[56]);
  buf(\xm8051_golden_model_1.n0983 [153], input_sha_func_11[57]);
  buf(\xm8051_golden_model_1.n0983 [154], input_sha_func_11[58]);
  buf(\xm8051_golden_model_1.n0983 [155], input_sha_func_11[59]);
  buf(\xm8051_golden_model_1.n0983 [156], input_sha_func_11[60]);
  buf(\xm8051_golden_model_1.n0983 [157], input_sha_func_11[61]);
  buf(\xm8051_golden_model_1.n0983 [158], input_sha_func_11[62]);
  buf(\xm8051_golden_model_1.n0983 [159], input_sha_func_11[63]);
  buf(\xm8051_golden_model_1.n0099 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0099 [1], \xm8051_golden_model_1.n0187 [1]);
  buf(\xm8051_golden_model_1.n0099 [2], \xm8051_golden_model_1.n0187 [2]);
  buf(\xm8051_golden_model_1.n0973 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0973 [1], \xm8051_golden_model_1.aes_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0973 [2], \xm8051_golden_model_1.aes_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n0973 [3], \xm8051_golden_model_1.aes_bytes_processed [3]);
  buf(\xm8051_golden_model_1.n0086 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0086 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0086 [2], \xm8051_golden_model_1.n0473 [2]);
  buf(\xm8051_golden_model_1.n0086 [3], \xm8051_golden_model_1.n0433 [3]);
  buf(\xm8051_golden_model_1.n0086 [4], \xm8051_golden_model_1.n0341 [4]);
  buf(\xm8051_golden_model_1.n0972 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0972 [1], \xm8051_golden_model_1.aes_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0972 [2], \xm8051_golden_model_1.aes_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n0972 [3], \xm8051_golden_model_1.aes_bytes_processed [3]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [0], ABINPUT000[1]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [1], ABINPUT000[2]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [2], ABINPUT000[3]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [3], ABINPUT000[4]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [4], ABINPUT000[5]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [5], ABINPUT000[6]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [6], ABINPUT000[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [7], ABINPUT000[8]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [8], ABINPUT000[9]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [9], ABINPUT000[10]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [10], ABINPUT000[11]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [11], ABINPUT000[12]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [12], ABINPUT000[13]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [13], ABINPUT000[14]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [14], ABINPUT000[15]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [15], ABINPUT000[16]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [16], ABINPUT000[17]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [17], ABINPUT000[18]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [18], ABINPUT000[19]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [19], ABINPUT000[20]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [20], ABINPUT000[21]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [21], ABINPUT000[22]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [22], ABINPUT000[23]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [23], ABINPUT000[24]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [24], ABINPUT000[25]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [25], ABINPUT000[26]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [26], ABINPUT000[27]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [27], ABINPUT000[28]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [28], ABINPUT000[29]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [29], ABINPUT000[30]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [30], ABINPUT000[31]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [31], ABINPUT000[32]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [32], ABINPUT000[33]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [33], ABINPUT000[34]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [34], ABINPUT000[35]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [35], ABINPUT000[36]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [36], ABINPUT000[37]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [37], ABINPUT000[38]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [38], ABINPUT000[39]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [39], ABINPUT000[40]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [40], ABINPUT000[41]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [41], ABINPUT000[42]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [42], ABINPUT000[43]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [43], ABINPUT000[44]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [44], ABINPUT000[45]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [45], ABINPUT000[46]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [46], ABINPUT000[47]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [47], ABINPUT000[48]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [48], ABINPUT000[49]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [49], ABINPUT000[50]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [50], ABINPUT000[51]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [51], ABINPUT000[52]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [52], ABINPUT000[53]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [53], ABINPUT000[54]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [54], ABINPUT000[55]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [55], ABINPUT000[56]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [56], ABINPUT000[57]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [57], ABINPUT000[58]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [58], ABINPUT000[59]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [59], ABINPUT000[60]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [60], ABINPUT000[61]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [61], ABINPUT000[62]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [62], ABINPUT000[63]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [63], ABINPUT000[64]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [64], ABINPUT000[65]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [65], ABINPUT000[66]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [66], ABINPUT000[67]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [67], ABINPUT000[68]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [68], ABINPUT000[69]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [69], ABINPUT000[70]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [70], ABINPUT000[71]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [71], ABINPUT000[72]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [72], ABINPUT000[73]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [73], ABINPUT000[74]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [74], ABINPUT000[75]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [75], ABINPUT000[76]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [76], ABINPUT000[77]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [77], ABINPUT000[78]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [78], ABINPUT000[79]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [79], ABINPUT000[80]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [80], ABINPUT000[81]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [81], ABINPUT000[82]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [82], ABINPUT000[83]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [83], ABINPUT000[84]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [84], ABINPUT000[85]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [85], ABINPUT000[86]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [86], ABINPUT000[87]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [87], ABINPUT000[88]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [88], ABINPUT000[89]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [89], ABINPUT000[90]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [90], ABINPUT000[91]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [91], ABINPUT000[92]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [92], ABINPUT000[93]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [93], ABINPUT000[94]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [94], ABINPUT000[95]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [95], ABINPUT000[96]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [96], ABINPUT000[97]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [97], ABINPUT000[98]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [98], ABINPUT000[99]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [99], ABINPUT000[100]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [100], ABINPUT000[101]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [101], ABINPUT000[102]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [102], ABINPUT000[103]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [103], ABINPUT000[104]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [104], ABINPUT000[105]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [105], ABINPUT000[106]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [106], ABINPUT000[107]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [107], ABINPUT000[108]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [108], ABINPUT000[109]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [109], ABINPUT000[110]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [110], ABINPUT000[111]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [111], ABINPUT000[112]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [112], ABINPUT000[113]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [113], ABINPUT000[114]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [114], ABINPUT000[115]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [115], ABINPUT000[116]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [116], ABINPUT000[117]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [117], ABINPUT000[118]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [118], ABINPUT000[119]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [119], ABINPUT000[120]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [120], ABINPUT000[121]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [121], ABINPUT000[122]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [122], ABINPUT000[123]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [123], ABINPUT000[124]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [124], ABINPUT000[125]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [125], ABINPUT000[126]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [126], ABINPUT000[127]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [127], ABINPUT000[128]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [128], ABINPUT000[129]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [129], ABINPUT000[130]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [130], ABINPUT000[131]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [131], ABINPUT000[132]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [132], ABINPUT000[133]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [133], ABINPUT000[134]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [134], ABINPUT000[135]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [135], ABINPUT000[136]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [136], ABINPUT000[137]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [137], ABINPUT000[138]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [138], ABINPUT000[139]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [139], ABINPUT000[140]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [140], ABINPUT000[141]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [141], ABINPUT000[142]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [142], ABINPUT000[143]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [143], ABINPUT000[144]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [144], ABINPUT000[145]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [145], ABINPUT000[146]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [146], ABINPUT000[147]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [147], ABINPUT000[148]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [148], ABINPUT000[149]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [149], ABINPUT000[150]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [150], ABINPUT000[151]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [151], ABINPUT000[152]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [152], ABINPUT000[153]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [153], ABINPUT000[154]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [154], ABINPUT000[155]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [155], ABINPUT000[156]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [156], ABINPUT000[157]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [157], ABINPUT000[158]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [158], ABINPUT000[159]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest [159], ABINPUT000[160]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_digest_valid , ABINPUT000[161]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_core_ready , ABINPUT000[0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [0], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [1], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [1]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [2], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [2]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [3], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [3]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [4], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [4]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [5], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [5]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [6], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [6]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [7], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [8], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [8]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [9], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [9]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [10], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [10]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [11], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [11]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [12], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [12]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [13], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [13]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [14], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [14]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_reg_len [15], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [15]);
  buf(\xm8051_golden_model_1.n0968 [0], input_sha_func_10[0]);
  buf(\xm8051_golden_model_1.n0968 [1], input_sha_func_10[1]);
  buf(\xm8051_golden_model_1.n0968 [2], input_sha_func_10[2]);
  buf(\xm8051_golden_model_1.n0968 [3], input_sha_func_10[3]);
  buf(\xm8051_golden_model_1.n0968 [4], input_sha_func_10[4]);
  buf(\xm8051_golden_model_1.n0968 [5], input_sha_func_10[5]);
  buf(\xm8051_golden_model_1.n0968 [6], input_sha_func_10[6]);
  buf(\xm8051_golden_model_1.n0968 [7], input_sha_func_10[7]);
  buf(\xm8051_golden_model_1.n0968 [8], input_sha_func_10[8]);
  buf(\xm8051_golden_model_1.n0968 [9], input_sha_func_10[9]);
  buf(\xm8051_golden_model_1.n0968 [10], input_sha_func_10[10]);
  buf(\xm8051_golden_model_1.n0968 [11], input_sha_func_10[11]);
  buf(\xm8051_golden_model_1.n0968 [12], input_sha_func_10[12]);
  buf(\xm8051_golden_model_1.n0968 [13], input_sha_func_10[13]);
  buf(\xm8051_golden_model_1.n0968 [14], input_sha_func_10[14]);
  buf(\xm8051_golden_model_1.n0968 [15], input_sha_func_10[15]);
  buf(\xm8051_golden_model_1.n0968 [16], input_sha_func_10[16]);
  buf(\xm8051_golden_model_1.n0968 [17], input_sha_func_10[17]);
  buf(\xm8051_golden_model_1.n0968 [18], input_sha_func_10[18]);
  buf(\xm8051_golden_model_1.n0968 [19], input_sha_func_10[19]);
  buf(\xm8051_golden_model_1.n0968 [20], input_sha_func_10[20]);
  buf(\xm8051_golden_model_1.n0968 [21], input_sha_func_10[21]);
  buf(\xm8051_golden_model_1.n0968 [22], input_sha_func_10[22]);
  buf(\xm8051_golden_model_1.n0968 [23], input_sha_func_10[23]);
  buf(\xm8051_golden_model_1.n0968 [24], input_sha_func_10[24]);
  buf(\xm8051_golden_model_1.n0968 [25], input_sha_func_10[25]);
  buf(\xm8051_golden_model_1.n0968 [26], input_sha_func_10[26]);
  buf(\xm8051_golden_model_1.n0968 [27], input_sha_func_10[27]);
  buf(\xm8051_golden_model_1.n0968 [28], input_sha_func_10[28]);
  buf(\xm8051_golden_model_1.n0968 [29], input_sha_func_10[29]);
  buf(\xm8051_golden_model_1.n0968 [30], input_sha_func_10[30]);
  buf(\xm8051_golden_model_1.n0968 [31], input_sha_func_10[31]);
  buf(\xm8051_golden_model_1.n0968 [32], input_sha_func_9[0]);
  buf(\xm8051_golden_model_1.n0968 [33], input_sha_func_9[1]);
  buf(\xm8051_golden_model_1.n0968 [34], input_sha_func_9[2]);
  buf(\xm8051_golden_model_1.n0968 [35], input_sha_func_9[3]);
  buf(\xm8051_golden_model_1.n0968 [36], input_sha_func_9[4]);
  buf(\xm8051_golden_model_1.n0968 [37], input_sha_func_9[5]);
  buf(\xm8051_golden_model_1.n0968 [38], input_sha_func_9[6]);
  buf(\xm8051_golden_model_1.n0968 [39], input_sha_func_9[7]);
  buf(\xm8051_golden_model_1.n0968 [40], input_sha_func_9[8]);
  buf(\xm8051_golden_model_1.n0968 [41], input_sha_func_9[9]);
  buf(\xm8051_golden_model_1.n0968 [42], input_sha_func_9[10]);
  buf(\xm8051_golden_model_1.n0968 [43], input_sha_func_9[11]);
  buf(\xm8051_golden_model_1.n0968 [44], input_sha_func_9[12]);
  buf(\xm8051_golden_model_1.n0968 [45], input_sha_func_9[13]);
  buf(\xm8051_golden_model_1.n0968 [46], input_sha_func_9[14]);
  buf(\xm8051_golden_model_1.n0968 [47], input_sha_func_9[15]);
  buf(\xm8051_golden_model_1.n0968 [48], input_sha_func_9[16]);
  buf(\xm8051_golden_model_1.n0968 [49], input_sha_func_9[17]);
  buf(\xm8051_golden_model_1.n0968 [50], input_sha_func_9[18]);
  buf(\xm8051_golden_model_1.n0968 [51], input_sha_func_9[19]);
  buf(\xm8051_golden_model_1.n0968 [52], input_sha_func_9[20]);
  buf(\xm8051_golden_model_1.n0968 [53], input_sha_func_9[21]);
  buf(\xm8051_golden_model_1.n0968 [54], input_sha_func_9[22]);
  buf(\xm8051_golden_model_1.n0968 [55], input_sha_func_9[23]);
  buf(\xm8051_golden_model_1.n0968 [56], input_sha_func_9[24]);
  buf(\xm8051_golden_model_1.n0968 [57], input_sha_func_9[25]);
  buf(\xm8051_golden_model_1.n0968 [58], input_sha_func_9[26]);
  buf(\xm8051_golden_model_1.n0968 [59], input_sha_func_9[27]);
  buf(\xm8051_golden_model_1.n0968 [60], input_sha_func_9[28]);
  buf(\xm8051_golden_model_1.n0968 [61], input_sha_func_9[29]);
  buf(\xm8051_golden_model_1.n0968 [62], input_sha_func_9[30]);
  buf(\xm8051_golden_model_1.n0968 [63], input_sha_func_9[31]);
  buf(\xm8051_golden_model_1.n0968 [64], input_sha_func_9[32]);
  buf(\xm8051_golden_model_1.n0968 [65], input_sha_func_9[33]);
  buf(\xm8051_golden_model_1.n0968 [66], input_sha_func_9[34]);
  buf(\xm8051_golden_model_1.n0968 [67], input_sha_func_9[35]);
  buf(\xm8051_golden_model_1.n0968 [68], input_sha_func_9[36]);
  buf(\xm8051_golden_model_1.n0968 [69], input_sha_func_9[37]);
  buf(\xm8051_golden_model_1.n0968 [70], input_sha_func_9[38]);
  buf(\xm8051_golden_model_1.n0968 [71], input_sha_func_9[39]);
  buf(\xm8051_golden_model_1.n0968 [72], input_sha_func_9[40]);
  buf(\xm8051_golden_model_1.n0968 [73], input_sha_func_9[41]);
  buf(\xm8051_golden_model_1.n0968 [74], input_sha_func_9[42]);
  buf(\xm8051_golden_model_1.n0968 [75], input_sha_func_9[43]);
  buf(\xm8051_golden_model_1.n0968 [76], input_sha_func_9[44]);
  buf(\xm8051_golden_model_1.n0968 [77], input_sha_func_9[45]);
  buf(\xm8051_golden_model_1.n0968 [78], input_sha_func_9[46]);
  buf(\xm8051_golden_model_1.n0968 [79], input_sha_func_9[47]);
  buf(\xm8051_golden_model_1.n0968 [80], input_sha_func_9[48]);
  buf(\xm8051_golden_model_1.n0968 [81], input_sha_func_9[49]);
  buf(\xm8051_golden_model_1.n0968 [82], input_sha_func_9[50]);
  buf(\xm8051_golden_model_1.n0968 [83], input_sha_func_9[51]);
  buf(\xm8051_golden_model_1.n0968 [84], input_sha_func_9[52]);
  buf(\xm8051_golden_model_1.n0968 [85], input_sha_func_9[53]);
  buf(\xm8051_golden_model_1.n0968 [86], input_sha_func_9[54]);
  buf(\xm8051_golden_model_1.n0968 [87], input_sha_func_9[55]);
  buf(\xm8051_golden_model_1.n0968 [88], input_sha_func_9[56]);
  buf(\xm8051_golden_model_1.n0968 [89], input_sha_func_9[57]);
  buf(\xm8051_golden_model_1.n0968 [90], input_sha_func_9[58]);
  buf(\xm8051_golden_model_1.n0968 [91], input_sha_func_9[59]);
  buf(\xm8051_golden_model_1.n0968 [92], input_sha_func_9[60]);
  buf(\xm8051_golden_model_1.n0968 [93], input_sha_func_9[61]);
  buf(\xm8051_golden_model_1.n0968 [94], input_sha_func_9[62]);
  buf(\xm8051_golden_model_1.n0968 [95], input_sha_func_9[63]);
  buf(\xm8051_golden_model_1.n0968 [96], input_sha_func_8[0]);
  buf(\xm8051_golden_model_1.n0968 [97], input_sha_func_8[1]);
  buf(\xm8051_golden_model_1.n0968 [98], input_sha_func_8[2]);
  buf(\xm8051_golden_model_1.n0968 [99], input_sha_func_8[3]);
  buf(\xm8051_golden_model_1.n0968 [100], input_sha_func_8[4]);
  buf(\xm8051_golden_model_1.n0968 [101], input_sha_func_8[5]);
  buf(\xm8051_golden_model_1.n0968 [102], input_sha_func_8[6]);
  buf(\xm8051_golden_model_1.n0968 [103], input_sha_func_8[7]);
  buf(\xm8051_golden_model_1.n0968 [104], input_sha_func_8[8]);
  buf(\xm8051_golden_model_1.n0968 [105], input_sha_func_8[9]);
  buf(\xm8051_golden_model_1.n0968 [106], input_sha_func_8[10]);
  buf(\xm8051_golden_model_1.n0968 [107], input_sha_func_8[11]);
  buf(\xm8051_golden_model_1.n0968 [108], input_sha_func_8[12]);
  buf(\xm8051_golden_model_1.n0968 [109], input_sha_func_8[13]);
  buf(\xm8051_golden_model_1.n0968 [110], input_sha_func_8[14]);
  buf(\xm8051_golden_model_1.n0968 [111], input_sha_func_8[15]);
  buf(\xm8051_golden_model_1.n0968 [112], input_sha_func_8[16]);
  buf(\xm8051_golden_model_1.n0968 [113], input_sha_func_8[17]);
  buf(\xm8051_golden_model_1.n0968 [114], input_sha_func_8[18]);
  buf(\xm8051_golden_model_1.n0968 [115], input_sha_func_8[19]);
  buf(\xm8051_golden_model_1.n0968 [116], input_sha_func_8[20]);
  buf(\xm8051_golden_model_1.n0968 [117], input_sha_func_8[21]);
  buf(\xm8051_golden_model_1.n0968 [118], input_sha_func_8[22]);
  buf(\xm8051_golden_model_1.n0968 [119], input_sha_func_8[23]);
  buf(\xm8051_golden_model_1.n0968 [120], input_sha_func_8[24]);
  buf(\xm8051_golden_model_1.n0968 [121], input_sha_func_8[25]);
  buf(\xm8051_golden_model_1.n0968 [122], input_sha_func_8[26]);
  buf(\xm8051_golden_model_1.n0968 [123], input_sha_func_8[27]);
  buf(\xm8051_golden_model_1.n0968 [124], input_sha_func_8[28]);
  buf(\xm8051_golden_model_1.n0968 [125], input_sha_func_8[29]);
  buf(\xm8051_golden_model_1.n0968 [126], input_sha_func_8[30]);
  buf(\xm8051_golden_model_1.n0968 [127], input_sha_func_8[31]);
  buf(\xm8051_golden_model_1.n0968 [128], input_sha_func_8[32]);
  buf(\xm8051_golden_model_1.n0968 [129], input_sha_func_8[33]);
  buf(\xm8051_golden_model_1.n0968 [130], input_sha_func_8[34]);
  buf(\xm8051_golden_model_1.n0968 [131], input_sha_func_8[35]);
  buf(\xm8051_golden_model_1.n0968 [132], input_sha_func_8[36]);
  buf(\xm8051_golden_model_1.n0968 [133], input_sha_func_8[37]);
  buf(\xm8051_golden_model_1.n0968 [134], input_sha_func_8[38]);
  buf(\xm8051_golden_model_1.n0968 [135], input_sha_func_8[39]);
  buf(\xm8051_golden_model_1.n0968 [136], input_sha_func_8[40]);
  buf(\xm8051_golden_model_1.n0968 [137], input_sha_func_8[41]);
  buf(\xm8051_golden_model_1.n0968 [138], input_sha_func_8[42]);
  buf(\xm8051_golden_model_1.n0968 [139], input_sha_func_8[43]);
  buf(\xm8051_golden_model_1.n0968 [140], input_sha_func_8[44]);
  buf(\xm8051_golden_model_1.n0968 [141], input_sha_func_8[45]);
  buf(\xm8051_golden_model_1.n0968 [142], input_sha_func_8[46]);
  buf(\xm8051_golden_model_1.n0968 [143], input_sha_func_8[47]);
  buf(\xm8051_golden_model_1.n0968 [144], input_sha_func_8[48]);
  buf(\xm8051_golden_model_1.n0968 [145], input_sha_func_8[49]);
  buf(\xm8051_golden_model_1.n0968 [146], input_sha_func_8[50]);
  buf(\xm8051_golden_model_1.n0968 [147], input_sha_func_8[51]);
  buf(\xm8051_golden_model_1.n0968 [148], input_sha_func_8[52]);
  buf(\xm8051_golden_model_1.n0968 [149], input_sha_func_8[53]);
  buf(\xm8051_golden_model_1.n0968 [150], input_sha_func_8[54]);
  buf(\xm8051_golden_model_1.n0968 [151], input_sha_func_8[55]);
  buf(\xm8051_golden_model_1.n0968 [152], input_sha_func_8[56]);
  buf(\xm8051_golden_model_1.n0968 [153], input_sha_func_8[57]);
  buf(\xm8051_golden_model_1.n0968 [154], input_sha_func_8[58]);
  buf(\xm8051_golden_model_1.n0968 [155], input_sha_func_8[59]);
  buf(\xm8051_golden_model_1.n0968 [156], input_sha_func_8[60]);
  buf(\xm8051_golden_model_1.n0968 [157], input_sha_func_8[61]);
  buf(\xm8051_golden_model_1.n0968 [158], input_sha_func_8[62]);
  buf(\xm8051_golden_model_1.n0968 [159], input_sha_func_8[63]);
  buf(\xm8051_golden_model_1.n0966 [0], input_aes_func_7[0]);
  buf(\xm8051_golden_model_1.n0966 [1], input_aes_func_7[1]);
  buf(\xm8051_golden_model_1.n0966 [2], input_aes_func_7[2]);
  buf(\xm8051_golden_model_1.n0966 [3], input_aes_func_7[3]);
  buf(\xm8051_golden_model_1.n0966 [4], input_aes_func_7[4]);
  buf(\xm8051_golden_model_1.n0966 [5], input_aes_func_7[5]);
  buf(\xm8051_golden_model_1.n0966 [6], input_aes_func_7[6]);
  buf(\xm8051_golden_model_1.n0966 [7], input_aes_func_7[7]);
  buf(\xm8051_golden_model_1.n0966 [8], input_aes_func_7[8]);
  buf(\xm8051_golden_model_1.n0966 [9], input_aes_func_7[9]);
  buf(\xm8051_golden_model_1.n0966 [10], input_aes_func_7[10]);
  buf(\xm8051_golden_model_1.n0966 [11], input_aes_func_7[11]);
  buf(\xm8051_golden_model_1.n0966 [12], input_aes_func_7[12]);
  buf(\xm8051_golden_model_1.n0966 [13], input_aes_func_7[13]);
  buf(\xm8051_golden_model_1.n0966 [14], input_aes_func_7[14]);
  buf(\xm8051_golden_model_1.n0966 [15], input_aes_func_7[15]);
  buf(\xm8051_golden_model_1.n0966 [16], input_aes_func_7[16]);
  buf(\xm8051_golden_model_1.n0966 [17], input_aes_func_7[17]);
  buf(\xm8051_golden_model_1.n0966 [18], input_aes_func_7[18]);
  buf(\xm8051_golden_model_1.n0966 [19], input_aes_func_7[19]);
  buf(\xm8051_golden_model_1.n0966 [20], input_aes_func_7[20]);
  buf(\xm8051_golden_model_1.n0966 [21], input_aes_func_7[21]);
  buf(\xm8051_golden_model_1.n0966 [22], input_aes_func_7[22]);
  buf(\xm8051_golden_model_1.n0966 [23], input_aes_func_7[23]);
  buf(\xm8051_golden_model_1.n0966 [24], input_aes_func_7[24]);
  buf(\xm8051_golden_model_1.n0966 [25], input_aes_func_7[25]);
  buf(\xm8051_golden_model_1.n0966 [26], input_aes_func_7[26]);
  buf(\xm8051_golden_model_1.n0966 [27], input_aes_func_7[27]);
  buf(\xm8051_golden_model_1.n0966 [28], input_aes_func_7[28]);
  buf(\xm8051_golden_model_1.n0966 [29], input_aes_func_7[29]);
  buf(\xm8051_golden_model_1.n0966 [30], input_aes_func_7[30]);
  buf(\xm8051_golden_model_1.n0966 [31], input_aes_func_7[31]);
  buf(\xm8051_golden_model_1.n0966 [32], input_aes_func_7[32]);
  buf(\xm8051_golden_model_1.n0966 [33], input_aes_func_7[33]);
  buf(\xm8051_golden_model_1.n0966 [34], input_aes_func_7[34]);
  buf(\xm8051_golden_model_1.n0966 [35], input_aes_func_7[35]);
  buf(\xm8051_golden_model_1.n0966 [36], input_aes_func_7[36]);
  buf(\xm8051_golden_model_1.n0966 [37], input_aes_func_7[37]);
  buf(\xm8051_golden_model_1.n0966 [38], input_aes_func_7[38]);
  buf(\xm8051_golden_model_1.n0966 [39], input_aes_func_7[39]);
  buf(\xm8051_golden_model_1.n0966 [40], input_aes_func_7[40]);
  buf(\xm8051_golden_model_1.n0966 [41], input_aes_func_7[41]);
  buf(\xm8051_golden_model_1.n0966 [42], input_aes_func_7[42]);
  buf(\xm8051_golden_model_1.n0966 [43], input_aes_func_7[43]);
  buf(\xm8051_golden_model_1.n0966 [44], input_aes_func_7[44]);
  buf(\xm8051_golden_model_1.n0966 [45], input_aes_func_7[45]);
  buf(\xm8051_golden_model_1.n0966 [46], input_aes_func_7[46]);
  buf(\xm8051_golden_model_1.n0966 [47], input_aes_func_7[47]);
  buf(\xm8051_golden_model_1.n0966 [48], input_aes_func_7[48]);
  buf(\xm8051_golden_model_1.n0966 [49], input_aes_func_7[49]);
  buf(\xm8051_golden_model_1.n0966 [50], input_aes_func_7[50]);
  buf(\xm8051_golden_model_1.n0966 [51], input_aes_func_7[51]);
  buf(\xm8051_golden_model_1.n0966 [52], input_aes_func_7[52]);
  buf(\xm8051_golden_model_1.n0966 [53], input_aes_func_7[53]);
  buf(\xm8051_golden_model_1.n0966 [54], input_aes_func_7[54]);
  buf(\xm8051_golden_model_1.n0966 [55], input_aes_func_7[55]);
  buf(\xm8051_golden_model_1.n0966 [56], input_aes_func_7[56]);
  buf(\xm8051_golden_model_1.n0966 [57], input_aes_func_7[57]);
  buf(\xm8051_golden_model_1.n0966 [58], input_aes_func_7[58]);
  buf(\xm8051_golden_model_1.n0966 [59], input_aes_func_7[59]);
  buf(\xm8051_golden_model_1.n0966 [60], input_aes_func_7[60]);
  buf(\xm8051_golden_model_1.n0966 [61], input_aes_func_7[61]);
  buf(\xm8051_golden_model_1.n0966 [62], input_aes_func_7[62]);
  buf(\xm8051_golden_model_1.n0966 [63], input_aes_func_7[63]);
  buf(\xm8051_golden_model_1.n0966 [64], input_aes_func_6[0]);
  buf(\xm8051_golden_model_1.n0966 [65], input_aes_func_6[1]);
  buf(\xm8051_golden_model_1.n0966 [66], input_aes_func_6[2]);
  buf(\xm8051_golden_model_1.n0966 [67], input_aes_func_6[3]);
  buf(\xm8051_golden_model_1.n0966 [68], input_aes_func_6[4]);
  buf(\xm8051_golden_model_1.n0966 [69], input_aes_func_6[5]);
  buf(\xm8051_golden_model_1.n0966 [70], input_aes_func_6[6]);
  buf(\xm8051_golden_model_1.n0966 [71], input_aes_func_6[7]);
  buf(\xm8051_golden_model_1.n0966 [72], input_aes_func_6[8]);
  buf(\xm8051_golden_model_1.n0966 [73], input_aes_func_6[9]);
  buf(\xm8051_golden_model_1.n0966 [74], input_aes_func_6[10]);
  buf(\xm8051_golden_model_1.n0966 [75], input_aes_func_6[11]);
  buf(\xm8051_golden_model_1.n0966 [76], input_aes_func_6[12]);
  buf(\xm8051_golden_model_1.n0966 [77], input_aes_func_6[13]);
  buf(\xm8051_golden_model_1.n0966 [78], input_aes_func_6[14]);
  buf(\xm8051_golden_model_1.n0966 [79], input_aes_func_6[15]);
  buf(\xm8051_golden_model_1.n0966 [80], input_aes_func_6[16]);
  buf(\xm8051_golden_model_1.n0966 [81], input_aes_func_6[17]);
  buf(\xm8051_golden_model_1.n0966 [82], input_aes_func_6[18]);
  buf(\xm8051_golden_model_1.n0966 [83], input_aes_func_6[19]);
  buf(\xm8051_golden_model_1.n0966 [84], input_aes_func_6[20]);
  buf(\xm8051_golden_model_1.n0966 [85], input_aes_func_6[21]);
  buf(\xm8051_golden_model_1.n0966 [86], input_aes_func_6[22]);
  buf(\xm8051_golden_model_1.n0966 [87], input_aes_func_6[23]);
  buf(\xm8051_golden_model_1.n0966 [88], input_aes_func_6[24]);
  buf(\xm8051_golden_model_1.n0966 [89], input_aes_func_6[25]);
  buf(\xm8051_golden_model_1.n0966 [90], input_aes_func_6[26]);
  buf(\xm8051_golden_model_1.n0966 [91], input_aes_func_6[27]);
  buf(\xm8051_golden_model_1.n0966 [92], input_aes_func_6[28]);
  buf(\xm8051_golden_model_1.n0966 [93], input_aes_func_6[29]);
  buf(\xm8051_golden_model_1.n0966 [94], input_aes_func_6[30]);
  buf(\xm8051_golden_model_1.n0966 [95], input_aes_func_6[31]);
  buf(\xm8051_golden_model_1.n0966 [96], input_aes_func_6[32]);
  buf(\xm8051_golden_model_1.n0966 [97], input_aes_func_6[33]);
  buf(\xm8051_golden_model_1.n0966 [98], input_aes_func_6[34]);
  buf(\xm8051_golden_model_1.n0966 [99], input_aes_func_6[35]);
  buf(\xm8051_golden_model_1.n0966 [100], input_aes_func_6[36]);
  buf(\xm8051_golden_model_1.n0966 [101], input_aes_func_6[37]);
  buf(\xm8051_golden_model_1.n0966 [102], input_aes_func_6[38]);
  buf(\xm8051_golden_model_1.n0966 [103], input_aes_func_6[39]);
  buf(\xm8051_golden_model_1.n0966 [104], input_aes_func_6[40]);
  buf(\xm8051_golden_model_1.n0966 [105], input_aes_func_6[41]);
  buf(\xm8051_golden_model_1.n0966 [106], input_aes_func_6[42]);
  buf(\xm8051_golden_model_1.n0966 [107], input_aes_func_6[43]);
  buf(\xm8051_golden_model_1.n0966 [108], input_aes_func_6[44]);
  buf(\xm8051_golden_model_1.n0966 [109], input_aes_func_6[45]);
  buf(\xm8051_golden_model_1.n0966 [110], input_aes_func_6[46]);
  buf(\xm8051_golden_model_1.n0966 [111], input_aes_func_6[47]);
  buf(\xm8051_golden_model_1.n0966 [112], input_aes_func_6[48]);
  buf(\xm8051_golden_model_1.n0966 [113], input_aes_func_6[49]);
  buf(\xm8051_golden_model_1.n0966 [114], input_aes_func_6[50]);
  buf(\xm8051_golden_model_1.n0966 [115], input_aes_func_6[51]);
  buf(\xm8051_golden_model_1.n0966 [116], input_aes_func_6[52]);
  buf(\xm8051_golden_model_1.n0966 [117], input_aes_func_6[53]);
  buf(\xm8051_golden_model_1.n0966 [118], input_aes_func_6[54]);
  buf(\xm8051_golden_model_1.n0966 [119], input_aes_func_6[55]);
  buf(\xm8051_golden_model_1.n0966 [120], input_aes_func_6[56]);
  buf(\xm8051_golden_model_1.n0966 [121], input_aes_func_6[57]);
  buf(\xm8051_golden_model_1.n0966 [122], input_aes_func_6[58]);
  buf(\xm8051_golden_model_1.n0966 [123], input_aes_func_6[59]);
  buf(\xm8051_golden_model_1.n0966 [124], input_aes_func_6[60]);
  buf(\xm8051_golden_model_1.n0966 [125], input_aes_func_6[61]);
  buf(\xm8051_golden_model_1.n0966 [126], input_aes_func_6[62]);
  buf(\xm8051_golden_model_1.n0966 [127], input_aes_func_6[63]);
  buf(\xm8051_golden_model_1.n0077 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0077 [1], \xm8051_golden_model_1.aes_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0077 [2], \xm8051_golden_model_1.n0165 [2]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_out_state [0], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_out_state [1], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [1]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_out_state [2], 1'b0);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_out_state [3], 1'b0);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_out_state [4], 1'b0);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_out_state [5], 1'b0);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_out_state [6], 1'b0);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_out_state [7], 1'b0);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.data_in [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.data_in [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.data_in [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.data_in [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.data_in [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.data_in [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.data_in [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.data_in [7], proc_data_in[7]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.addr [0], proc_addr[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.addr [1], proc_addr[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.addr [2], proc_addr[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.addr [3], proc_addr[3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.rst , rst);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key0_i.clk , clk);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [0], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [1], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [1]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [2], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [2]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [3], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [3]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [4], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [4]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [5], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [5]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [6], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [6]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [7], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [8], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [8]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [9], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [9]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [10], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [10]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [11], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [11]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [12], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [12]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [13], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [13]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [14], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [14]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_len [15], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [15]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_state [0], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.sha_state [1], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [1]);
  buf(\xm8051_golden_model_1.n0958 [0], input_sha_func_5[0]);
  buf(\xm8051_golden_model_1.n0958 [1], input_sha_func_5[1]);
  buf(\xm8051_golden_model_1.n0958 [2], input_sha_func_5[2]);
  buf(\xm8051_golden_model_1.n0958 [3], input_sha_func_5[3]);
  buf(\xm8051_golden_model_1.n0958 [4], input_sha_func_5[4]);
  buf(\xm8051_golden_model_1.n0958 [5], input_sha_func_5[5]);
  buf(\xm8051_golden_model_1.n0958 [6], input_sha_func_5[6]);
  buf(\xm8051_golden_model_1.n0958 [7], input_sha_func_5[7]);
  buf(\xm8051_golden_model_1.n0958 [8], input_sha_func_5[8]);
  buf(\xm8051_golden_model_1.n0958 [9], input_sha_func_5[9]);
  buf(\xm8051_golden_model_1.n0958 [10], input_sha_func_5[10]);
  buf(\xm8051_golden_model_1.n0958 [11], input_sha_func_5[11]);
  buf(\xm8051_golden_model_1.n0958 [12], input_sha_func_5[12]);
  buf(\xm8051_golden_model_1.n0958 [13], input_sha_func_5[13]);
  buf(\xm8051_golden_model_1.n0958 [14], input_sha_func_5[14]);
  buf(\xm8051_golden_model_1.n0958 [15], input_sha_func_5[15]);
  buf(\xm8051_golden_model_1.n0958 [16], input_sha_func_5[16]);
  buf(\xm8051_golden_model_1.n0958 [17], input_sha_func_5[17]);
  buf(\xm8051_golden_model_1.n0958 [18], input_sha_func_5[18]);
  buf(\xm8051_golden_model_1.n0958 [19], input_sha_func_5[19]);
  buf(\xm8051_golden_model_1.n0958 [20], input_sha_func_5[20]);
  buf(\xm8051_golden_model_1.n0958 [21], input_sha_func_5[21]);
  buf(\xm8051_golden_model_1.n0958 [22], input_sha_func_5[22]);
  buf(\xm8051_golden_model_1.n0958 [23], input_sha_func_5[23]);
  buf(\xm8051_golden_model_1.n0958 [24], input_sha_func_5[24]);
  buf(\xm8051_golden_model_1.n0958 [25], input_sha_func_5[25]);
  buf(\xm8051_golden_model_1.n0958 [26], input_sha_func_5[26]);
  buf(\xm8051_golden_model_1.n0958 [27], input_sha_func_5[27]);
  buf(\xm8051_golden_model_1.n0958 [28], input_sha_func_5[28]);
  buf(\xm8051_golden_model_1.n0958 [29], input_sha_func_5[29]);
  buf(\xm8051_golden_model_1.n0958 [30], input_sha_func_5[30]);
  buf(\xm8051_golden_model_1.n0958 [31], input_sha_func_5[31]);
  buf(\xm8051_golden_model_1.n0958 [32], input_sha_func_4[0]);
  buf(\xm8051_golden_model_1.n0958 [33], input_sha_func_4[1]);
  buf(\xm8051_golden_model_1.n0958 [34], input_sha_func_4[2]);
  buf(\xm8051_golden_model_1.n0958 [35], input_sha_func_4[3]);
  buf(\xm8051_golden_model_1.n0958 [36], input_sha_func_4[4]);
  buf(\xm8051_golden_model_1.n0958 [37], input_sha_func_4[5]);
  buf(\xm8051_golden_model_1.n0958 [38], input_sha_func_4[6]);
  buf(\xm8051_golden_model_1.n0958 [39], input_sha_func_4[7]);
  buf(\xm8051_golden_model_1.n0958 [40], input_sha_func_4[8]);
  buf(\xm8051_golden_model_1.n0958 [41], input_sha_func_4[9]);
  buf(\xm8051_golden_model_1.n0958 [42], input_sha_func_4[10]);
  buf(\xm8051_golden_model_1.n0958 [43], input_sha_func_4[11]);
  buf(\xm8051_golden_model_1.n0958 [44], input_sha_func_4[12]);
  buf(\xm8051_golden_model_1.n0958 [45], input_sha_func_4[13]);
  buf(\xm8051_golden_model_1.n0958 [46], input_sha_func_4[14]);
  buf(\xm8051_golden_model_1.n0958 [47], input_sha_func_4[15]);
  buf(\xm8051_golden_model_1.n0958 [48], input_sha_func_4[16]);
  buf(\xm8051_golden_model_1.n0958 [49], input_sha_func_4[17]);
  buf(\xm8051_golden_model_1.n0958 [50], input_sha_func_4[18]);
  buf(\xm8051_golden_model_1.n0958 [51], input_sha_func_4[19]);
  buf(\xm8051_golden_model_1.n0958 [52], input_sha_func_4[20]);
  buf(\xm8051_golden_model_1.n0958 [53], input_sha_func_4[21]);
  buf(\xm8051_golden_model_1.n0958 [54], input_sha_func_4[22]);
  buf(\xm8051_golden_model_1.n0958 [55], input_sha_func_4[23]);
  buf(\xm8051_golden_model_1.n0958 [56], input_sha_func_4[24]);
  buf(\xm8051_golden_model_1.n0958 [57], input_sha_func_4[25]);
  buf(\xm8051_golden_model_1.n0958 [58], input_sha_func_4[26]);
  buf(\xm8051_golden_model_1.n0958 [59], input_sha_func_4[27]);
  buf(\xm8051_golden_model_1.n0958 [60], input_sha_func_4[28]);
  buf(\xm8051_golden_model_1.n0958 [61], input_sha_func_4[29]);
  buf(\xm8051_golden_model_1.n0958 [62], input_sha_func_4[30]);
  buf(\xm8051_golden_model_1.n0958 [63], input_sha_func_4[31]);
  buf(\xm8051_golden_model_1.n0958 [64], input_sha_func_4[32]);
  buf(\xm8051_golden_model_1.n0958 [65], input_sha_func_4[33]);
  buf(\xm8051_golden_model_1.n0958 [66], input_sha_func_4[34]);
  buf(\xm8051_golden_model_1.n0958 [67], input_sha_func_4[35]);
  buf(\xm8051_golden_model_1.n0958 [68], input_sha_func_4[36]);
  buf(\xm8051_golden_model_1.n0958 [69], input_sha_func_4[37]);
  buf(\xm8051_golden_model_1.n0958 [70], input_sha_func_4[38]);
  buf(\xm8051_golden_model_1.n0958 [71], input_sha_func_4[39]);
  buf(\xm8051_golden_model_1.n0958 [72], input_sha_func_4[40]);
  buf(\xm8051_golden_model_1.n0958 [73], input_sha_func_4[41]);
  buf(\xm8051_golden_model_1.n0958 [74], input_sha_func_4[42]);
  buf(\xm8051_golden_model_1.n0958 [75], input_sha_func_4[43]);
  buf(\xm8051_golden_model_1.n0958 [76], input_sha_func_4[44]);
  buf(\xm8051_golden_model_1.n0958 [77], input_sha_func_4[45]);
  buf(\xm8051_golden_model_1.n0958 [78], input_sha_func_4[46]);
  buf(\xm8051_golden_model_1.n0958 [79], input_sha_func_4[47]);
  buf(\xm8051_golden_model_1.n0958 [80], input_sha_func_4[48]);
  buf(\xm8051_golden_model_1.n0958 [81], input_sha_func_4[49]);
  buf(\xm8051_golden_model_1.n0958 [82], input_sha_func_4[50]);
  buf(\xm8051_golden_model_1.n0958 [83], input_sha_func_4[51]);
  buf(\xm8051_golden_model_1.n0958 [84], input_sha_func_4[52]);
  buf(\xm8051_golden_model_1.n0958 [85], input_sha_func_4[53]);
  buf(\xm8051_golden_model_1.n0958 [86], input_sha_func_4[54]);
  buf(\xm8051_golden_model_1.n0958 [87], input_sha_func_4[55]);
  buf(\xm8051_golden_model_1.n0958 [88], input_sha_func_4[56]);
  buf(\xm8051_golden_model_1.n0958 [89], input_sha_func_4[57]);
  buf(\xm8051_golden_model_1.n0958 [90], input_sha_func_4[58]);
  buf(\xm8051_golden_model_1.n0958 [91], input_sha_func_4[59]);
  buf(\xm8051_golden_model_1.n0958 [92], input_sha_func_4[60]);
  buf(\xm8051_golden_model_1.n0958 [93], input_sha_func_4[61]);
  buf(\xm8051_golden_model_1.n0958 [94], input_sha_func_4[62]);
  buf(\xm8051_golden_model_1.n0958 [95], input_sha_func_4[63]);
  buf(\xm8051_golden_model_1.n0958 [96], input_sha_func_3[0]);
  buf(\xm8051_golden_model_1.n0958 [97], input_sha_func_3[1]);
  buf(\xm8051_golden_model_1.n0958 [98], input_sha_func_3[2]);
  buf(\xm8051_golden_model_1.n0958 [99], input_sha_func_3[3]);
  buf(\xm8051_golden_model_1.n0958 [100], input_sha_func_3[4]);
  buf(\xm8051_golden_model_1.n0958 [101], input_sha_func_3[5]);
  buf(\xm8051_golden_model_1.n0958 [102], input_sha_func_3[6]);
  buf(\xm8051_golden_model_1.n0958 [103], input_sha_func_3[7]);
  buf(\xm8051_golden_model_1.n0958 [104], input_sha_func_3[8]);
  buf(\xm8051_golden_model_1.n0958 [105], input_sha_func_3[9]);
  buf(\xm8051_golden_model_1.n0958 [106], input_sha_func_3[10]);
  buf(\xm8051_golden_model_1.n0958 [107], input_sha_func_3[11]);
  buf(\xm8051_golden_model_1.n0958 [108], input_sha_func_3[12]);
  buf(\xm8051_golden_model_1.n0958 [109], input_sha_func_3[13]);
  buf(\xm8051_golden_model_1.n0958 [110], input_sha_func_3[14]);
  buf(\xm8051_golden_model_1.n0958 [111], input_sha_func_3[15]);
  buf(\xm8051_golden_model_1.n0958 [112], input_sha_func_3[16]);
  buf(\xm8051_golden_model_1.n0958 [113], input_sha_func_3[17]);
  buf(\xm8051_golden_model_1.n0958 [114], input_sha_func_3[18]);
  buf(\xm8051_golden_model_1.n0958 [115], input_sha_func_3[19]);
  buf(\xm8051_golden_model_1.n0958 [116], input_sha_func_3[20]);
  buf(\xm8051_golden_model_1.n0958 [117], input_sha_func_3[21]);
  buf(\xm8051_golden_model_1.n0958 [118], input_sha_func_3[22]);
  buf(\xm8051_golden_model_1.n0958 [119], input_sha_func_3[23]);
  buf(\xm8051_golden_model_1.n0958 [120], input_sha_func_3[24]);
  buf(\xm8051_golden_model_1.n0958 [121], input_sha_func_3[25]);
  buf(\xm8051_golden_model_1.n0958 [122], input_sha_func_3[26]);
  buf(\xm8051_golden_model_1.n0958 [123], input_sha_func_3[27]);
  buf(\xm8051_golden_model_1.n0958 [124], input_sha_func_3[28]);
  buf(\xm8051_golden_model_1.n0958 [125], input_sha_func_3[29]);
  buf(\xm8051_golden_model_1.n0958 [126], input_sha_func_3[30]);
  buf(\xm8051_golden_model_1.n0958 [127], input_sha_func_3[31]);
  buf(\xm8051_golden_model_1.n0958 [128], input_sha_func_3[32]);
  buf(\xm8051_golden_model_1.n0958 [129], input_sha_func_3[33]);
  buf(\xm8051_golden_model_1.n0958 [130], input_sha_func_3[34]);
  buf(\xm8051_golden_model_1.n0958 [131], input_sha_func_3[35]);
  buf(\xm8051_golden_model_1.n0958 [132], input_sha_func_3[36]);
  buf(\xm8051_golden_model_1.n0958 [133], input_sha_func_3[37]);
  buf(\xm8051_golden_model_1.n0958 [134], input_sha_func_3[38]);
  buf(\xm8051_golden_model_1.n0958 [135], input_sha_func_3[39]);
  buf(\xm8051_golden_model_1.n0958 [136], input_sha_func_3[40]);
  buf(\xm8051_golden_model_1.n0958 [137], input_sha_func_3[41]);
  buf(\xm8051_golden_model_1.n0958 [138], input_sha_func_3[42]);
  buf(\xm8051_golden_model_1.n0958 [139], input_sha_func_3[43]);
  buf(\xm8051_golden_model_1.n0958 [140], input_sha_func_3[44]);
  buf(\xm8051_golden_model_1.n0958 [141], input_sha_func_3[45]);
  buf(\xm8051_golden_model_1.n0958 [142], input_sha_func_3[46]);
  buf(\xm8051_golden_model_1.n0958 [143], input_sha_func_3[47]);
  buf(\xm8051_golden_model_1.n0958 [144], input_sha_func_3[48]);
  buf(\xm8051_golden_model_1.n0958 [145], input_sha_func_3[49]);
  buf(\xm8051_golden_model_1.n0958 [146], input_sha_func_3[50]);
  buf(\xm8051_golden_model_1.n0958 [147], input_sha_func_3[51]);
  buf(\xm8051_golden_model_1.n0958 [148], input_sha_func_3[52]);
  buf(\xm8051_golden_model_1.n0958 [149], input_sha_func_3[53]);
  buf(\xm8051_golden_model_1.n0958 [150], input_sha_func_3[54]);
  buf(\xm8051_golden_model_1.n0958 [151], input_sha_func_3[55]);
  buf(\xm8051_golden_model_1.n0958 [152], input_sha_func_3[56]);
  buf(\xm8051_golden_model_1.n0958 [153], input_sha_func_3[57]);
  buf(\xm8051_golden_model_1.n0958 [154], input_sha_func_3[58]);
  buf(\xm8051_golden_model_1.n0958 [155], input_sha_func_3[59]);
  buf(\xm8051_golden_model_1.n0958 [156], input_sha_func_3[60]);
  buf(\xm8051_golden_model_1.n0958 [157], input_sha_func_3[61]);
  buf(\xm8051_golden_model_1.n0958 [158], input_sha_func_3[62]);
  buf(\xm8051_golden_model_1.n0958 [159], input_sha_func_3[63]);
  buf(\xm8051_golden_model_1.n0956 [0], RD_xram_16[0]);
  buf(\xm8051_golden_model_1.n0956 [1], RD_xram_16[1]);
  buf(\xm8051_golden_model_1.n0956 [2], RD_xram_16[2]);
  buf(\xm8051_golden_model_1.n0956 [3], RD_xram_16[3]);
  buf(\xm8051_golden_model_1.n0956 [4], RD_xram_16[4]);
  buf(\xm8051_golden_model_1.n0956 [5], RD_xram_16[5]);
  buf(\xm8051_golden_model_1.n0956 [6], RD_xram_16[6]);
  buf(\xm8051_golden_model_1.n0956 [7], RD_xram_16[7]);
  buf(\xm8051_golden_model_1.n0956 [8], RD_xram_15[0]);
  buf(\xm8051_golden_model_1.n0956 [9], RD_xram_15[1]);
  buf(\xm8051_golden_model_1.n0956 [10], RD_xram_15[2]);
  buf(\xm8051_golden_model_1.n0956 [11], RD_xram_15[3]);
  buf(\xm8051_golden_model_1.n0956 [12], RD_xram_15[4]);
  buf(\xm8051_golden_model_1.n0956 [13], RD_xram_15[5]);
  buf(\xm8051_golden_model_1.n0956 [14], RD_xram_15[6]);
  buf(\xm8051_golden_model_1.n0956 [15], RD_xram_15[7]);
  buf(\xm8051_golden_model_1.n0956 [16], RD_xram_14[0]);
  buf(\xm8051_golden_model_1.n0956 [17], RD_xram_14[1]);
  buf(\xm8051_golden_model_1.n0956 [18], RD_xram_14[2]);
  buf(\xm8051_golden_model_1.n0956 [19], RD_xram_14[3]);
  buf(\xm8051_golden_model_1.n0956 [20], RD_xram_14[4]);
  buf(\xm8051_golden_model_1.n0956 [21], RD_xram_14[5]);
  buf(\xm8051_golden_model_1.n0956 [22], RD_xram_14[6]);
  buf(\xm8051_golden_model_1.n0956 [23], RD_xram_14[7]);
  buf(\xm8051_golden_model_1.n0956 [24], RD_xram_13[0]);
  buf(\xm8051_golden_model_1.n0956 [25], RD_xram_13[1]);
  buf(\xm8051_golden_model_1.n0956 [26], RD_xram_13[2]);
  buf(\xm8051_golden_model_1.n0956 [27], RD_xram_13[3]);
  buf(\xm8051_golden_model_1.n0956 [28], RD_xram_13[4]);
  buf(\xm8051_golden_model_1.n0956 [29], RD_xram_13[5]);
  buf(\xm8051_golden_model_1.n0956 [30], RD_xram_13[6]);
  buf(\xm8051_golden_model_1.n0956 [31], RD_xram_13[7]);
  buf(\xm8051_golden_model_1.n0956 [32], RD_xram_12[0]);
  buf(\xm8051_golden_model_1.n0956 [33], RD_xram_12[1]);
  buf(\xm8051_golden_model_1.n0956 [34], RD_xram_12[2]);
  buf(\xm8051_golden_model_1.n0956 [35], RD_xram_12[3]);
  buf(\xm8051_golden_model_1.n0956 [36], RD_xram_12[4]);
  buf(\xm8051_golden_model_1.n0956 [37], RD_xram_12[5]);
  buf(\xm8051_golden_model_1.n0956 [38], RD_xram_12[6]);
  buf(\xm8051_golden_model_1.n0956 [39], RD_xram_12[7]);
  buf(\xm8051_golden_model_1.n0956 [40], RD_xram_11[0]);
  buf(\xm8051_golden_model_1.n0956 [41], RD_xram_11[1]);
  buf(\xm8051_golden_model_1.n0956 [42], RD_xram_11[2]);
  buf(\xm8051_golden_model_1.n0956 [43], RD_xram_11[3]);
  buf(\xm8051_golden_model_1.n0956 [44], RD_xram_11[4]);
  buf(\xm8051_golden_model_1.n0956 [45], RD_xram_11[5]);
  buf(\xm8051_golden_model_1.n0956 [46], RD_xram_11[6]);
  buf(\xm8051_golden_model_1.n0956 [47], RD_xram_11[7]);
  buf(\xm8051_golden_model_1.n0956 [48], RD_xram_10[0]);
  buf(\xm8051_golden_model_1.n0956 [49], RD_xram_10[1]);
  buf(\xm8051_golden_model_1.n0956 [50], RD_xram_10[2]);
  buf(\xm8051_golden_model_1.n0956 [51], RD_xram_10[3]);
  buf(\xm8051_golden_model_1.n0956 [52], RD_xram_10[4]);
  buf(\xm8051_golden_model_1.n0956 [53], RD_xram_10[5]);
  buf(\xm8051_golden_model_1.n0956 [54], RD_xram_10[6]);
  buf(\xm8051_golden_model_1.n0956 [55], RD_xram_10[7]);
  buf(\xm8051_golden_model_1.n0956 [56], RD_xram_9[0]);
  buf(\xm8051_golden_model_1.n0956 [57], RD_xram_9[1]);
  buf(\xm8051_golden_model_1.n0956 [58], RD_xram_9[2]);
  buf(\xm8051_golden_model_1.n0956 [59], RD_xram_9[3]);
  buf(\xm8051_golden_model_1.n0956 [60], RD_xram_9[4]);
  buf(\xm8051_golden_model_1.n0956 [61], RD_xram_9[5]);
  buf(\xm8051_golden_model_1.n0956 [62], RD_xram_9[6]);
  buf(\xm8051_golden_model_1.n0956 [63], RD_xram_9[7]);
  buf(\xm8051_golden_model_1.n0956 [64], RD_xram_8[0]);
  buf(\xm8051_golden_model_1.n0956 [65], RD_xram_8[1]);
  buf(\xm8051_golden_model_1.n0956 [66], RD_xram_8[2]);
  buf(\xm8051_golden_model_1.n0956 [67], RD_xram_8[3]);
  buf(\xm8051_golden_model_1.n0956 [68], RD_xram_8[4]);
  buf(\xm8051_golden_model_1.n0956 [69], RD_xram_8[5]);
  buf(\xm8051_golden_model_1.n0956 [70], RD_xram_8[6]);
  buf(\xm8051_golden_model_1.n0956 [71], RD_xram_8[7]);
  buf(\xm8051_golden_model_1.n0956 [72], RD_xram_7[0]);
  buf(\xm8051_golden_model_1.n0956 [73], RD_xram_7[1]);
  buf(\xm8051_golden_model_1.n0956 [74], RD_xram_7[2]);
  buf(\xm8051_golden_model_1.n0956 [75], RD_xram_7[3]);
  buf(\xm8051_golden_model_1.n0956 [76], RD_xram_7[4]);
  buf(\xm8051_golden_model_1.n0956 [77], RD_xram_7[5]);
  buf(\xm8051_golden_model_1.n0956 [78], RD_xram_7[6]);
  buf(\xm8051_golden_model_1.n0956 [79], RD_xram_7[7]);
  buf(\xm8051_golden_model_1.n0956 [80], RD_xram_6[0]);
  buf(\xm8051_golden_model_1.n0956 [81], RD_xram_6[1]);
  buf(\xm8051_golden_model_1.n0956 [82], RD_xram_6[2]);
  buf(\xm8051_golden_model_1.n0956 [83], RD_xram_6[3]);
  buf(\xm8051_golden_model_1.n0956 [84], RD_xram_6[4]);
  buf(\xm8051_golden_model_1.n0956 [85], RD_xram_6[5]);
  buf(\xm8051_golden_model_1.n0956 [86], RD_xram_6[6]);
  buf(\xm8051_golden_model_1.n0956 [87], RD_xram_6[7]);
  buf(\xm8051_golden_model_1.n0956 [88], RD_xram_5[0]);
  buf(\xm8051_golden_model_1.n0956 [89], RD_xram_5[1]);
  buf(\xm8051_golden_model_1.n0956 [90], RD_xram_5[2]);
  buf(\xm8051_golden_model_1.n0956 [91], RD_xram_5[3]);
  buf(\xm8051_golden_model_1.n0956 [92], RD_xram_5[4]);
  buf(\xm8051_golden_model_1.n0956 [93], RD_xram_5[5]);
  buf(\xm8051_golden_model_1.n0956 [94], RD_xram_5[6]);
  buf(\xm8051_golden_model_1.n0956 [95], RD_xram_5[7]);
  buf(\xm8051_golden_model_1.n0956 [96], RD_xram_4[0]);
  buf(\xm8051_golden_model_1.n0956 [97], RD_xram_4[1]);
  buf(\xm8051_golden_model_1.n0956 [98], RD_xram_4[2]);
  buf(\xm8051_golden_model_1.n0956 [99], RD_xram_4[3]);
  buf(\xm8051_golden_model_1.n0956 [100], RD_xram_4[4]);
  buf(\xm8051_golden_model_1.n0956 [101], RD_xram_4[5]);
  buf(\xm8051_golden_model_1.n0956 [102], RD_xram_4[6]);
  buf(\xm8051_golden_model_1.n0956 [103], RD_xram_4[7]);
  buf(\xm8051_golden_model_1.n0956 [104], RD_xram_3[0]);
  buf(\xm8051_golden_model_1.n0956 [105], RD_xram_3[1]);
  buf(\xm8051_golden_model_1.n0956 [106], RD_xram_3[2]);
  buf(\xm8051_golden_model_1.n0956 [107], RD_xram_3[3]);
  buf(\xm8051_golden_model_1.n0956 [108], RD_xram_3[4]);
  buf(\xm8051_golden_model_1.n0956 [109], RD_xram_3[5]);
  buf(\xm8051_golden_model_1.n0956 [110], RD_xram_3[6]);
  buf(\xm8051_golden_model_1.n0956 [111], RD_xram_3[7]);
  buf(\xm8051_golden_model_1.n0956 [112], RD_xram_2[0]);
  buf(\xm8051_golden_model_1.n0956 [113], RD_xram_2[1]);
  buf(\xm8051_golden_model_1.n0956 [114], RD_xram_2[2]);
  buf(\xm8051_golden_model_1.n0956 [115], RD_xram_2[3]);
  buf(\xm8051_golden_model_1.n0956 [116], RD_xram_2[4]);
  buf(\xm8051_golden_model_1.n0956 [117], RD_xram_2[5]);
  buf(\xm8051_golden_model_1.n0956 [118], RD_xram_2[6]);
  buf(\xm8051_golden_model_1.n0956 [119], RD_xram_2[7]);
  buf(\xm8051_golden_model_1.n0956 [120], RD_xram_1[0]);
  buf(\xm8051_golden_model_1.n0956 [121], RD_xram_1[1]);
  buf(\xm8051_golden_model_1.n0956 [122], RD_xram_1[2]);
  buf(\xm8051_golden_model_1.n0956 [123], RD_xram_1[3]);
  buf(\xm8051_golden_model_1.n0956 [124], RD_xram_1[4]);
  buf(\xm8051_golden_model_1.n0956 [125], RD_xram_1[5]);
  buf(\xm8051_golden_model_1.n0956 [126], RD_xram_1[6]);
  buf(\xm8051_golden_model_1.n0956 [127], RD_xram_1[7]);
  buf(\xm8051_golden_model_1.n0064 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0064 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0064 [2], \xm8051_golden_model_1.n0463 [2]);
  buf(\xm8051_golden_model_1.n0064 [3], \xm8051_golden_model_1.n0423 [3]);
  buf(\xm8051_golden_model_1.n0064 [4], \xm8051_golden_model_1.n0329 [4]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [0], proc_addr[0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [1], proc_addr[1]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [2], proc_addr[2]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [3], proc_addr[3]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [4], proc_addr[4]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [5], proc_addr[5]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [6], proc_addr[6]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [7], proc_addr[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [8], proc_addr[8]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [9], proc_addr[9]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [10], proc_addr[10]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [11], proc_addr[11]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [12], proc_addr[12]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [13], proc_addr[13]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [14], proc_addr[14]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.addr [15], proc_addr[15]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_in [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_in [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_in [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_in [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_in [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_in [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_in [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.data_in [7], proc_data_in[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.rst , rst);
  buf(\oc8051_xiommu_impl_1.sha_top_i.clk , clk);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [0], ABINPUT000[0]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [1], ABINPUT000[1]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [2], ABINPUT000[2]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [3], ABINPUT000[3]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [4], ABINPUT000[4]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [5], ABINPUT000[5]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [6], ABINPUT000[6]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [7], ABINPUT000[7]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [8], ABINPUT000[8]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [9], ABINPUT000[9]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [10], ABINPUT000[10]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [11], ABINPUT000[11]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [12], ABINPUT000[12]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [13], ABINPUT000[13]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [14], ABINPUT000[14]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [15], ABINPUT000[15]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [16], ABINPUT000[16]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [17], ABINPUT000[17]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [18], ABINPUT000[18]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [19], ABINPUT000[19]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [20], ABINPUT000[20]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [21], ABINPUT000[21]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [22], ABINPUT000[22]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [23], ABINPUT000[23]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [24], ABINPUT000[24]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [25], ABINPUT000[25]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [26], ABINPUT000[26]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [27], ABINPUT000[27]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [28], ABINPUT000[28]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [29], ABINPUT000[29]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [30], ABINPUT000[30]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [31], ABINPUT000[31]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [32], ABINPUT000[32]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [33], ABINPUT000[33]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [34], ABINPUT000[34]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [35], ABINPUT000[35]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [36], ABINPUT000[36]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [37], ABINPUT000[37]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [38], ABINPUT000[38]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [39], ABINPUT000[39]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [40], ABINPUT000[40]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [41], ABINPUT000[41]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [42], ABINPUT000[42]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [43], ABINPUT000[43]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [44], ABINPUT000[44]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [45], ABINPUT000[45]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [46], ABINPUT000[46]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [47], ABINPUT000[47]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [48], ABINPUT000[48]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [49], ABINPUT000[49]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [50], ABINPUT000[50]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [51], ABINPUT000[51]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [52], ABINPUT000[52]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [53], ABINPUT000[53]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [54], ABINPUT000[54]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [55], ABINPUT000[55]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [56], ABINPUT000[56]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [57], ABINPUT000[57]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [58], ABINPUT000[58]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [59], ABINPUT000[59]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [60], ABINPUT000[60]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [61], ABINPUT000[61]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [62], ABINPUT000[62]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [63], ABINPUT000[63]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [64], ABINPUT000[64]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [65], ABINPUT000[65]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [66], ABINPUT000[66]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [67], ABINPUT000[67]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [68], ABINPUT000[68]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [69], ABINPUT000[69]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [70], ABINPUT000[70]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [71], ABINPUT000[71]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [72], ABINPUT000[72]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [73], ABINPUT000[73]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [74], ABINPUT000[74]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [75], ABINPUT000[75]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [76], ABINPUT000[76]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [77], ABINPUT000[77]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [78], ABINPUT000[78]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [79], ABINPUT000[79]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [80], ABINPUT000[80]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [81], ABINPUT000[81]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [82], ABINPUT000[82]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [83], ABINPUT000[83]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [84], ABINPUT000[84]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [85], ABINPUT000[85]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [86], ABINPUT000[86]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [87], ABINPUT000[87]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [88], ABINPUT000[88]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [89], ABINPUT000[89]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [90], ABINPUT000[90]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [91], ABINPUT000[91]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [92], ABINPUT000[92]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [93], ABINPUT000[93]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [94], ABINPUT000[94]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [95], ABINPUT000[95]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [96], ABINPUT000[96]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [97], ABINPUT000[97]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [98], ABINPUT000[98]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [99], ABINPUT000[99]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [100], ABINPUT000[100]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [101], ABINPUT000[101]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [102], ABINPUT000[102]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [103], ABINPUT000[103]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [104], ABINPUT000[104]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [105], ABINPUT000[105]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [106], ABINPUT000[106]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [107], ABINPUT000[107]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [108], ABINPUT000[108]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [109], ABINPUT000[109]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [110], ABINPUT000[110]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [111], ABINPUT000[111]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [112], ABINPUT000[112]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [113], ABINPUT000[113]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [114], ABINPUT000[114]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [115], ABINPUT000[115]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [116], ABINPUT000[116]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [117], ABINPUT000[117]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [118], ABINPUT000[118]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [119], ABINPUT000[119]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [120], ABINPUT000[120]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [121], ABINPUT000[121]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [122], ABINPUT000[122]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [123], ABINPUT000[123]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [124], ABINPUT000[124]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [125], ABINPUT000[125]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [126], ABINPUT000[126]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [127], ABINPUT000[127]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [128], ABINPUT000[128]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [129], ABINPUT000[129]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [130], ABINPUT000[130]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [131], ABINPUT000[131]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [132], ABINPUT000[132]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [133], ABINPUT000[133]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [134], ABINPUT000[134]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [135], ABINPUT000[135]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [136], ABINPUT000[136]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [137], ABINPUT000[137]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [138], ABINPUT000[138]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [139], ABINPUT000[139]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [140], ABINPUT000[140]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [141], ABINPUT000[141]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [142], ABINPUT000[142]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [143], ABINPUT000[143]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [144], ABINPUT000[144]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [145], ABINPUT000[145]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [146], ABINPUT000[146]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [147], ABINPUT000[147]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [148], ABINPUT000[148]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [149], ABINPUT000[149]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [150], ABINPUT000[150]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [151], ABINPUT000[151]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [152], ABINPUT000[152]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [153], ABINPUT000[153]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [154], ABINPUT000[154]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [155], ABINPUT000[155]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [156], ABINPUT000[156]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [157], ABINPUT000[157]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [158], ABINPUT000[158]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [159], ABINPUT000[159]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [160], ABINPUT000[160]);
  buf(\oc8051_xiommu_impl_1.sha_top_i.ABINPUT [161], ABINPUT000[161]);
  buf(\xm8051_golden_model_1.n0055 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0055 [1], \xm8051_golden_model_1.n0187 [1]);
  buf(\xm8051_golden_model_1.n0055 [2], \xm8051_golden_model_1.n0143 [2]);
  buf(\xm8051_golden_model_1.n1305 [0], input_sha_func_55[0]);
  buf(\xm8051_golden_model_1.n1305 [1], input_sha_func_55[1]);
  buf(\xm8051_golden_model_1.n1305 [2], input_sha_func_55[2]);
  buf(\xm8051_golden_model_1.n1305 [3], input_sha_func_55[3]);
  buf(\xm8051_golden_model_1.n1305 [4], input_sha_func_55[4]);
  buf(\xm8051_golden_model_1.n1305 [5], input_sha_func_55[5]);
  buf(\xm8051_golden_model_1.n1305 [6], input_sha_func_55[6]);
  buf(\xm8051_golden_model_1.n1305 [7], input_sha_func_55[7]);
  buf(\xm8051_golden_model_1.n1305 [8], input_sha_func_55[8]);
  buf(\xm8051_golden_model_1.n1305 [9], input_sha_func_55[9]);
  buf(\xm8051_golden_model_1.n1305 [10], input_sha_func_55[10]);
  buf(\xm8051_golden_model_1.n1305 [11], input_sha_func_55[11]);
  buf(\xm8051_golden_model_1.n1305 [12], input_sha_func_55[12]);
  buf(\xm8051_golden_model_1.n1305 [13], input_sha_func_55[13]);
  buf(\xm8051_golden_model_1.n1305 [14], input_sha_func_55[14]);
  buf(\xm8051_golden_model_1.n1305 [15], input_sha_func_55[15]);
  buf(\xm8051_golden_model_1.n1305 [16], input_sha_func_55[16]);
  buf(\xm8051_golden_model_1.n1305 [17], input_sha_func_55[17]);
  buf(\xm8051_golden_model_1.n1305 [18], input_sha_func_55[18]);
  buf(\xm8051_golden_model_1.n1305 [19], input_sha_func_55[19]);
  buf(\xm8051_golden_model_1.n1305 [20], input_sha_func_55[20]);
  buf(\xm8051_golden_model_1.n1305 [21], input_sha_func_55[21]);
  buf(\xm8051_golden_model_1.n1305 [22], input_sha_func_55[22]);
  buf(\xm8051_golden_model_1.n1305 [23], input_sha_func_55[23]);
  buf(\xm8051_golden_model_1.n1305 [24], input_sha_func_55[24]);
  buf(\xm8051_golden_model_1.n1305 [25], input_sha_func_55[25]);
  buf(\xm8051_golden_model_1.n1305 [26], input_sha_func_55[26]);
  buf(\xm8051_golden_model_1.n1305 [27], input_sha_func_55[27]);
  buf(\xm8051_golden_model_1.n1305 [28], input_sha_func_55[28]);
  buf(\xm8051_golden_model_1.n1305 [29], input_sha_func_55[29]);
  buf(\xm8051_golden_model_1.n1305 [30], input_sha_func_55[30]);
  buf(\xm8051_golden_model_1.n1305 [31], input_sha_func_55[31]);
  buf(\xm8051_golden_model_1.n1305 [32], input_sha_func_54[0]);
  buf(\xm8051_golden_model_1.n1305 [33], input_sha_func_54[1]);
  buf(\xm8051_golden_model_1.n1305 [34], input_sha_func_54[2]);
  buf(\xm8051_golden_model_1.n1305 [35], input_sha_func_54[3]);
  buf(\xm8051_golden_model_1.n1305 [36], input_sha_func_54[4]);
  buf(\xm8051_golden_model_1.n1305 [37], input_sha_func_54[5]);
  buf(\xm8051_golden_model_1.n1305 [38], input_sha_func_54[6]);
  buf(\xm8051_golden_model_1.n1305 [39], input_sha_func_54[7]);
  buf(\xm8051_golden_model_1.n1305 [40], input_sha_func_54[8]);
  buf(\xm8051_golden_model_1.n1305 [41], input_sha_func_54[9]);
  buf(\xm8051_golden_model_1.n1305 [42], input_sha_func_54[10]);
  buf(\xm8051_golden_model_1.n1305 [43], input_sha_func_54[11]);
  buf(\xm8051_golden_model_1.n1305 [44], input_sha_func_54[12]);
  buf(\xm8051_golden_model_1.n1305 [45], input_sha_func_54[13]);
  buf(\xm8051_golden_model_1.n1305 [46], input_sha_func_54[14]);
  buf(\xm8051_golden_model_1.n1305 [47], input_sha_func_54[15]);
  buf(\xm8051_golden_model_1.n1305 [48], input_sha_func_54[16]);
  buf(\xm8051_golden_model_1.n1305 [49], input_sha_func_54[17]);
  buf(\xm8051_golden_model_1.n1305 [50], input_sha_func_54[18]);
  buf(\xm8051_golden_model_1.n1305 [51], input_sha_func_54[19]);
  buf(\xm8051_golden_model_1.n1305 [52], input_sha_func_54[20]);
  buf(\xm8051_golden_model_1.n1305 [53], input_sha_func_54[21]);
  buf(\xm8051_golden_model_1.n1305 [54], input_sha_func_54[22]);
  buf(\xm8051_golden_model_1.n1305 [55], input_sha_func_54[23]);
  buf(\xm8051_golden_model_1.n1305 [56], input_sha_func_54[24]);
  buf(\xm8051_golden_model_1.n1305 [57], input_sha_func_54[25]);
  buf(\xm8051_golden_model_1.n1305 [58], input_sha_func_54[26]);
  buf(\xm8051_golden_model_1.n1305 [59], input_sha_func_54[27]);
  buf(\xm8051_golden_model_1.n1305 [60], input_sha_func_54[28]);
  buf(\xm8051_golden_model_1.n1305 [61], input_sha_func_54[29]);
  buf(\xm8051_golden_model_1.n1305 [62], input_sha_func_54[30]);
  buf(\xm8051_golden_model_1.n1305 [63], input_sha_func_54[31]);
  buf(\xm8051_golden_model_1.n1305 [64], input_sha_func_54[32]);
  buf(\xm8051_golden_model_1.n1305 [65], input_sha_func_54[33]);
  buf(\xm8051_golden_model_1.n1305 [66], input_sha_func_54[34]);
  buf(\xm8051_golden_model_1.n1305 [67], input_sha_func_54[35]);
  buf(\xm8051_golden_model_1.n1305 [68], input_sha_func_54[36]);
  buf(\xm8051_golden_model_1.n1305 [69], input_sha_func_54[37]);
  buf(\xm8051_golden_model_1.n1305 [70], input_sha_func_54[38]);
  buf(\xm8051_golden_model_1.n1305 [71], input_sha_func_54[39]);
  buf(\xm8051_golden_model_1.n1305 [72], input_sha_func_54[40]);
  buf(\xm8051_golden_model_1.n1305 [73], input_sha_func_54[41]);
  buf(\xm8051_golden_model_1.n1305 [74], input_sha_func_54[42]);
  buf(\xm8051_golden_model_1.n1305 [75], input_sha_func_54[43]);
  buf(\xm8051_golden_model_1.n1305 [76], input_sha_func_54[44]);
  buf(\xm8051_golden_model_1.n1305 [77], input_sha_func_54[45]);
  buf(\xm8051_golden_model_1.n1305 [78], input_sha_func_54[46]);
  buf(\xm8051_golden_model_1.n1305 [79], input_sha_func_54[47]);
  buf(\xm8051_golden_model_1.n1305 [80], input_sha_func_54[48]);
  buf(\xm8051_golden_model_1.n1305 [81], input_sha_func_54[49]);
  buf(\xm8051_golden_model_1.n1305 [82], input_sha_func_54[50]);
  buf(\xm8051_golden_model_1.n1305 [83], input_sha_func_54[51]);
  buf(\xm8051_golden_model_1.n1305 [84], input_sha_func_54[52]);
  buf(\xm8051_golden_model_1.n1305 [85], input_sha_func_54[53]);
  buf(\xm8051_golden_model_1.n1305 [86], input_sha_func_54[54]);
  buf(\xm8051_golden_model_1.n1305 [87], input_sha_func_54[55]);
  buf(\xm8051_golden_model_1.n1305 [88], input_sha_func_54[56]);
  buf(\xm8051_golden_model_1.n1305 [89], input_sha_func_54[57]);
  buf(\xm8051_golden_model_1.n1305 [90], input_sha_func_54[58]);
  buf(\xm8051_golden_model_1.n1305 [91], input_sha_func_54[59]);
  buf(\xm8051_golden_model_1.n1305 [92], input_sha_func_54[60]);
  buf(\xm8051_golden_model_1.n1305 [93], input_sha_func_54[61]);
  buf(\xm8051_golden_model_1.n1305 [94], input_sha_func_54[62]);
  buf(\xm8051_golden_model_1.n1305 [95], input_sha_func_54[63]);
  buf(\xm8051_golden_model_1.n1305 [96], input_sha_func_53[0]);
  buf(\xm8051_golden_model_1.n1305 [97], input_sha_func_53[1]);
  buf(\xm8051_golden_model_1.n1305 [98], input_sha_func_53[2]);
  buf(\xm8051_golden_model_1.n1305 [99], input_sha_func_53[3]);
  buf(\xm8051_golden_model_1.n1305 [100], input_sha_func_53[4]);
  buf(\xm8051_golden_model_1.n1305 [101], input_sha_func_53[5]);
  buf(\xm8051_golden_model_1.n1305 [102], input_sha_func_53[6]);
  buf(\xm8051_golden_model_1.n1305 [103], input_sha_func_53[7]);
  buf(\xm8051_golden_model_1.n1305 [104], input_sha_func_53[8]);
  buf(\xm8051_golden_model_1.n1305 [105], input_sha_func_53[9]);
  buf(\xm8051_golden_model_1.n1305 [106], input_sha_func_53[10]);
  buf(\xm8051_golden_model_1.n1305 [107], input_sha_func_53[11]);
  buf(\xm8051_golden_model_1.n1305 [108], input_sha_func_53[12]);
  buf(\xm8051_golden_model_1.n1305 [109], input_sha_func_53[13]);
  buf(\xm8051_golden_model_1.n1305 [110], input_sha_func_53[14]);
  buf(\xm8051_golden_model_1.n1305 [111], input_sha_func_53[15]);
  buf(\xm8051_golden_model_1.n1305 [112], input_sha_func_53[16]);
  buf(\xm8051_golden_model_1.n1305 [113], input_sha_func_53[17]);
  buf(\xm8051_golden_model_1.n1305 [114], input_sha_func_53[18]);
  buf(\xm8051_golden_model_1.n1305 [115], input_sha_func_53[19]);
  buf(\xm8051_golden_model_1.n1305 [116], input_sha_func_53[20]);
  buf(\xm8051_golden_model_1.n1305 [117], input_sha_func_53[21]);
  buf(\xm8051_golden_model_1.n1305 [118], input_sha_func_53[22]);
  buf(\xm8051_golden_model_1.n1305 [119], input_sha_func_53[23]);
  buf(\xm8051_golden_model_1.n1305 [120], input_sha_func_53[24]);
  buf(\xm8051_golden_model_1.n1305 [121], input_sha_func_53[25]);
  buf(\xm8051_golden_model_1.n1305 [122], input_sha_func_53[26]);
  buf(\xm8051_golden_model_1.n1305 [123], input_sha_func_53[27]);
  buf(\xm8051_golden_model_1.n1305 [124], input_sha_func_53[28]);
  buf(\xm8051_golden_model_1.n1305 [125], input_sha_func_53[29]);
  buf(\xm8051_golden_model_1.n1305 [126], input_sha_func_53[30]);
  buf(\xm8051_golden_model_1.n1305 [127], input_sha_func_53[31]);
  buf(\xm8051_golden_model_1.n1305 [128], input_sha_func_53[32]);
  buf(\xm8051_golden_model_1.n1305 [129], input_sha_func_53[33]);
  buf(\xm8051_golden_model_1.n1305 [130], input_sha_func_53[34]);
  buf(\xm8051_golden_model_1.n1305 [131], input_sha_func_53[35]);
  buf(\xm8051_golden_model_1.n1305 [132], input_sha_func_53[36]);
  buf(\xm8051_golden_model_1.n1305 [133], input_sha_func_53[37]);
  buf(\xm8051_golden_model_1.n1305 [134], input_sha_func_53[38]);
  buf(\xm8051_golden_model_1.n1305 [135], input_sha_func_53[39]);
  buf(\xm8051_golden_model_1.n1305 [136], input_sha_func_53[40]);
  buf(\xm8051_golden_model_1.n1305 [137], input_sha_func_53[41]);
  buf(\xm8051_golden_model_1.n1305 [138], input_sha_func_53[42]);
  buf(\xm8051_golden_model_1.n1305 [139], input_sha_func_53[43]);
  buf(\xm8051_golden_model_1.n1305 [140], input_sha_func_53[44]);
  buf(\xm8051_golden_model_1.n1305 [141], input_sha_func_53[45]);
  buf(\xm8051_golden_model_1.n1305 [142], input_sha_func_53[46]);
  buf(\xm8051_golden_model_1.n1305 [143], input_sha_func_53[47]);
  buf(\xm8051_golden_model_1.n1305 [144], input_sha_func_53[48]);
  buf(\xm8051_golden_model_1.n1305 [145], input_sha_func_53[49]);
  buf(\xm8051_golden_model_1.n1305 [146], input_sha_func_53[50]);
  buf(\xm8051_golden_model_1.n1305 [147], input_sha_func_53[51]);
  buf(\xm8051_golden_model_1.n1305 [148], input_sha_func_53[52]);
  buf(\xm8051_golden_model_1.n1305 [149], input_sha_func_53[53]);
  buf(\xm8051_golden_model_1.n1305 [150], input_sha_func_53[54]);
  buf(\xm8051_golden_model_1.n1305 [151], input_sha_func_53[55]);
  buf(\xm8051_golden_model_1.n1305 [152], input_sha_func_53[56]);
  buf(\xm8051_golden_model_1.n1305 [153], input_sha_func_53[57]);
  buf(\xm8051_golden_model_1.n1305 [154], input_sha_func_53[58]);
  buf(\xm8051_golden_model_1.n1305 [155], input_sha_func_53[59]);
  buf(\xm8051_golden_model_1.n1305 [156], input_sha_func_53[60]);
  buf(\xm8051_golden_model_1.n1305 [157], input_sha_func_53[61]);
  buf(\xm8051_golden_model_1.n1305 [158], input_sha_func_53[62]);
  buf(\xm8051_golden_model_1.n1305 [159], input_sha_func_53[63]);
  buf(\xm8051_golden_model_1.n1303 [0], input_aes_func_52[0]);
  buf(\xm8051_golden_model_1.n1303 [1], input_aes_func_52[1]);
  buf(\xm8051_golden_model_1.n1303 [2], input_aes_func_52[2]);
  buf(\xm8051_golden_model_1.n1303 [3], input_aes_func_52[3]);
  buf(\xm8051_golden_model_1.n1303 [4], input_aes_func_52[4]);
  buf(\xm8051_golden_model_1.n1303 [5], input_aes_func_52[5]);
  buf(\xm8051_golden_model_1.n1303 [6], input_aes_func_52[6]);
  buf(\xm8051_golden_model_1.n1303 [7], input_aes_func_52[7]);
  buf(\xm8051_golden_model_1.n1303 [8], input_aes_func_52[8]);
  buf(\xm8051_golden_model_1.n1303 [9], input_aes_func_52[9]);
  buf(\xm8051_golden_model_1.n1303 [10], input_aes_func_52[10]);
  buf(\xm8051_golden_model_1.n1303 [11], input_aes_func_52[11]);
  buf(\xm8051_golden_model_1.n1303 [12], input_aes_func_52[12]);
  buf(\xm8051_golden_model_1.n1303 [13], input_aes_func_52[13]);
  buf(\xm8051_golden_model_1.n1303 [14], input_aes_func_52[14]);
  buf(\xm8051_golden_model_1.n1303 [15], input_aes_func_52[15]);
  buf(\xm8051_golden_model_1.n1303 [16], input_aes_func_52[16]);
  buf(\xm8051_golden_model_1.n1303 [17], input_aes_func_52[17]);
  buf(\xm8051_golden_model_1.n1303 [18], input_aes_func_52[18]);
  buf(\xm8051_golden_model_1.n1303 [19], input_aes_func_52[19]);
  buf(\xm8051_golden_model_1.n1303 [20], input_aes_func_52[20]);
  buf(\xm8051_golden_model_1.n1303 [21], input_aes_func_52[21]);
  buf(\xm8051_golden_model_1.n1303 [22], input_aes_func_52[22]);
  buf(\xm8051_golden_model_1.n1303 [23], input_aes_func_52[23]);
  buf(\xm8051_golden_model_1.n1303 [24], input_aes_func_52[24]);
  buf(\xm8051_golden_model_1.n1303 [25], input_aes_func_52[25]);
  buf(\xm8051_golden_model_1.n1303 [26], input_aes_func_52[26]);
  buf(\xm8051_golden_model_1.n1303 [27], input_aes_func_52[27]);
  buf(\xm8051_golden_model_1.n1303 [28], input_aes_func_52[28]);
  buf(\xm8051_golden_model_1.n1303 [29], input_aes_func_52[29]);
  buf(\xm8051_golden_model_1.n1303 [30], input_aes_func_52[30]);
  buf(\xm8051_golden_model_1.n1303 [31], input_aes_func_52[31]);
  buf(\xm8051_golden_model_1.n1303 [32], input_aes_func_52[32]);
  buf(\xm8051_golden_model_1.n1303 [33], input_aes_func_52[33]);
  buf(\xm8051_golden_model_1.n1303 [34], input_aes_func_52[34]);
  buf(\xm8051_golden_model_1.n1303 [35], input_aes_func_52[35]);
  buf(\xm8051_golden_model_1.n1303 [36], input_aes_func_52[36]);
  buf(\xm8051_golden_model_1.n1303 [37], input_aes_func_52[37]);
  buf(\xm8051_golden_model_1.n1303 [38], input_aes_func_52[38]);
  buf(\xm8051_golden_model_1.n1303 [39], input_aes_func_52[39]);
  buf(\xm8051_golden_model_1.n1303 [40], input_aes_func_52[40]);
  buf(\xm8051_golden_model_1.n1303 [41], input_aes_func_52[41]);
  buf(\xm8051_golden_model_1.n1303 [42], input_aes_func_52[42]);
  buf(\xm8051_golden_model_1.n1303 [43], input_aes_func_52[43]);
  buf(\xm8051_golden_model_1.n1303 [44], input_aes_func_52[44]);
  buf(\xm8051_golden_model_1.n1303 [45], input_aes_func_52[45]);
  buf(\xm8051_golden_model_1.n1303 [46], input_aes_func_52[46]);
  buf(\xm8051_golden_model_1.n1303 [47], input_aes_func_52[47]);
  buf(\xm8051_golden_model_1.n1303 [48], input_aes_func_52[48]);
  buf(\xm8051_golden_model_1.n1303 [49], input_aes_func_52[49]);
  buf(\xm8051_golden_model_1.n1303 [50], input_aes_func_52[50]);
  buf(\xm8051_golden_model_1.n1303 [51], input_aes_func_52[51]);
  buf(\xm8051_golden_model_1.n1303 [52], input_aes_func_52[52]);
  buf(\xm8051_golden_model_1.n1303 [53], input_aes_func_52[53]);
  buf(\xm8051_golden_model_1.n1303 [54], input_aes_func_52[54]);
  buf(\xm8051_golden_model_1.n1303 [55], input_aes_func_52[55]);
  buf(\xm8051_golden_model_1.n1303 [56], input_aes_func_52[56]);
  buf(\xm8051_golden_model_1.n1303 [57], input_aes_func_52[57]);
  buf(\xm8051_golden_model_1.n1303 [58], input_aes_func_52[58]);
  buf(\xm8051_golden_model_1.n1303 [59], input_aes_func_52[59]);
  buf(\xm8051_golden_model_1.n1303 [60], input_aes_func_52[60]);
  buf(\xm8051_golden_model_1.n1303 [61], input_aes_func_52[61]);
  buf(\xm8051_golden_model_1.n1303 [62], input_aes_func_52[62]);
  buf(\xm8051_golden_model_1.n1303 [63], input_aes_func_52[63]);
  buf(\xm8051_golden_model_1.n1303 [64], input_aes_func_51[0]);
  buf(\xm8051_golden_model_1.n1303 [65], input_aes_func_51[1]);
  buf(\xm8051_golden_model_1.n1303 [66], input_aes_func_51[2]);
  buf(\xm8051_golden_model_1.n1303 [67], input_aes_func_51[3]);
  buf(\xm8051_golden_model_1.n1303 [68], input_aes_func_51[4]);
  buf(\xm8051_golden_model_1.n1303 [69], input_aes_func_51[5]);
  buf(\xm8051_golden_model_1.n1303 [70], input_aes_func_51[6]);
  buf(\xm8051_golden_model_1.n1303 [71], input_aes_func_51[7]);
  buf(\xm8051_golden_model_1.n1303 [72], input_aes_func_51[8]);
  buf(\xm8051_golden_model_1.n1303 [73], input_aes_func_51[9]);
  buf(\xm8051_golden_model_1.n1303 [74], input_aes_func_51[10]);
  buf(\xm8051_golden_model_1.n1303 [75], input_aes_func_51[11]);
  buf(\xm8051_golden_model_1.n1303 [76], input_aes_func_51[12]);
  buf(\xm8051_golden_model_1.n1303 [77], input_aes_func_51[13]);
  buf(\xm8051_golden_model_1.n1303 [78], input_aes_func_51[14]);
  buf(\xm8051_golden_model_1.n1303 [79], input_aes_func_51[15]);
  buf(\xm8051_golden_model_1.n1303 [80], input_aes_func_51[16]);
  buf(\xm8051_golden_model_1.n1303 [81], input_aes_func_51[17]);
  buf(\xm8051_golden_model_1.n1303 [82], input_aes_func_51[18]);
  buf(\xm8051_golden_model_1.n1303 [83], input_aes_func_51[19]);
  buf(\xm8051_golden_model_1.n1303 [84], input_aes_func_51[20]);
  buf(\xm8051_golden_model_1.n1303 [85], input_aes_func_51[21]);
  buf(\xm8051_golden_model_1.n1303 [86], input_aes_func_51[22]);
  buf(\xm8051_golden_model_1.n1303 [87], input_aes_func_51[23]);
  buf(\xm8051_golden_model_1.n1303 [88], input_aes_func_51[24]);
  buf(\xm8051_golden_model_1.n1303 [89], input_aes_func_51[25]);
  buf(\xm8051_golden_model_1.n1303 [90], input_aes_func_51[26]);
  buf(\xm8051_golden_model_1.n1303 [91], input_aes_func_51[27]);
  buf(\xm8051_golden_model_1.n1303 [92], input_aes_func_51[28]);
  buf(\xm8051_golden_model_1.n1303 [93], input_aes_func_51[29]);
  buf(\xm8051_golden_model_1.n1303 [94], input_aes_func_51[30]);
  buf(\xm8051_golden_model_1.n1303 [95], input_aes_func_51[31]);
  buf(\xm8051_golden_model_1.n1303 [96], input_aes_func_51[32]);
  buf(\xm8051_golden_model_1.n1303 [97], input_aes_func_51[33]);
  buf(\xm8051_golden_model_1.n1303 [98], input_aes_func_51[34]);
  buf(\xm8051_golden_model_1.n1303 [99], input_aes_func_51[35]);
  buf(\xm8051_golden_model_1.n1303 [100], input_aes_func_51[36]);
  buf(\xm8051_golden_model_1.n1303 [101], input_aes_func_51[37]);
  buf(\xm8051_golden_model_1.n1303 [102], input_aes_func_51[38]);
  buf(\xm8051_golden_model_1.n1303 [103], input_aes_func_51[39]);
  buf(\xm8051_golden_model_1.n1303 [104], input_aes_func_51[40]);
  buf(\xm8051_golden_model_1.n1303 [105], input_aes_func_51[41]);
  buf(\xm8051_golden_model_1.n1303 [106], input_aes_func_51[42]);
  buf(\xm8051_golden_model_1.n1303 [107], input_aes_func_51[43]);
  buf(\xm8051_golden_model_1.n1303 [108], input_aes_func_51[44]);
  buf(\xm8051_golden_model_1.n1303 [109], input_aes_func_51[45]);
  buf(\xm8051_golden_model_1.n1303 [110], input_aes_func_51[46]);
  buf(\xm8051_golden_model_1.n1303 [111], input_aes_func_51[47]);
  buf(\xm8051_golden_model_1.n1303 [112], input_aes_func_51[48]);
  buf(\xm8051_golden_model_1.n1303 [113], input_aes_func_51[49]);
  buf(\xm8051_golden_model_1.n1303 [114], input_aes_func_51[50]);
  buf(\xm8051_golden_model_1.n1303 [115], input_aes_func_51[51]);
  buf(\xm8051_golden_model_1.n1303 [116], input_aes_func_51[52]);
  buf(\xm8051_golden_model_1.n1303 [117], input_aes_func_51[53]);
  buf(\xm8051_golden_model_1.n1303 [118], input_aes_func_51[54]);
  buf(\xm8051_golden_model_1.n1303 [119], input_aes_func_51[55]);
  buf(\xm8051_golden_model_1.n1303 [120], input_aes_func_51[56]);
  buf(\xm8051_golden_model_1.n1303 [121], input_aes_func_51[57]);
  buf(\xm8051_golden_model_1.n1303 [122], input_aes_func_51[58]);
  buf(\xm8051_golden_model_1.n1303 [123], input_aes_func_51[59]);
  buf(\xm8051_golden_model_1.n1303 [124], input_aes_func_51[60]);
  buf(\xm8051_golden_model_1.n1303 [125], input_aes_func_51[61]);
  buf(\xm8051_golden_model_1.n1303 [126], input_aes_func_51[62]);
  buf(\xm8051_golden_model_1.n1303 [127], input_aes_func_51[63]);
  buf(\xm8051_golden_model_1.n0532 [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.n0532 [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.n0532 [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.n0532 [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.n0529 [0], 1'b0);
  buf(\xm8051_golden_model_1.n0529 [1], 1'b0);
  buf(\xm8051_golden_model_1.n0529 [2], 1'b0);
  buf(\xm8051_golden_model_1.n0529 [3], 1'b0);
  buf(\xm8051_golden_model_1.n0529 [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.n0529 [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.n0529 [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.n0529 [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.n0529 [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.n0529 [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.n0529 [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.n0529 [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.n0529 [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.n0529 [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.n0529 [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.n0529 [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.n0527 [0], proc_addr[4]);
  buf(\xm8051_golden_model_1.n0527 [1], proc_addr[5]);
  buf(\xm8051_golden_model_1.n0527 [2], proc_addr[6]);
  buf(\xm8051_golden_model_1.n0527 [3], proc_addr[7]);
  buf(\xm8051_golden_model_1.n0527 [4], proc_addr[8]);
  buf(\xm8051_golden_model_1.n0527 [5], proc_addr[9]);
  buf(\xm8051_golden_model_1.n0527 [6], proc_addr[10]);
  buf(\xm8051_golden_model_1.n0527 [7], proc_addr[11]);
  buf(\xm8051_golden_model_1.n0527 [8], proc_addr[12]);
  buf(\xm8051_golden_model_1.n0527 [9], proc_addr[13]);
  buf(\xm8051_golden_model_1.n0527 [10], proc_addr[14]);
  buf(\xm8051_golden_model_1.n0527 [11], proc_addr[15]);
  buf(\xm8051_golden_model_1.n0037 [0], proc_addr[0]);
  buf(\xm8051_golden_model_1.n0037 [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.n0037 [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.n0037 [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.n0037 [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.n0037 [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.n0037 [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.n0037 [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.n0037 [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.n0037 [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.n0037 [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.n0037 [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.n0037 [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.n0037 [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.n0037 [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.n0037 [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.n1299 [0], input_sha_func_50[0]);
  buf(\xm8051_golden_model_1.n1299 [1], input_sha_func_50[1]);
  buf(\xm8051_golden_model_1.n1299 [2], input_sha_func_50[2]);
  buf(\xm8051_golden_model_1.n1299 [3], input_sha_func_50[3]);
  buf(\xm8051_golden_model_1.n1299 [4], input_sha_func_50[4]);
  buf(\xm8051_golden_model_1.n1299 [5], input_sha_func_50[5]);
  buf(\xm8051_golden_model_1.n1299 [6], input_sha_func_50[6]);
  buf(\xm8051_golden_model_1.n1299 [7], input_sha_func_50[7]);
  buf(\xm8051_golden_model_1.n1299 [8], input_sha_func_50[8]);
  buf(\xm8051_golden_model_1.n1299 [9], input_sha_func_50[9]);
  buf(\xm8051_golden_model_1.n1299 [10], input_sha_func_50[10]);
  buf(\xm8051_golden_model_1.n1299 [11], input_sha_func_50[11]);
  buf(\xm8051_golden_model_1.n1299 [12], input_sha_func_50[12]);
  buf(\xm8051_golden_model_1.n1299 [13], input_sha_func_50[13]);
  buf(\xm8051_golden_model_1.n1299 [14], input_sha_func_50[14]);
  buf(\xm8051_golden_model_1.n1299 [15], input_sha_func_50[15]);
  buf(\xm8051_golden_model_1.n1299 [16], input_sha_func_50[16]);
  buf(\xm8051_golden_model_1.n1299 [17], input_sha_func_50[17]);
  buf(\xm8051_golden_model_1.n1299 [18], input_sha_func_50[18]);
  buf(\xm8051_golden_model_1.n1299 [19], input_sha_func_50[19]);
  buf(\xm8051_golden_model_1.n1299 [20], input_sha_func_50[20]);
  buf(\xm8051_golden_model_1.n1299 [21], input_sha_func_50[21]);
  buf(\xm8051_golden_model_1.n1299 [22], input_sha_func_50[22]);
  buf(\xm8051_golden_model_1.n1299 [23], input_sha_func_50[23]);
  buf(\xm8051_golden_model_1.n1299 [24], input_sha_func_50[24]);
  buf(\xm8051_golden_model_1.n1299 [25], input_sha_func_50[25]);
  buf(\xm8051_golden_model_1.n1299 [26], input_sha_func_50[26]);
  buf(\xm8051_golden_model_1.n1299 [27], input_sha_func_50[27]);
  buf(\xm8051_golden_model_1.n1299 [28], input_sha_func_50[28]);
  buf(\xm8051_golden_model_1.n1299 [29], input_sha_func_50[29]);
  buf(\xm8051_golden_model_1.n1299 [30], input_sha_func_50[30]);
  buf(\xm8051_golden_model_1.n1299 [31], input_sha_func_50[31]);
  buf(\xm8051_golden_model_1.n1299 [32], input_sha_func_49[0]);
  buf(\xm8051_golden_model_1.n1299 [33], input_sha_func_49[1]);
  buf(\xm8051_golden_model_1.n1299 [34], input_sha_func_49[2]);
  buf(\xm8051_golden_model_1.n1299 [35], input_sha_func_49[3]);
  buf(\xm8051_golden_model_1.n1299 [36], input_sha_func_49[4]);
  buf(\xm8051_golden_model_1.n1299 [37], input_sha_func_49[5]);
  buf(\xm8051_golden_model_1.n1299 [38], input_sha_func_49[6]);
  buf(\xm8051_golden_model_1.n1299 [39], input_sha_func_49[7]);
  buf(\xm8051_golden_model_1.n1299 [40], input_sha_func_49[8]);
  buf(\xm8051_golden_model_1.n1299 [41], input_sha_func_49[9]);
  buf(\xm8051_golden_model_1.n1299 [42], input_sha_func_49[10]);
  buf(\xm8051_golden_model_1.n1299 [43], input_sha_func_49[11]);
  buf(\xm8051_golden_model_1.n1299 [44], input_sha_func_49[12]);
  buf(\xm8051_golden_model_1.n1299 [45], input_sha_func_49[13]);
  buf(\xm8051_golden_model_1.n1299 [46], input_sha_func_49[14]);
  buf(\xm8051_golden_model_1.n1299 [47], input_sha_func_49[15]);
  buf(\xm8051_golden_model_1.n1299 [48], input_sha_func_49[16]);
  buf(\xm8051_golden_model_1.n1299 [49], input_sha_func_49[17]);
  buf(\xm8051_golden_model_1.n1299 [50], input_sha_func_49[18]);
  buf(\xm8051_golden_model_1.n1299 [51], input_sha_func_49[19]);
  buf(\xm8051_golden_model_1.n1299 [52], input_sha_func_49[20]);
  buf(\xm8051_golden_model_1.n1299 [53], input_sha_func_49[21]);
  buf(\xm8051_golden_model_1.n1299 [54], input_sha_func_49[22]);
  buf(\xm8051_golden_model_1.n1299 [55], input_sha_func_49[23]);
  buf(\xm8051_golden_model_1.n1299 [56], input_sha_func_49[24]);
  buf(\xm8051_golden_model_1.n1299 [57], input_sha_func_49[25]);
  buf(\xm8051_golden_model_1.n1299 [58], input_sha_func_49[26]);
  buf(\xm8051_golden_model_1.n1299 [59], input_sha_func_49[27]);
  buf(\xm8051_golden_model_1.n1299 [60], input_sha_func_49[28]);
  buf(\xm8051_golden_model_1.n1299 [61], input_sha_func_49[29]);
  buf(\xm8051_golden_model_1.n1299 [62], input_sha_func_49[30]);
  buf(\xm8051_golden_model_1.n1299 [63], input_sha_func_49[31]);
  buf(\xm8051_golden_model_1.n1299 [64], input_sha_func_49[32]);
  buf(\xm8051_golden_model_1.n1299 [65], input_sha_func_49[33]);
  buf(\xm8051_golden_model_1.n1299 [66], input_sha_func_49[34]);
  buf(\xm8051_golden_model_1.n1299 [67], input_sha_func_49[35]);
  buf(\xm8051_golden_model_1.n1299 [68], input_sha_func_49[36]);
  buf(\xm8051_golden_model_1.n1299 [69], input_sha_func_49[37]);
  buf(\xm8051_golden_model_1.n1299 [70], input_sha_func_49[38]);
  buf(\xm8051_golden_model_1.n1299 [71], input_sha_func_49[39]);
  buf(\xm8051_golden_model_1.n1299 [72], input_sha_func_49[40]);
  buf(\xm8051_golden_model_1.n1299 [73], input_sha_func_49[41]);
  buf(\xm8051_golden_model_1.n1299 [74], input_sha_func_49[42]);
  buf(\xm8051_golden_model_1.n1299 [75], input_sha_func_49[43]);
  buf(\xm8051_golden_model_1.n1299 [76], input_sha_func_49[44]);
  buf(\xm8051_golden_model_1.n1299 [77], input_sha_func_49[45]);
  buf(\xm8051_golden_model_1.n1299 [78], input_sha_func_49[46]);
  buf(\xm8051_golden_model_1.n1299 [79], input_sha_func_49[47]);
  buf(\xm8051_golden_model_1.n1299 [80], input_sha_func_49[48]);
  buf(\xm8051_golden_model_1.n1299 [81], input_sha_func_49[49]);
  buf(\xm8051_golden_model_1.n1299 [82], input_sha_func_49[50]);
  buf(\xm8051_golden_model_1.n1299 [83], input_sha_func_49[51]);
  buf(\xm8051_golden_model_1.n1299 [84], input_sha_func_49[52]);
  buf(\xm8051_golden_model_1.n1299 [85], input_sha_func_49[53]);
  buf(\xm8051_golden_model_1.n1299 [86], input_sha_func_49[54]);
  buf(\xm8051_golden_model_1.n1299 [87], input_sha_func_49[55]);
  buf(\xm8051_golden_model_1.n1299 [88], input_sha_func_49[56]);
  buf(\xm8051_golden_model_1.n1299 [89], input_sha_func_49[57]);
  buf(\xm8051_golden_model_1.n1299 [90], input_sha_func_49[58]);
  buf(\xm8051_golden_model_1.n1299 [91], input_sha_func_49[59]);
  buf(\xm8051_golden_model_1.n1299 [92], input_sha_func_49[60]);
  buf(\xm8051_golden_model_1.n1299 [93], input_sha_func_49[61]);
  buf(\xm8051_golden_model_1.n1299 [94], input_sha_func_49[62]);
  buf(\xm8051_golden_model_1.n1299 [95], input_sha_func_49[63]);
  buf(\xm8051_golden_model_1.n1299 [96], input_sha_func_48[0]);
  buf(\xm8051_golden_model_1.n1299 [97], input_sha_func_48[1]);
  buf(\xm8051_golden_model_1.n1299 [98], input_sha_func_48[2]);
  buf(\xm8051_golden_model_1.n1299 [99], input_sha_func_48[3]);
  buf(\xm8051_golden_model_1.n1299 [100], input_sha_func_48[4]);
  buf(\xm8051_golden_model_1.n1299 [101], input_sha_func_48[5]);
  buf(\xm8051_golden_model_1.n1299 [102], input_sha_func_48[6]);
  buf(\xm8051_golden_model_1.n1299 [103], input_sha_func_48[7]);
  buf(\xm8051_golden_model_1.n1299 [104], input_sha_func_48[8]);
  buf(\xm8051_golden_model_1.n1299 [105], input_sha_func_48[9]);
  buf(\xm8051_golden_model_1.n1299 [106], input_sha_func_48[10]);
  buf(\xm8051_golden_model_1.n1299 [107], input_sha_func_48[11]);
  buf(\xm8051_golden_model_1.n1299 [108], input_sha_func_48[12]);
  buf(\xm8051_golden_model_1.n1299 [109], input_sha_func_48[13]);
  buf(\xm8051_golden_model_1.n1299 [110], input_sha_func_48[14]);
  buf(\xm8051_golden_model_1.n1299 [111], input_sha_func_48[15]);
  buf(\xm8051_golden_model_1.n1299 [112], input_sha_func_48[16]);
  buf(\xm8051_golden_model_1.n1299 [113], input_sha_func_48[17]);
  buf(\xm8051_golden_model_1.n1299 [114], input_sha_func_48[18]);
  buf(\xm8051_golden_model_1.n1299 [115], input_sha_func_48[19]);
  buf(\xm8051_golden_model_1.n1299 [116], input_sha_func_48[20]);
  buf(\xm8051_golden_model_1.n1299 [117], input_sha_func_48[21]);
  buf(\xm8051_golden_model_1.n1299 [118], input_sha_func_48[22]);
  buf(\xm8051_golden_model_1.n1299 [119], input_sha_func_48[23]);
  buf(\xm8051_golden_model_1.n1299 [120], input_sha_func_48[24]);
  buf(\xm8051_golden_model_1.n1299 [121], input_sha_func_48[25]);
  buf(\xm8051_golden_model_1.n1299 [122], input_sha_func_48[26]);
  buf(\xm8051_golden_model_1.n1299 [123], input_sha_func_48[27]);
  buf(\xm8051_golden_model_1.n1299 [124], input_sha_func_48[28]);
  buf(\xm8051_golden_model_1.n1299 [125], input_sha_func_48[29]);
  buf(\xm8051_golden_model_1.n1299 [126], input_sha_func_48[30]);
  buf(\xm8051_golden_model_1.n1299 [127], input_sha_func_48[31]);
  buf(\xm8051_golden_model_1.n1299 [128], input_sha_func_48[32]);
  buf(\xm8051_golden_model_1.n1299 [129], input_sha_func_48[33]);
  buf(\xm8051_golden_model_1.n1299 [130], input_sha_func_48[34]);
  buf(\xm8051_golden_model_1.n1299 [131], input_sha_func_48[35]);
  buf(\xm8051_golden_model_1.n1299 [132], input_sha_func_48[36]);
  buf(\xm8051_golden_model_1.n1299 [133], input_sha_func_48[37]);
  buf(\xm8051_golden_model_1.n1299 [134], input_sha_func_48[38]);
  buf(\xm8051_golden_model_1.n1299 [135], input_sha_func_48[39]);
  buf(\xm8051_golden_model_1.n1299 [136], input_sha_func_48[40]);
  buf(\xm8051_golden_model_1.n1299 [137], input_sha_func_48[41]);
  buf(\xm8051_golden_model_1.n1299 [138], input_sha_func_48[42]);
  buf(\xm8051_golden_model_1.n1299 [139], input_sha_func_48[43]);
  buf(\xm8051_golden_model_1.n1299 [140], input_sha_func_48[44]);
  buf(\xm8051_golden_model_1.n1299 [141], input_sha_func_48[45]);
  buf(\xm8051_golden_model_1.n1299 [142], input_sha_func_48[46]);
  buf(\xm8051_golden_model_1.n1299 [143], input_sha_func_48[47]);
  buf(\xm8051_golden_model_1.n1299 [144], input_sha_func_48[48]);
  buf(\xm8051_golden_model_1.n1299 [145], input_sha_func_48[49]);
  buf(\xm8051_golden_model_1.n1299 [146], input_sha_func_48[50]);
  buf(\xm8051_golden_model_1.n1299 [147], input_sha_func_48[51]);
  buf(\xm8051_golden_model_1.n1299 [148], input_sha_func_48[52]);
  buf(\xm8051_golden_model_1.n1299 [149], input_sha_func_48[53]);
  buf(\xm8051_golden_model_1.n1299 [150], input_sha_func_48[54]);
  buf(\xm8051_golden_model_1.n1299 [151], input_sha_func_48[55]);
  buf(\xm8051_golden_model_1.n1299 [152], input_sha_func_48[56]);
  buf(\xm8051_golden_model_1.n1299 [153], input_sha_func_48[57]);
  buf(\xm8051_golden_model_1.n1299 [154], input_sha_func_48[58]);
  buf(\xm8051_golden_model_1.n1299 [155], input_sha_func_48[59]);
  buf(\xm8051_golden_model_1.n1299 [156], input_sha_func_48[60]);
  buf(\xm8051_golden_model_1.n1299 [157], input_sha_func_48[61]);
  buf(\xm8051_golden_model_1.n1299 [158], input_sha_func_48[62]);
  buf(\xm8051_golden_model_1.n1299 [159], input_sha_func_48[63]);
  buf(\xm8051_golden_model_1.n0524 [0], \xm8051_golden_model_1.aes_len [8]);
  buf(\xm8051_golden_model_1.n0524 [1], \xm8051_golden_model_1.aes_len [9]);
  buf(\xm8051_golden_model_1.n0524 [2], \xm8051_golden_model_1.aes_len [10]);
  buf(\xm8051_golden_model_1.n0524 [3], \xm8051_golden_model_1.aes_len [11]);
  buf(\xm8051_golden_model_1.n0524 [4], \xm8051_golden_model_1.aes_len [12]);
  buf(\xm8051_golden_model_1.n0524 [5], \xm8051_golden_model_1.aes_len [13]);
  buf(\xm8051_golden_model_1.n0524 [6], \xm8051_golden_model_1.aes_len [14]);
  buf(\xm8051_golden_model_1.n0524 [7], \xm8051_golden_model_1.aes_len [15]);
  buf(\xm8051_golden_model_1.n0523 [0], \xm8051_golden_model_1.aes_len [0]);
  buf(\xm8051_golden_model_1.n0523 [1], \xm8051_golden_model_1.aes_len [1]);
  buf(\xm8051_golden_model_1.n0523 [2], \xm8051_golden_model_1.aes_len [2]);
  buf(\xm8051_golden_model_1.n0523 [3], \xm8051_golden_model_1.aes_len [3]);
  buf(\xm8051_golden_model_1.n0523 [4], \xm8051_golden_model_1.aes_len [4]);
  buf(\xm8051_golden_model_1.n0523 [5], \xm8051_golden_model_1.aes_len [5]);
  buf(\xm8051_golden_model_1.n0523 [6], \xm8051_golden_model_1.aes_len [6]);
  buf(\xm8051_golden_model_1.n0523 [7], \xm8051_golden_model_1.aes_len [7]);
  buf(\xm8051_golden_model_1.n0931 [0], input_sha_func_2[0]);
  buf(\xm8051_golden_model_1.n0931 [1], input_sha_func_2[1]);
  buf(\xm8051_golden_model_1.n0931 [2], input_sha_func_2[2]);
  buf(\xm8051_golden_model_1.n0931 [3], input_sha_func_2[3]);
  buf(\xm8051_golden_model_1.n0931 [4], input_sha_func_2[4]);
  buf(\xm8051_golden_model_1.n0931 [5], input_sha_func_2[5]);
  buf(\xm8051_golden_model_1.n0931 [6], input_sha_func_2[6]);
  buf(\xm8051_golden_model_1.n0931 [7], input_sha_func_2[7]);
  buf(\xm8051_golden_model_1.n0931 [8], input_sha_func_2[8]);
  buf(\xm8051_golden_model_1.n0931 [9], input_sha_func_2[9]);
  buf(\xm8051_golden_model_1.n0931 [10], input_sha_func_2[10]);
  buf(\xm8051_golden_model_1.n0931 [11], input_sha_func_2[11]);
  buf(\xm8051_golden_model_1.n0931 [12], input_sha_func_2[12]);
  buf(\xm8051_golden_model_1.n0931 [13], input_sha_func_2[13]);
  buf(\xm8051_golden_model_1.n0931 [14], input_sha_func_2[14]);
  buf(\xm8051_golden_model_1.n0931 [15], input_sha_func_2[15]);
  buf(\xm8051_golden_model_1.n0931 [16], input_sha_func_2[16]);
  buf(\xm8051_golden_model_1.n0931 [17], input_sha_func_2[17]);
  buf(\xm8051_golden_model_1.n0931 [18], input_sha_func_2[18]);
  buf(\xm8051_golden_model_1.n0931 [19], input_sha_func_2[19]);
  buf(\xm8051_golden_model_1.n0931 [20], input_sha_func_2[20]);
  buf(\xm8051_golden_model_1.n0931 [21], input_sha_func_2[21]);
  buf(\xm8051_golden_model_1.n0931 [22], input_sha_func_2[22]);
  buf(\xm8051_golden_model_1.n0931 [23], input_sha_func_2[23]);
  buf(\xm8051_golden_model_1.n0931 [24], input_sha_func_2[24]);
  buf(\xm8051_golden_model_1.n0931 [25], input_sha_func_2[25]);
  buf(\xm8051_golden_model_1.n0931 [26], input_sha_func_2[26]);
  buf(\xm8051_golden_model_1.n0931 [27], input_sha_func_2[27]);
  buf(\xm8051_golden_model_1.n0931 [28], input_sha_func_2[28]);
  buf(\xm8051_golden_model_1.n0931 [29], input_sha_func_2[29]);
  buf(\xm8051_golden_model_1.n0931 [30], input_sha_func_2[30]);
  buf(\xm8051_golden_model_1.n0931 [31], input_sha_func_2[31]);
  buf(\xm8051_golden_model_1.n0931 [32], input_sha_func_1[0]);
  buf(\xm8051_golden_model_1.n0931 [33], input_sha_func_1[1]);
  buf(\xm8051_golden_model_1.n0931 [34], input_sha_func_1[2]);
  buf(\xm8051_golden_model_1.n0931 [35], input_sha_func_1[3]);
  buf(\xm8051_golden_model_1.n0931 [36], input_sha_func_1[4]);
  buf(\xm8051_golden_model_1.n0931 [37], input_sha_func_1[5]);
  buf(\xm8051_golden_model_1.n0931 [38], input_sha_func_1[6]);
  buf(\xm8051_golden_model_1.n0931 [39], input_sha_func_1[7]);
  buf(\xm8051_golden_model_1.n0931 [40], input_sha_func_1[8]);
  buf(\xm8051_golden_model_1.n0931 [41], input_sha_func_1[9]);
  buf(\xm8051_golden_model_1.n0931 [42], input_sha_func_1[10]);
  buf(\xm8051_golden_model_1.n0931 [43], input_sha_func_1[11]);
  buf(\xm8051_golden_model_1.n0931 [44], input_sha_func_1[12]);
  buf(\xm8051_golden_model_1.n0931 [45], input_sha_func_1[13]);
  buf(\xm8051_golden_model_1.n0931 [46], input_sha_func_1[14]);
  buf(\xm8051_golden_model_1.n0931 [47], input_sha_func_1[15]);
  buf(\xm8051_golden_model_1.n0931 [48], input_sha_func_1[16]);
  buf(\xm8051_golden_model_1.n0931 [49], input_sha_func_1[17]);
  buf(\xm8051_golden_model_1.n0931 [50], input_sha_func_1[18]);
  buf(\xm8051_golden_model_1.n0931 [51], input_sha_func_1[19]);
  buf(\xm8051_golden_model_1.n0931 [52], input_sha_func_1[20]);
  buf(\xm8051_golden_model_1.n0931 [53], input_sha_func_1[21]);
  buf(\xm8051_golden_model_1.n0931 [54], input_sha_func_1[22]);
  buf(\xm8051_golden_model_1.n0931 [55], input_sha_func_1[23]);
  buf(\xm8051_golden_model_1.n0931 [56], input_sha_func_1[24]);
  buf(\xm8051_golden_model_1.n0931 [57], input_sha_func_1[25]);
  buf(\xm8051_golden_model_1.n0931 [58], input_sha_func_1[26]);
  buf(\xm8051_golden_model_1.n0931 [59], input_sha_func_1[27]);
  buf(\xm8051_golden_model_1.n0931 [60], input_sha_func_1[28]);
  buf(\xm8051_golden_model_1.n0931 [61], input_sha_func_1[29]);
  buf(\xm8051_golden_model_1.n0931 [62], input_sha_func_1[30]);
  buf(\xm8051_golden_model_1.n0931 [63], input_sha_func_1[31]);
  buf(\xm8051_golden_model_1.n0931 [64], input_sha_func_1[32]);
  buf(\xm8051_golden_model_1.n0931 [65], input_sha_func_1[33]);
  buf(\xm8051_golden_model_1.n0931 [66], input_sha_func_1[34]);
  buf(\xm8051_golden_model_1.n0931 [67], input_sha_func_1[35]);
  buf(\xm8051_golden_model_1.n0931 [68], input_sha_func_1[36]);
  buf(\xm8051_golden_model_1.n0931 [69], input_sha_func_1[37]);
  buf(\xm8051_golden_model_1.n0931 [70], input_sha_func_1[38]);
  buf(\xm8051_golden_model_1.n0931 [71], input_sha_func_1[39]);
  buf(\xm8051_golden_model_1.n0931 [72], input_sha_func_1[40]);
  buf(\xm8051_golden_model_1.n0931 [73], input_sha_func_1[41]);
  buf(\xm8051_golden_model_1.n0931 [74], input_sha_func_1[42]);
  buf(\xm8051_golden_model_1.n0931 [75], input_sha_func_1[43]);
  buf(\xm8051_golden_model_1.n0931 [76], input_sha_func_1[44]);
  buf(\xm8051_golden_model_1.n0931 [77], input_sha_func_1[45]);
  buf(\xm8051_golden_model_1.n0931 [78], input_sha_func_1[46]);
  buf(\xm8051_golden_model_1.n0931 [79], input_sha_func_1[47]);
  buf(\xm8051_golden_model_1.n0931 [80], input_sha_func_1[48]);
  buf(\xm8051_golden_model_1.n0931 [81], input_sha_func_1[49]);
  buf(\xm8051_golden_model_1.n0931 [82], input_sha_func_1[50]);
  buf(\xm8051_golden_model_1.n0931 [83], input_sha_func_1[51]);
  buf(\xm8051_golden_model_1.n0931 [84], input_sha_func_1[52]);
  buf(\xm8051_golden_model_1.n0931 [85], input_sha_func_1[53]);
  buf(\xm8051_golden_model_1.n0931 [86], input_sha_func_1[54]);
  buf(\xm8051_golden_model_1.n0931 [87], input_sha_func_1[55]);
  buf(\xm8051_golden_model_1.n0931 [88], input_sha_func_1[56]);
  buf(\xm8051_golden_model_1.n0931 [89], input_sha_func_1[57]);
  buf(\xm8051_golden_model_1.n0931 [90], input_sha_func_1[58]);
  buf(\xm8051_golden_model_1.n0931 [91], input_sha_func_1[59]);
  buf(\xm8051_golden_model_1.n0931 [92], input_sha_func_1[60]);
  buf(\xm8051_golden_model_1.n0931 [93], input_sha_func_1[61]);
  buf(\xm8051_golden_model_1.n0931 [94], input_sha_func_1[62]);
  buf(\xm8051_golden_model_1.n0931 [95], input_sha_func_1[63]);
  buf(\xm8051_golden_model_1.n0931 [96], input_sha_func_0[0]);
  buf(\xm8051_golden_model_1.n0931 [97], input_sha_func_0[1]);
  buf(\xm8051_golden_model_1.n0931 [98], input_sha_func_0[2]);
  buf(\xm8051_golden_model_1.n0931 [99], input_sha_func_0[3]);
  buf(\xm8051_golden_model_1.n0931 [100], input_sha_func_0[4]);
  buf(\xm8051_golden_model_1.n0931 [101], input_sha_func_0[5]);
  buf(\xm8051_golden_model_1.n0931 [102], input_sha_func_0[6]);
  buf(\xm8051_golden_model_1.n0931 [103], input_sha_func_0[7]);
  buf(\xm8051_golden_model_1.n0931 [104], input_sha_func_0[8]);
  buf(\xm8051_golden_model_1.n0931 [105], input_sha_func_0[9]);
  buf(\xm8051_golden_model_1.n0931 [106], input_sha_func_0[10]);
  buf(\xm8051_golden_model_1.n0931 [107], input_sha_func_0[11]);
  buf(\xm8051_golden_model_1.n0931 [108], input_sha_func_0[12]);
  buf(\xm8051_golden_model_1.n0931 [109], input_sha_func_0[13]);
  buf(\xm8051_golden_model_1.n0931 [110], input_sha_func_0[14]);
  buf(\xm8051_golden_model_1.n0931 [111], input_sha_func_0[15]);
  buf(\xm8051_golden_model_1.n0931 [112], input_sha_func_0[16]);
  buf(\xm8051_golden_model_1.n0931 [113], input_sha_func_0[17]);
  buf(\xm8051_golden_model_1.n0931 [114], input_sha_func_0[18]);
  buf(\xm8051_golden_model_1.n0931 [115], input_sha_func_0[19]);
  buf(\xm8051_golden_model_1.n0931 [116], input_sha_func_0[20]);
  buf(\xm8051_golden_model_1.n0931 [117], input_sha_func_0[21]);
  buf(\xm8051_golden_model_1.n0931 [118], input_sha_func_0[22]);
  buf(\xm8051_golden_model_1.n0931 [119], input_sha_func_0[23]);
  buf(\xm8051_golden_model_1.n0931 [120], input_sha_func_0[24]);
  buf(\xm8051_golden_model_1.n0931 [121], input_sha_func_0[25]);
  buf(\xm8051_golden_model_1.n0931 [122], input_sha_func_0[26]);
  buf(\xm8051_golden_model_1.n0931 [123], input_sha_func_0[27]);
  buf(\xm8051_golden_model_1.n0931 [124], input_sha_func_0[28]);
  buf(\xm8051_golden_model_1.n0931 [125], input_sha_func_0[29]);
  buf(\xm8051_golden_model_1.n0931 [126], input_sha_func_0[30]);
  buf(\xm8051_golden_model_1.n0931 [127], input_sha_func_0[31]);
  buf(\xm8051_golden_model_1.n0931 [128], input_sha_func_0[32]);
  buf(\xm8051_golden_model_1.n0931 [129], input_sha_func_0[33]);
  buf(\xm8051_golden_model_1.n0931 [130], input_sha_func_0[34]);
  buf(\xm8051_golden_model_1.n0931 [131], input_sha_func_0[35]);
  buf(\xm8051_golden_model_1.n0931 [132], input_sha_func_0[36]);
  buf(\xm8051_golden_model_1.n0931 [133], input_sha_func_0[37]);
  buf(\xm8051_golden_model_1.n0931 [134], input_sha_func_0[38]);
  buf(\xm8051_golden_model_1.n0931 [135], input_sha_func_0[39]);
  buf(\xm8051_golden_model_1.n0931 [136], input_sha_func_0[40]);
  buf(\xm8051_golden_model_1.n0931 [137], input_sha_func_0[41]);
  buf(\xm8051_golden_model_1.n0931 [138], input_sha_func_0[42]);
  buf(\xm8051_golden_model_1.n0931 [139], input_sha_func_0[43]);
  buf(\xm8051_golden_model_1.n0931 [140], input_sha_func_0[44]);
  buf(\xm8051_golden_model_1.n0931 [141], input_sha_func_0[45]);
  buf(\xm8051_golden_model_1.n0931 [142], input_sha_func_0[46]);
  buf(\xm8051_golden_model_1.n0931 [143], input_sha_func_0[47]);
  buf(\xm8051_golden_model_1.n0931 [144], input_sha_func_0[48]);
  buf(\xm8051_golden_model_1.n0931 [145], input_sha_func_0[49]);
  buf(\xm8051_golden_model_1.n0931 [146], input_sha_func_0[50]);
  buf(\xm8051_golden_model_1.n0931 [147], input_sha_func_0[51]);
  buf(\xm8051_golden_model_1.n0931 [148], input_sha_func_0[52]);
  buf(\xm8051_golden_model_1.n0931 [149], input_sha_func_0[53]);
  buf(\xm8051_golden_model_1.n0931 [150], input_sha_func_0[54]);
  buf(\xm8051_golden_model_1.n0931 [151], input_sha_func_0[55]);
  buf(\xm8051_golden_model_1.n0931 [152], input_sha_func_0[56]);
  buf(\xm8051_golden_model_1.n0931 [153], input_sha_func_0[57]);
  buf(\xm8051_golden_model_1.n0931 [154], input_sha_func_0[58]);
  buf(\xm8051_golden_model_1.n0931 [155], input_sha_func_0[59]);
  buf(\xm8051_golden_model_1.n0931 [156], input_sha_func_0[60]);
  buf(\xm8051_golden_model_1.n0931 [157], input_sha_func_0[61]);
  buf(\xm8051_golden_model_1.n0931 [158], input_sha_func_0[62]);
  buf(\xm8051_golden_model_1.n0931 [159], input_sha_func_0[63]);
  buf(\xm8051_golden_model_1.n0515 , proc_addr[0]);
  buf(\xm8051_golden_model_1.n1295 [0], input_sha_func_47[0]);
  buf(\xm8051_golden_model_1.n1295 [1], input_sha_func_47[1]);
  buf(\xm8051_golden_model_1.n1295 [2], input_sha_func_47[2]);
  buf(\xm8051_golden_model_1.n1295 [3], input_sha_func_47[3]);
  buf(\xm8051_golden_model_1.n1295 [4], input_sha_func_47[4]);
  buf(\xm8051_golden_model_1.n1295 [5], input_sha_func_47[5]);
  buf(\xm8051_golden_model_1.n1295 [6], input_sha_func_47[6]);
  buf(\xm8051_golden_model_1.n1295 [7], input_sha_func_47[7]);
  buf(\xm8051_golden_model_1.n1295 [8], input_sha_func_47[8]);
  buf(\xm8051_golden_model_1.n1295 [9], input_sha_func_47[9]);
  buf(\xm8051_golden_model_1.n1295 [10], input_sha_func_47[10]);
  buf(\xm8051_golden_model_1.n1295 [11], input_sha_func_47[11]);
  buf(\xm8051_golden_model_1.n1295 [12], input_sha_func_47[12]);
  buf(\xm8051_golden_model_1.n1295 [13], input_sha_func_47[13]);
  buf(\xm8051_golden_model_1.n1295 [14], input_sha_func_47[14]);
  buf(\xm8051_golden_model_1.n1295 [15], input_sha_func_47[15]);
  buf(\xm8051_golden_model_1.n1295 [16], input_sha_func_47[16]);
  buf(\xm8051_golden_model_1.n1295 [17], input_sha_func_47[17]);
  buf(\xm8051_golden_model_1.n1295 [18], input_sha_func_47[18]);
  buf(\xm8051_golden_model_1.n1295 [19], input_sha_func_47[19]);
  buf(\xm8051_golden_model_1.n1295 [20], input_sha_func_47[20]);
  buf(\xm8051_golden_model_1.n1295 [21], input_sha_func_47[21]);
  buf(\xm8051_golden_model_1.n1295 [22], input_sha_func_47[22]);
  buf(\xm8051_golden_model_1.n1295 [23], input_sha_func_47[23]);
  buf(\xm8051_golden_model_1.n1295 [24], input_sha_func_47[24]);
  buf(\xm8051_golden_model_1.n1295 [25], input_sha_func_47[25]);
  buf(\xm8051_golden_model_1.n1295 [26], input_sha_func_47[26]);
  buf(\xm8051_golden_model_1.n1295 [27], input_sha_func_47[27]);
  buf(\xm8051_golden_model_1.n1295 [28], input_sha_func_47[28]);
  buf(\xm8051_golden_model_1.n1295 [29], input_sha_func_47[29]);
  buf(\xm8051_golden_model_1.n1295 [30], input_sha_func_47[30]);
  buf(\xm8051_golden_model_1.n1295 [31], input_sha_func_47[31]);
  buf(\xm8051_golden_model_1.n1295 [32], input_sha_func_46[0]);
  buf(\xm8051_golden_model_1.n1295 [33], input_sha_func_46[1]);
  buf(\xm8051_golden_model_1.n1295 [34], input_sha_func_46[2]);
  buf(\xm8051_golden_model_1.n1295 [35], input_sha_func_46[3]);
  buf(\xm8051_golden_model_1.n1295 [36], input_sha_func_46[4]);
  buf(\xm8051_golden_model_1.n1295 [37], input_sha_func_46[5]);
  buf(\xm8051_golden_model_1.n1295 [38], input_sha_func_46[6]);
  buf(\xm8051_golden_model_1.n1295 [39], input_sha_func_46[7]);
  buf(\xm8051_golden_model_1.n1295 [40], input_sha_func_46[8]);
  buf(\xm8051_golden_model_1.n1295 [41], input_sha_func_46[9]);
  buf(\xm8051_golden_model_1.n1295 [42], input_sha_func_46[10]);
  buf(\xm8051_golden_model_1.n1295 [43], input_sha_func_46[11]);
  buf(\xm8051_golden_model_1.n1295 [44], input_sha_func_46[12]);
  buf(\xm8051_golden_model_1.n1295 [45], input_sha_func_46[13]);
  buf(\xm8051_golden_model_1.n1295 [46], input_sha_func_46[14]);
  buf(\xm8051_golden_model_1.n1295 [47], input_sha_func_46[15]);
  buf(\xm8051_golden_model_1.n1295 [48], input_sha_func_46[16]);
  buf(\xm8051_golden_model_1.n1295 [49], input_sha_func_46[17]);
  buf(\xm8051_golden_model_1.n1295 [50], input_sha_func_46[18]);
  buf(\xm8051_golden_model_1.n1295 [51], input_sha_func_46[19]);
  buf(\xm8051_golden_model_1.n1295 [52], input_sha_func_46[20]);
  buf(\xm8051_golden_model_1.n1295 [53], input_sha_func_46[21]);
  buf(\xm8051_golden_model_1.n1295 [54], input_sha_func_46[22]);
  buf(\xm8051_golden_model_1.n1295 [55], input_sha_func_46[23]);
  buf(\xm8051_golden_model_1.n1295 [56], input_sha_func_46[24]);
  buf(\xm8051_golden_model_1.n1295 [57], input_sha_func_46[25]);
  buf(\xm8051_golden_model_1.n1295 [58], input_sha_func_46[26]);
  buf(\xm8051_golden_model_1.n1295 [59], input_sha_func_46[27]);
  buf(\xm8051_golden_model_1.n1295 [60], input_sha_func_46[28]);
  buf(\xm8051_golden_model_1.n1295 [61], input_sha_func_46[29]);
  buf(\xm8051_golden_model_1.n1295 [62], input_sha_func_46[30]);
  buf(\xm8051_golden_model_1.n1295 [63], input_sha_func_46[31]);
  buf(\xm8051_golden_model_1.n1295 [64], input_sha_func_46[32]);
  buf(\xm8051_golden_model_1.n1295 [65], input_sha_func_46[33]);
  buf(\xm8051_golden_model_1.n1295 [66], input_sha_func_46[34]);
  buf(\xm8051_golden_model_1.n1295 [67], input_sha_func_46[35]);
  buf(\xm8051_golden_model_1.n1295 [68], input_sha_func_46[36]);
  buf(\xm8051_golden_model_1.n1295 [69], input_sha_func_46[37]);
  buf(\xm8051_golden_model_1.n1295 [70], input_sha_func_46[38]);
  buf(\xm8051_golden_model_1.n1295 [71], input_sha_func_46[39]);
  buf(\xm8051_golden_model_1.n1295 [72], input_sha_func_46[40]);
  buf(\xm8051_golden_model_1.n1295 [73], input_sha_func_46[41]);
  buf(\xm8051_golden_model_1.n1295 [74], input_sha_func_46[42]);
  buf(\xm8051_golden_model_1.n1295 [75], input_sha_func_46[43]);
  buf(\xm8051_golden_model_1.n1295 [76], input_sha_func_46[44]);
  buf(\xm8051_golden_model_1.n1295 [77], input_sha_func_46[45]);
  buf(\xm8051_golden_model_1.n1295 [78], input_sha_func_46[46]);
  buf(\xm8051_golden_model_1.n1295 [79], input_sha_func_46[47]);
  buf(\xm8051_golden_model_1.n1295 [80], input_sha_func_46[48]);
  buf(\xm8051_golden_model_1.n1295 [81], input_sha_func_46[49]);
  buf(\xm8051_golden_model_1.n1295 [82], input_sha_func_46[50]);
  buf(\xm8051_golden_model_1.n1295 [83], input_sha_func_46[51]);
  buf(\xm8051_golden_model_1.n1295 [84], input_sha_func_46[52]);
  buf(\xm8051_golden_model_1.n1295 [85], input_sha_func_46[53]);
  buf(\xm8051_golden_model_1.n1295 [86], input_sha_func_46[54]);
  buf(\xm8051_golden_model_1.n1295 [87], input_sha_func_46[55]);
  buf(\xm8051_golden_model_1.n1295 [88], input_sha_func_46[56]);
  buf(\xm8051_golden_model_1.n1295 [89], input_sha_func_46[57]);
  buf(\xm8051_golden_model_1.n1295 [90], input_sha_func_46[58]);
  buf(\xm8051_golden_model_1.n1295 [91], input_sha_func_46[59]);
  buf(\xm8051_golden_model_1.n1295 [92], input_sha_func_46[60]);
  buf(\xm8051_golden_model_1.n1295 [93], input_sha_func_46[61]);
  buf(\xm8051_golden_model_1.n1295 [94], input_sha_func_46[62]);
  buf(\xm8051_golden_model_1.n1295 [95], input_sha_func_46[63]);
  buf(\xm8051_golden_model_1.n1295 [96], input_sha_func_45[0]);
  buf(\xm8051_golden_model_1.n1295 [97], input_sha_func_45[1]);
  buf(\xm8051_golden_model_1.n1295 [98], input_sha_func_45[2]);
  buf(\xm8051_golden_model_1.n1295 [99], input_sha_func_45[3]);
  buf(\xm8051_golden_model_1.n1295 [100], input_sha_func_45[4]);
  buf(\xm8051_golden_model_1.n1295 [101], input_sha_func_45[5]);
  buf(\xm8051_golden_model_1.n1295 [102], input_sha_func_45[6]);
  buf(\xm8051_golden_model_1.n1295 [103], input_sha_func_45[7]);
  buf(\xm8051_golden_model_1.n1295 [104], input_sha_func_45[8]);
  buf(\xm8051_golden_model_1.n1295 [105], input_sha_func_45[9]);
  buf(\xm8051_golden_model_1.n1295 [106], input_sha_func_45[10]);
  buf(\xm8051_golden_model_1.n1295 [107], input_sha_func_45[11]);
  buf(\xm8051_golden_model_1.n1295 [108], input_sha_func_45[12]);
  buf(\xm8051_golden_model_1.n1295 [109], input_sha_func_45[13]);
  buf(\xm8051_golden_model_1.n1295 [110], input_sha_func_45[14]);
  buf(\xm8051_golden_model_1.n1295 [111], input_sha_func_45[15]);
  buf(\xm8051_golden_model_1.n1295 [112], input_sha_func_45[16]);
  buf(\xm8051_golden_model_1.n1295 [113], input_sha_func_45[17]);
  buf(\xm8051_golden_model_1.n1295 [114], input_sha_func_45[18]);
  buf(\xm8051_golden_model_1.n1295 [115], input_sha_func_45[19]);
  buf(\xm8051_golden_model_1.n1295 [116], input_sha_func_45[20]);
  buf(\xm8051_golden_model_1.n1295 [117], input_sha_func_45[21]);
  buf(\xm8051_golden_model_1.n1295 [118], input_sha_func_45[22]);
  buf(\xm8051_golden_model_1.n1295 [119], input_sha_func_45[23]);
  buf(\xm8051_golden_model_1.n1295 [120], input_sha_func_45[24]);
  buf(\xm8051_golden_model_1.n1295 [121], input_sha_func_45[25]);
  buf(\xm8051_golden_model_1.n1295 [122], input_sha_func_45[26]);
  buf(\xm8051_golden_model_1.n1295 [123], input_sha_func_45[27]);
  buf(\xm8051_golden_model_1.n1295 [124], input_sha_func_45[28]);
  buf(\xm8051_golden_model_1.n1295 [125], input_sha_func_45[29]);
  buf(\xm8051_golden_model_1.n1295 [126], input_sha_func_45[30]);
  buf(\xm8051_golden_model_1.n1295 [127], input_sha_func_45[31]);
  buf(\xm8051_golden_model_1.n1295 [128], input_sha_func_45[32]);
  buf(\xm8051_golden_model_1.n1295 [129], input_sha_func_45[33]);
  buf(\xm8051_golden_model_1.n1295 [130], input_sha_func_45[34]);
  buf(\xm8051_golden_model_1.n1295 [131], input_sha_func_45[35]);
  buf(\xm8051_golden_model_1.n1295 [132], input_sha_func_45[36]);
  buf(\xm8051_golden_model_1.n1295 [133], input_sha_func_45[37]);
  buf(\xm8051_golden_model_1.n1295 [134], input_sha_func_45[38]);
  buf(\xm8051_golden_model_1.n1295 [135], input_sha_func_45[39]);
  buf(\xm8051_golden_model_1.n1295 [136], input_sha_func_45[40]);
  buf(\xm8051_golden_model_1.n1295 [137], input_sha_func_45[41]);
  buf(\xm8051_golden_model_1.n1295 [138], input_sha_func_45[42]);
  buf(\xm8051_golden_model_1.n1295 [139], input_sha_func_45[43]);
  buf(\xm8051_golden_model_1.n1295 [140], input_sha_func_45[44]);
  buf(\xm8051_golden_model_1.n1295 [141], input_sha_func_45[45]);
  buf(\xm8051_golden_model_1.n1295 [142], input_sha_func_45[46]);
  buf(\xm8051_golden_model_1.n1295 [143], input_sha_func_45[47]);
  buf(\xm8051_golden_model_1.n1295 [144], input_sha_func_45[48]);
  buf(\xm8051_golden_model_1.n1295 [145], input_sha_func_45[49]);
  buf(\xm8051_golden_model_1.n1295 [146], input_sha_func_45[50]);
  buf(\xm8051_golden_model_1.n1295 [147], input_sha_func_45[51]);
  buf(\xm8051_golden_model_1.n1295 [148], input_sha_func_45[52]);
  buf(\xm8051_golden_model_1.n1295 [149], input_sha_func_45[53]);
  buf(\xm8051_golden_model_1.n1295 [150], input_sha_func_45[54]);
  buf(\xm8051_golden_model_1.n1295 [151], input_sha_func_45[55]);
  buf(\xm8051_golden_model_1.n1295 [152], input_sha_func_45[56]);
  buf(\xm8051_golden_model_1.n1295 [153], input_sha_func_45[57]);
  buf(\xm8051_golden_model_1.n1295 [154], input_sha_func_45[58]);
  buf(\xm8051_golden_model_1.n1295 [155], input_sha_func_45[59]);
  buf(\xm8051_golden_model_1.n1295 [156], input_sha_func_45[60]);
  buf(\xm8051_golden_model_1.n1295 [157], input_sha_func_45[61]);
  buf(\xm8051_golden_model_1.n1295 [158], input_sha_func_45[62]);
  buf(\xm8051_golden_model_1.n1295 [159], input_sha_func_45[63]);
  buf(\xm8051_golden_model_1.n0512 [0], 1'b0);
  buf(\xm8051_golden_model_1.n0512 [1], proc_addr[1]);
  buf(\xm8051_golden_model_1.n0512 [2], proc_addr[2]);
  buf(\xm8051_golden_model_1.n0512 [3], proc_addr[3]);
  buf(\xm8051_golden_model_1.n0512 [4], proc_addr[4]);
  buf(\xm8051_golden_model_1.n0512 [5], proc_addr[5]);
  buf(\xm8051_golden_model_1.n0512 [6], proc_addr[6]);
  buf(\xm8051_golden_model_1.n0512 [7], proc_addr[7]);
  buf(\xm8051_golden_model_1.n0512 [8], proc_addr[8]);
  buf(\xm8051_golden_model_1.n0512 [9], proc_addr[9]);
  buf(\xm8051_golden_model_1.n0512 [10], proc_addr[10]);
  buf(\xm8051_golden_model_1.n0512 [11], proc_addr[11]);
  buf(\xm8051_golden_model_1.n0512 [12], proc_addr[12]);
  buf(\xm8051_golden_model_1.n0512 [13], proc_addr[13]);
  buf(\xm8051_golden_model_1.n0512 [14], proc_addr[14]);
  buf(\xm8051_golden_model_1.n0512 [15], proc_addr[15]);
  buf(\xm8051_golden_model_1.n0510 [0], proc_addr[1]);
  buf(\xm8051_golden_model_1.n0510 [1], proc_addr[2]);
  buf(\xm8051_golden_model_1.n0510 [2], proc_addr[3]);
  buf(\xm8051_golden_model_1.n0510 [3], proc_addr[4]);
  buf(\xm8051_golden_model_1.n0510 [4], proc_addr[5]);
  buf(\xm8051_golden_model_1.n0510 [5], proc_addr[6]);
  buf(\xm8051_golden_model_1.n0510 [6], proc_addr[7]);
  buf(\xm8051_golden_model_1.n0510 [7], proc_addr[8]);
  buf(\xm8051_golden_model_1.n0510 [8], proc_addr[9]);
  buf(\xm8051_golden_model_1.n0510 [9], proc_addr[10]);
  buf(\xm8051_golden_model_1.n0510 [10], proc_addr[11]);
  buf(\xm8051_golden_model_1.n0510 [11], proc_addr[12]);
  buf(\xm8051_golden_model_1.n0510 [12], proc_addr[13]);
  buf(\xm8051_golden_model_1.n0510 [13], proc_addr[14]);
  buf(\xm8051_golden_model_1.n0510 [14], proc_addr[15]);
  buf(\xm8051_golden_model_1.n1290 [0], RD_xram_15[0]);
  buf(\xm8051_golden_model_1.n1290 [1], RD_xram_15[1]);
  buf(\xm8051_golden_model_1.n1290 [2], RD_xram_15[2]);
  buf(\xm8051_golden_model_1.n1290 [3], RD_xram_15[3]);
  buf(\xm8051_golden_model_1.n1290 [4], RD_xram_15[4]);
  buf(\xm8051_golden_model_1.n1290 [5], RD_xram_15[5]);
  buf(\xm8051_golden_model_1.n1290 [6], RD_xram_15[6]);
  buf(\xm8051_golden_model_1.n1290 [7], RD_xram_15[7]);
  buf(\xm8051_golden_model_1.n1290 [8], RD_xram_14[0]);
  buf(\xm8051_golden_model_1.n1290 [9], RD_xram_14[1]);
  buf(\xm8051_golden_model_1.n1290 [10], RD_xram_14[2]);
  buf(\xm8051_golden_model_1.n1290 [11], RD_xram_14[3]);
  buf(\xm8051_golden_model_1.n1290 [12], RD_xram_14[4]);
  buf(\xm8051_golden_model_1.n1290 [13], RD_xram_14[5]);
  buf(\xm8051_golden_model_1.n1290 [14], RD_xram_14[6]);
  buf(\xm8051_golden_model_1.n1290 [15], RD_xram_14[7]);
  buf(\xm8051_golden_model_1.n1290 [16], RD_xram_13[0]);
  buf(\xm8051_golden_model_1.n1290 [17], RD_xram_13[1]);
  buf(\xm8051_golden_model_1.n1290 [18], RD_xram_13[2]);
  buf(\xm8051_golden_model_1.n1290 [19], RD_xram_13[3]);
  buf(\xm8051_golden_model_1.n1290 [20], RD_xram_13[4]);
  buf(\xm8051_golden_model_1.n1290 [21], RD_xram_13[5]);
  buf(\xm8051_golden_model_1.n1290 [22], RD_xram_13[6]);
  buf(\xm8051_golden_model_1.n1290 [23], RD_xram_13[7]);
  buf(\xm8051_golden_model_1.n1290 [24], RD_xram_12[0]);
  buf(\xm8051_golden_model_1.n1290 [25], RD_xram_12[1]);
  buf(\xm8051_golden_model_1.n1290 [26], RD_xram_12[2]);
  buf(\xm8051_golden_model_1.n1290 [27], RD_xram_12[3]);
  buf(\xm8051_golden_model_1.n1290 [28], RD_xram_12[4]);
  buf(\xm8051_golden_model_1.n1290 [29], RD_xram_12[5]);
  buf(\xm8051_golden_model_1.n1290 [30], RD_xram_12[6]);
  buf(\xm8051_golden_model_1.n1290 [31], RD_xram_12[7]);
  buf(\xm8051_golden_model_1.n1290 [32], RD_xram_11[0]);
  buf(\xm8051_golden_model_1.n1290 [33], RD_xram_11[1]);
  buf(\xm8051_golden_model_1.n1290 [34], RD_xram_11[2]);
  buf(\xm8051_golden_model_1.n1290 [35], RD_xram_11[3]);
  buf(\xm8051_golden_model_1.n1290 [36], RD_xram_11[4]);
  buf(\xm8051_golden_model_1.n1290 [37], RD_xram_11[5]);
  buf(\xm8051_golden_model_1.n1290 [38], RD_xram_11[6]);
  buf(\xm8051_golden_model_1.n1290 [39], RD_xram_11[7]);
  buf(\xm8051_golden_model_1.n1290 [40], RD_xram_10[0]);
  buf(\xm8051_golden_model_1.n1290 [41], RD_xram_10[1]);
  buf(\xm8051_golden_model_1.n1290 [42], RD_xram_10[2]);
  buf(\xm8051_golden_model_1.n1290 [43], RD_xram_10[3]);
  buf(\xm8051_golden_model_1.n1290 [44], RD_xram_10[4]);
  buf(\xm8051_golden_model_1.n1290 [45], RD_xram_10[5]);
  buf(\xm8051_golden_model_1.n1290 [46], RD_xram_10[6]);
  buf(\xm8051_golden_model_1.n1290 [47], RD_xram_10[7]);
  buf(\xm8051_golden_model_1.n1290 [48], RD_xram_9[0]);
  buf(\xm8051_golden_model_1.n1290 [49], RD_xram_9[1]);
  buf(\xm8051_golden_model_1.n1290 [50], RD_xram_9[2]);
  buf(\xm8051_golden_model_1.n1290 [51], RD_xram_9[3]);
  buf(\xm8051_golden_model_1.n1290 [52], RD_xram_9[4]);
  buf(\xm8051_golden_model_1.n1290 [53], RD_xram_9[5]);
  buf(\xm8051_golden_model_1.n1290 [54], RD_xram_9[6]);
  buf(\xm8051_golden_model_1.n1290 [55], RD_xram_9[7]);
  buf(\xm8051_golden_model_1.n1290 [56], RD_xram_8[0]);
  buf(\xm8051_golden_model_1.n1290 [57], RD_xram_8[1]);
  buf(\xm8051_golden_model_1.n1290 [58], RD_xram_8[2]);
  buf(\xm8051_golden_model_1.n1290 [59], RD_xram_8[3]);
  buf(\xm8051_golden_model_1.n1290 [60], RD_xram_8[4]);
  buf(\xm8051_golden_model_1.n1290 [61], RD_xram_8[5]);
  buf(\xm8051_golden_model_1.n1290 [62], RD_xram_8[6]);
  buf(\xm8051_golden_model_1.n1290 [63], RD_xram_8[7]);
  buf(\xm8051_golden_model_1.n1290 [64], RD_xram_7[0]);
  buf(\xm8051_golden_model_1.n1290 [65], RD_xram_7[1]);
  buf(\xm8051_golden_model_1.n1290 [66], RD_xram_7[2]);
  buf(\xm8051_golden_model_1.n1290 [67], RD_xram_7[3]);
  buf(\xm8051_golden_model_1.n1290 [68], RD_xram_7[4]);
  buf(\xm8051_golden_model_1.n1290 [69], RD_xram_7[5]);
  buf(\xm8051_golden_model_1.n1290 [70], RD_xram_7[6]);
  buf(\xm8051_golden_model_1.n1290 [71], RD_xram_7[7]);
  buf(\xm8051_golden_model_1.n1290 [72], RD_xram_6[0]);
  buf(\xm8051_golden_model_1.n1290 [73], RD_xram_6[1]);
  buf(\xm8051_golden_model_1.n1290 [74], RD_xram_6[2]);
  buf(\xm8051_golden_model_1.n1290 [75], RD_xram_6[3]);
  buf(\xm8051_golden_model_1.n1290 [76], RD_xram_6[4]);
  buf(\xm8051_golden_model_1.n1290 [77], RD_xram_6[5]);
  buf(\xm8051_golden_model_1.n1290 [78], RD_xram_6[6]);
  buf(\xm8051_golden_model_1.n1290 [79], RD_xram_6[7]);
  buf(\xm8051_golden_model_1.n1290 [80], RD_xram_5[0]);
  buf(\xm8051_golden_model_1.n1290 [81], RD_xram_5[1]);
  buf(\xm8051_golden_model_1.n1290 [82], RD_xram_5[2]);
  buf(\xm8051_golden_model_1.n1290 [83], RD_xram_5[3]);
  buf(\xm8051_golden_model_1.n1290 [84], RD_xram_5[4]);
  buf(\xm8051_golden_model_1.n1290 [85], RD_xram_5[5]);
  buf(\xm8051_golden_model_1.n1290 [86], RD_xram_5[6]);
  buf(\xm8051_golden_model_1.n1290 [87], RD_xram_5[7]);
  buf(\xm8051_golden_model_1.n1290 [88], RD_xram_4[0]);
  buf(\xm8051_golden_model_1.n1290 [89], RD_xram_4[1]);
  buf(\xm8051_golden_model_1.n1290 [90], RD_xram_4[2]);
  buf(\xm8051_golden_model_1.n1290 [91], RD_xram_4[3]);
  buf(\xm8051_golden_model_1.n1290 [92], RD_xram_4[4]);
  buf(\xm8051_golden_model_1.n1290 [93], RD_xram_4[5]);
  buf(\xm8051_golden_model_1.n1290 [94], RD_xram_4[6]);
  buf(\xm8051_golden_model_1.n1290 [95], RD_xram_4[7]);
  buf(\xm8051_golden_model_1.n1290 [96], RD_xram_3[0]);
  buf(\xm8051_golden_model_1.n1290 [97], RD_xram_3[1]);
  buf(\xm8051_golden_model_1.n1290 [98], RD_xram_3[2]);
  buf(\xm8051_golden_model_1.n1290 [99], RD_xram_3[3]);
  buf(\xm8051_golden_model_1.n1290 [100], RD_xram_3[4]);
  buf(\xm8051_golden_model_1.n1290 [101], RD_xram_3[5]);
  buf(\xm8051_golden_model_1.n1290 [102], RD_xram_3[6]);
  buf(\xm8051_golden_model_1.n1290 [103], RD_xram_3[7]);
  buf(\xm8051_golden_model_1.n1290 [104], RD_xram_2[0]);
  buf(\xm8051_golden_model_1.n1290 [105], RD_xram_2[1]);
  buf(\xm8051_golden_model_1.n1290 [106], RD_xram_2[2]);
  buf(\xm8051_golden_model_1.n1290 [107], RD_xram_2[3]);
  buf(\xm8051_golden_model_1.n1290 [108], RD_xram_2[4]);
  buf(\xm8051_golden_model_1.n1290 [109], RD_xram_2[5]);
  buf(\xm8051_golden_model_1.n1290 [110], RD_xram_2[6]);
  buf(\xm8051_golden_model_1.n1290 [111], RD_xram_2[7]);
  buf(\xm8051_golden_model_1.n1290 [112], RD_xram_1[0]);
  buf(\xm8051_golden_model_1.n1290 [113], RD_xram_1[1]);
  buf(\xm8051_golden_model_1.n1290 [114], RD_xram_1[2]);
  buf(\xm8051_golden_model_1.n1290 [115], RD_xram_1[3]);
  buf(\xm8051_golden_model_1.n1290 [116], RD_xram_1[4]);
  buf(\xm8051_golden_model_1.n1290 [117], RD_xram_1[5]);
  buf(\xm8051_golden_model_1.n1290 [118], RD_xram_1[6]);
  buf(\xm8051_golden_model_1.n1290 [119], RD_xram_1[7]);
  buf(\xm8051_golden_model_1.n1290 [120], RD_xram_0[0]);
  buf(\xm8051_golden_model_1.n1290 [121], RD_xram_0[1]);
  buf(\xm8051_golden_model_1.n1290 [122], RD_xram_0[2]);
  buf(\xm8051_golden_model_1.n1290 [123], RD_xram_0[3]);
  buf(\xm8051_golden_model_1.n1290 [124], RD_xram_0[4]);
  buf(\xm8051_golden_model_1.n1290 [125], RD_xram_0[5]);
  buf(\xm8051_golden_model_1.n1290 [126], RD_xram_0[6]);
  buf(\xm8051_golden_model_1.n1290 [127], RD_xram_0[7]);
  buf(\xm8051_golden_model_1.n0921 [0], sha_wraddr_gm[0]);
  buf(\xm8051_golden_model_1.n0921 [1], sha_wraddr_gm[1]);
  buf(\xm8051_golden_model_1.n0921 [2], sha_wraddr_gm[2]);
  buf(\xm8051_golden_model_1.n0921 [3], sha_wraddr_gm[3]);
  buf(\xm8051_golden_model_1.n0921 [4], sha_wraddr_gm[4]);
  buf(\xm8051_golden_model_1.n0921 [5], sha_wraddr_gm[5]);
  buf(\xm8051_golden_model_1.n0921 [6], sha_wraddr_gm[6]);
  buf(\xm8051_golden_model_1.n0921 [7], sha_wraddr_gm[7]);
  buf(\xm8051_golden_model_1.n0921 [8], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0921 [9], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0921 [10], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0921 [11], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0921 [12], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0921 [13], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0921 [14], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0921 [15], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0003 [0], \xm8051_golden_model_1.aes_state [0]);
  buf(\xm8051_golden_model_1.n0003 [1], \xm8051_golden_model_1.aes_state [1]);
  buf(\xm8051_golden_model_1.n0003 [2], \xm8051_golden_model_1.sha_state [0]);
  buf(\xm8051_golden_model_1.n0003 [3], \xm8051_golden_model_1.sha_state [1]);
  buf(\xm8051_golden_model_1.n0002 [0], \xm8051_golden_model_1.aes_state [0]);
  buf(\xm8051_golden_model_1.n0002 [1], \xm8051_golden_model_1.aes_state [1]);
  buf(\xm8051_golden_model_1.n0001 [0], \xm8051_golden_model_1.sha_state [0]);
  buf(\xm8051_golden_model_1.n0001 [1], \xm8051_golden_model_1.sha_state [1]);
  buf(\xm8051_golden_model_1.n0920 [0], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0920 [1], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0920 [2], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0920 [3], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0920 [4], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0920 [5], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0920 [6], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0920 [7], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0920 [8], sha_wraddr_gm[8]);
  buf(\xm8051_golden_model_1.n0920 [9], sha_wraddr_gm[9]);
  buf(\xm8051_golden_model_1.n0920 [10], sha_wraddr_gm[10]);
  buf(\xm8051_golden_model_1.n0920 [11], sha_wraddr_gm[11]);
  buf(\xm8051_golden_model_1.n0920 [12], sha_wraddr_gm[12]);
  buf(\xm8051_golden_model_1.n0920 [13], sha_wraddr_gm[13]);
  buf(\xm8051_golden_model_1.n0920 [14], sha_wraddr_gm[14]);
  buf(\xm8051_golden_model_1.n0920 [15], sha_wraddr_gm[15]);
  buf(\xm8051_golden_model_1.n0493 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0493 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0493 [2], \xm8051_golden_model_1.sha_bytes_processed [2]);
  buf(\xm8051_golden_model_1.n0493 [3], \xm8051_golden_model_1.sha_bytes_processed [3]);
  buf(\xm8051_golden_model_1.n0493 [4], \xm8051_golden_model_1.sha_bytes_processed [4]);
  buf(\xm8051_golden_model_1.n0493 [5], \xm8051_golden_model_1.sha_bytes_processed [5]);
  buf(\xm8051_golden_model_1.n0493 [6], \xm8051_golden_model_1.sha_bytes_processed [6]);
  buf(\xm8051_golden_model_1.n0493 [7], \xm8051_golden_model_1.sha_bytes_processed [7]);
  buf(\xm8051_golden_model_1.n0493 [8], \xm8051_golden_model_1.sha_bytes_processed [8]);
  buf(\xm8051_golden_model_1.n0493 [9], \xm8051_golden_model_1.sha_bytes_processed [9]);
  buf(\xm8051_golden_model_1.n0493 [10], \xm8051_golden_model_1.sha_bytes_processed [10]);
  buf(\xm8051_golden_model_1.n0493 [11], \xm8051_golden_model_1.sha_bytes_processed [11]);
  buf(\xm8051_golden_model_1.n0493 [12], \xm8051_golden_model_1.sha_bytes_processed [12]);
  buf(\xm8051_golden_model_1.n0493 [13], \xm8051_golden_model_1.sha_bytes_processed [13]);
  buf(\xm8051_golden_model_1.n0493 [14], \xm8051_golden_model_1.sha_bytes_processed [14]);
  buf(\xm8051_golden_model_1.n0493 [15], \xm8051_golden_model_1.sha_bytes_processed [15]);
  buf(\xm8051_golden_model_1.n0910 [0], \xm8051_golden_model_1.aes_len [0]);
  buf(\xm8051_golden_model_1.n0910 [1], \xm8051_golden_model_1.aes_len [1]);
  buf(\xm8051_golden_model_1.n0910 [2], \xm8051_golden_model_1.aes_len [2]);
  buf(\xm8051_golden_model_1.n0910 [3], \xm8051_golden_model_1.aes_len [3]);
  buf(\xm8051_golden_model_1.n0910 [4], \xm8051_golden_model_1.aes_len [4]);
  buf(\xm8051_golden_model_1.n0910 [5], \xm8051_golden_model_1.aes_len [5]);
  buf(\xm8051_golden_model_1.n0910 [6], \xm8051_golden_model_1.aes_len [6]);
  buf(\xm8051_golden_model_1.n0910 [7], \xm8051_golden_model_1.aes_len [7]);
  buf(\xm8051_golden_model_1.n0910 [8], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0910 [9], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0910 [10], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0910 [11], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0910 [12], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0910 [13], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0910 [14], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0910 [15], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0909 [0], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0909 [1], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0909 [2], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0909 [3], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0909 [4], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0909 [5], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0909 [6], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0909 [7], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0909 [8], \xm8051_golden_model_1.aes_len [8]);
  buf(\xm8051_golden_model_1.n0909 [9], \xm8051_golden_model_1.aes_len [9]);
  buf(\xm8051_golden_model_1.n0909 [10], \xm8051_golden_model_1.aes_len [10]);
  buf(\xm8051_golden_model_1.n0909 [11], \xm8051_golden_model_1.aes_len [11]);
  buf(\xm8051_golden_model_1.n0909 [12], \xm8051_golden_model_1.aes_len [12]);
  buf(\xm8051_golden_model_1.n0909 [13], \xm8051_golden_model_1.aes_len [13]);
  buf(\xm8051_golden_model_1.n0909 [14], \xm8051_golden_model_1.aes_len [14]);
  buf(\xm8051_golden_model_1.n0909 [15], \xm8051_golden_model_1.aes_len [15]);
  buf(\xm8051_golden_model_1.n0483 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0904 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0904 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0904 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0904 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0904 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0904 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0904 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0904 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0903 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0903 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0903 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0903 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0903 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0903 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0903 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0903 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0903 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0903 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0903 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0903 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0903 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0903 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0903 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0903 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\oc8051_xiommu_impl_1.oc8051_xram_i.rst , rst);
  buf(\oc8051_xiommu_impl_1.oc8051_xram_i.clk , clk);
  buf(\xm8051_golden_model_1.n0902 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0902 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0902 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0902 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0902 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0902 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0902 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0902 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0902 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0902 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0902 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0902 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0902 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0902 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0902 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0902 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0902 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0902 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0902 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0902 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0902 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0902 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0902 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0902 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0901 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0901 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0901 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0901 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0901 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0901 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0901 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0901 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0901 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0901 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0901 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0901 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0901 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0901 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0901 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0901 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0901 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0901 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0901 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0901 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0901 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0901 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0901 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0901 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0901 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0901 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0901 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0901 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0901 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0901 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0901 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0901 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0900 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0900 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0900 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0900 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0900 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0900 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0900 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0900 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0900 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0900 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0900 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0900 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0900 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0900 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0900 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0900 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0900 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0900 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0900 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0900 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0900 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0900 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0900 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0900 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0900 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0900 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0900 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0900 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0900 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0900 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0900 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0900 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0900 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0900 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0900 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0900 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0900 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0900 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0900 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0900 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0899 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0899 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0899 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0899 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0899 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0899 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0899 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0899 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0899 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0899 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0899 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0899 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0899 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0899 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0899 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0899 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0899 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0899 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0899 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0899 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0899 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0899 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0899 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0899 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0899 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0899 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0899 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0899 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0899 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0899 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0899 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0899 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0899 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0899 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0899 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0899 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0899 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0899 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0899 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0899 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0899 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0899 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0899 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0899 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0899 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0899 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0899 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0899 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0898 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0898 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0898 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0898 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0898 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0898 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0898 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0898 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0898 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0898 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0898 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0898 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0898 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0898 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0898 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0898 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0898 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0898 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0898 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0898 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0898 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0898 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0898 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0898 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0898 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0898 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0898 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0898 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0898 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0898 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0898 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0898 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0898 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0898 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0898 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0898 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0898 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0898 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0898 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0898 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0898 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0898 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0898 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0898 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0898 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0898 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0898 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0898 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0898 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0898 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0898 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0898 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0898 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0898 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0898 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0898 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0473 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0473 [1], \xm8051_golden_model_1.sha_bytes_processed [1]);
  buf(\xm8051_golden_model_1.n0897 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0897 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0897 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0897 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0897 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0897 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0897 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0897 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0897 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0897 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0897 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0897 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0897 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0897 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0897 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0897 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0897 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0897 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0897 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0897 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0897 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0897 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0897 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0897 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0897 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0897 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0897 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0897 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0897 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0897 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0897 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0897 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0897 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0897 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0897 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0897 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0897 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0897 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0897 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0897 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0897 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0897 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0897 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0897 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0897 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0897 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0897 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0897 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0897 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0897 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0897 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0897 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0897 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0897 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0897 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0897 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0897 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0897 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0897 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0897 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0897 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0897 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0897 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0897 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0896 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0896 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0896 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0896 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0896 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0896 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0896 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0896 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0896 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0896 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0896 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0896 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0896 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0896 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0896 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0896 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0896 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0896 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0896 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0896 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0896 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0896 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0896 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0896 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0896 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0896 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0896 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0896 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0896 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0896 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0896 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0896 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0896 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0896 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0896 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0896 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0896 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0896 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0896 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0896 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0896 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0896 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0896 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0896 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0896 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0896 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0896 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0896 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0896 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0896 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0896 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0896 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0896 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0896 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0896 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0896 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0896 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0896 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0896 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0896 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0896 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0896 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0896 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0896 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0896 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0896 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0896 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0896 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0896 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0896 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0896 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0896 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0895 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0895 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0895 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0895 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0895 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0895 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0895 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0895 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0895 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0895 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0895 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0895 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0895 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0895 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0895 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0895 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0895 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0895 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0895 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0895 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0895 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0895 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0895 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0895 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0895 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0895 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0895 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0895 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0895 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0895 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0895 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0895 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0895 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0895 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0895 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0895 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0895 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0895 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0895 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0895 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0895 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0895 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0895 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0895 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0895 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0895 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0895 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0895 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0895 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0895 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0895 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0895 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0895 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0895 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0895 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0895 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0895 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0895 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0895 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0895 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0895 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0895 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0895 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0895 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0895 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0895 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0895 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0895 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0895 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0895 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0895 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0895 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0895 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0895 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0895 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0895 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0895 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0895 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0895 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0895 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0894 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0894 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0894 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0894 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0894 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0894 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0894 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0894 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0894 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0894 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0894 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0894 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0894 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0894 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0894 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0894 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0894 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0894 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0894 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0894 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0894 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0894 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0894 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0894 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0894 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0894 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0894 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0894 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0894 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0894 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0894 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0894 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0894 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0894 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0894 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0894 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0894 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0894 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0894 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0894 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0894 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0894 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0894 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0894 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0894 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0894 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0894 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0894 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0894 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0894 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0894 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0894 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0894 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0894 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0894 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0894 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0894 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0894 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0894 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0894 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0894 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0894 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0894 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0894 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0894 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0894 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0894 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0894 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0894 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0894 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0894 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0894 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0894 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0894 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0894 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0894 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0894 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0894 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0894 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0894 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0894 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0894 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0894 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0894 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0894 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0894 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0894 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0894 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0893 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0893 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0893 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0893 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0893 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0893 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0893 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0893 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0893 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0893 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0893 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0893 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0893 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0893 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0893 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0893 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0893 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0893 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0893 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0893 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0893 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0893 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0893 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0893 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0893 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0893 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0893 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0893 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0893 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0893 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0893 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0893 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0893 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0893 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0893 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0893 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0893 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0893 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0893 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0893 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0893 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0893 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0893 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0893 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0893 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0893 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0893 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0893 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0893 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0893 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0893 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0893 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0893 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0893 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0893 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0893 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0893 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0893 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0893 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0893 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0893 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0893 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0893 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0893 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0893 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0893 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0893 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0893 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0893 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0893 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0893 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0893 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0893 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0893 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0893 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0893 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0893 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0893 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0893 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0893 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0893 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0893 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0893 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0893 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0893 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0893 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0893 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0893 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0893 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0893 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0893 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0893 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0893 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0893 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0893 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0893 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0892 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0892 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0892 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0892 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0892 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0892 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0892 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0892 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0892 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0892 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0892 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0892 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0892 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0892 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0892 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0892 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0892 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0892 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0892 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0892 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0892 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0892 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0892 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0892 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0892 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0892 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0892 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0892 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0892 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0892 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0892 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0892 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0892 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0892 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0892 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0892 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0892 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0892 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0892 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0892 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0892 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0892 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0892 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0892 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0892 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0892 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0892 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0892 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0892 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0892 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0892 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0892 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0892 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0892 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0892 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0892 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0892 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0892 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0892 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0892 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0892 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0892 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0892 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0892 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0892 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0892 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0892 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0892 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0892 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0892 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0892 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0892 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0892 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0892 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0892 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0892 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0892 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0892 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0892 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0892 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0892 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0892 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0892 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0892 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0892 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0892 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0892 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0892 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0892 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0892 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0892 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0892 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0892 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0892 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0892 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0892 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0892 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0892 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0892 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0892 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0892 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0892 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0892 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0892 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0891 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0891 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0891 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0891 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0891 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0891 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0891 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0891 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0891 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0891 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0891 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0891 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0891 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0891 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0891 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0891 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0891 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0891 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0891 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0891 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0891 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0891 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0891 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0891 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0891 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0891 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0891 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0891 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0891 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0891 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0891 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0891 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0891 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0891 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0891 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0891 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0891 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0891 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0891 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0891 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0891 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0891 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0891 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0891 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0891 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0891 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0891 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0891 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0891 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0891 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0891 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0891 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0891 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0891 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0891 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0891 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0891 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0891 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0891 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0891 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0891 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0891 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0891 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0891 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0891 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0891 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0891 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0891 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0891 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0891 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0891 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0891 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0891 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0891 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0891 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0891 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0891 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0891 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0891 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0891 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0891 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0891 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0891 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0891 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0891 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0891 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0891 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0891 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0891 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0891 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0891 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0891 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0891 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0891 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0891 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0891 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0891 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0891 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0891 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0891 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0891 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0891 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0891 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0891 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0891 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0891 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0891 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0891 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0891 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0891 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0891 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0891 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0891 [120], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0891 [121], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0891 [122], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0891 [123], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0891 [124], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0891 [125], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0891 [126], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0891 [127], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0890 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0890 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0890 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0890 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0890 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0890 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0890 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0890 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0890 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0890 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0890 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0890 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0890 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0890 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0890 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0890 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0890 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0890 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0890 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0890 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0890 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0890 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0890 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0890 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0890 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0890 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0890 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0890 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0890 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0890 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0890 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0890 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0890 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0890 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0890 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0890 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0890 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0890 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0890 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0890 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0890 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0890 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0890 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0890 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0890 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0890 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0890 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0890 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0890 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0890 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0890 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0890 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0890 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0890 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0890 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0890 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0890 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0890 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0890 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0890 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0890 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0890 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0890 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0890 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0890 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0890 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0890 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0890 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0890 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0890 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0890 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0890 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0890 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0890 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0890 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0890 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0890 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0890 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0890 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0890 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0890 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0890 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0890 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0890 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0890 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0890 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0890 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0890 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0890 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0890 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0890 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0890 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0890 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0890 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0890 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0890 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0890 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0890 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0890 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0890 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0890 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0890 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0890 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0890 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0890 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0890 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0890 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0890 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0890 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0890 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0890 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0890 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0890 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0890 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0890 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0890 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0890 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0890 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0890 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0890 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [1], \xm8051_golden_model_1.aes_bytes_processed [1]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [2], \xm8051_golden_model_1.aes_bytes_processed [2]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [3], \xm8051_golden_model_1.aes_bytes_processed [3]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [4], \xm8051_golden_model_1.n0973 [4]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [5], \xm8051_golden_model_1.n0973 [5]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [6], \xm8051_golden_model_1.n0973 [6]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [7], \xm8051_golden_model_1.n0973 [7]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [8], \xm8051_golden_model_1.n0973 [8]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [9], \xm8051_golden_model_1.n0973 [9]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [10], \xm8051_golden_model_1.n0973 [10]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [11], \xm8051_golden_model_1.n0973 [11]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [12], \xm8051_golden_model_1.n0973 [12]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [13], \xm8051_golden_model_1.n0973 [13]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [14], \xm8051_golden_model_1.n0973 [14]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0f [15], \xm8051_golden_model_1.n0973 [15]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [1], \xm8051_golden_model_1.aes_bytes_processed [1]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [2], \xm8051_golden_model_1.aes_bytes_processed [2]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [3], \xm8051_golden_model_1.aes_bytes_processed [3]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [4], \xm8051_golden_model_1.n0973 [4]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [5], \xm8051_golden_model_1.n0973 [5]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [6], \xm8051_golden_model_1.n0973 [6]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [7], \xm8051_golden_model_1.n0973 [7]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [8], \xm8051_golden_model_1.n0973 [8]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [9], \xm8051_golden_model_1.n0973 [9]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [10], \xm8051_golden_model_1.n0973 [10]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [11], \xm8051_golden_model_1.n0973 [11]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [12], \xm8051_golden_model_1.n0973 [12]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [13], \xm8051_golden_model_1.n0973 [13]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [14], \xm8051_golden_model_1.n0973 [14]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_0b [15], \xm8051_golden_model_1.n0973 [15]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [1], \xm8051_golden_model_1.aes_bytes_processed [1]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [2], \xm8051_golden_model_1.aes_bytes_processed [2]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [3], \xm8051_golden_model_1.aes_bytes_processed [3]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [4], \xm8051_golden_model_1.n0973 [4]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [5], \xm8051_golden_model_1.n0973 [5]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [6], \xm8051_golden_model_1.n0973 [6]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [7], \xm8051_golden_model_1.n0973 [7]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [8], \xm8051_golden_model_1.n0973 [8]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [9], \xm8051_golden_model_1.n0973 [9]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [10], \xm8051_golden_model_1.n0973 [10]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [11], \xm8051_golden_model_1.n0973 [11]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [12], \xm8051_golden_model_1.n0973 [12]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [13], \xm8051_golden_model_1.n0973 [13]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [14], \xm8051_golden_model_1.n0973 [14]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_07 [15], \xm8051_golden_model_1.n0973 [15]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [0], \xm8051_golden_model_1.aes_bytes_processed [0]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [1], \xm8051_golden_model_1.aes_bytes_processed [1]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [2], \xm8051_golden_model_1.aes_bytes_processed [2]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [3], \xm8051_golden_model_1.aes_bytes_processed [3]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [4], \xm8051_golden_model_1.n0973 [4]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [5], \xm8051_golden_model_1.n0973 [5]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [6], \xm8051_golden_model_1.n0973 [6]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [7], \xm8051_golden_model_1.n0973 [7]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [8], \xm8051_golden_model_1.n0973 [8]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [9], \xm8051_golden_model_1.n0973 [9]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [10], \xm8051_golden_model_1.n0973 [10]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [11], \xm8051_golden_model_1.n0973 [11]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [12], \xm8051_golden_model_1.n0973 [12]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [13], \xm8051_golden_model_1.n0973 [13]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [14], \xm8051_golden_model_1.n0973 [14]);
  buf(\xm8051_golden_model_1.aes_bytes_processed_03 [15], \xm8051_golden_model_1.n0973 [15]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [9], ABINPUT[9]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [10], ABINPUT[10]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [11], ABINPUT[11]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [12], ABINPUT[12]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [13], ABINPUT[13]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [14], ABINPUT[14]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [15], ABINPUT[15]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [16], ABINPUT[16]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [17], ABINPUT[17]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [18], ABINPUT[18]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [19], ABINPUT[19]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [20], ABINPUT[20]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [21], ABINPUT[21]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [22], ABINPUT[22]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [23], ABINPUT[23]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [24], ABINPUT[24]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [25], ABINPUT[25]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [26], ABINPUT[26]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [27], ABINPUT[27]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [28], ABINPUT[28]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [29], ABINPUT[29]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [30], ABINPUT[30]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [31], ABINPUT[31]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [32], ABINPUT[32]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [33], ABINPUT[33]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [34], ABINPUT[34]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [35], ABINPUT[35]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [36], ABINPUT[36]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [37], ABINPUT[37]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [38], ABINPUT[38]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [39], ABINPUT[39]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [40], ABINPUT[40]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [41], ABINPUT[41]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [42], ABINPUT[42]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [43], ABINPUT[43]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [44], ABINPUT[44]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [45], ABINPUT[45]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [46], ABINPUT[46]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [47], ABINPUT[47]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [48], ABINPUT[48]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [49], ABINPUT[49]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [50], ABINPUT[50]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [51], ABINPUT[51]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [52], ABINPUT[52]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [53], ABINPUT[53]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [54], ABINPUT[54]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [55], ABINPUT[55]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [56], ABINPUT[56]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [57], ABINPUT[57]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [58], ABINPUT[58]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [59], ABINPUT[59]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [60], ABINPUT[60]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [61], ABINPUT[61]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [62], ABINPUT[62]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [63], ABINPUT[63]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [64], ABINPUT[64]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [65], ABINPUT[65]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [66], ABINPUT[66]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [67], ABINPUT[67]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [68], ABINPUT[68]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [69], ABINPUT[69]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [70], ABINPUT[70]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [71], ABINPUT[71]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [72], ABINPUT[72]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [73], ABINPUT[73]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [74], ABINPUT[74]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [75], ABINPUT[75]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [76], ABINPUT[76]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [77], ABINPUT[77]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [78], ABINPUT[78]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [79], ABINPUT[79]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [80], ABINPUT[80]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [81], ABINPUT[81]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [82], ABINPUT[82]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [83], ABINPUT[83]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [84], ABINPUT[84]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [85], ABINPUT[85]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [86], ABINPUT[86]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [87], ABINPUT[87]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [88], ABINPUT[88]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [89], ABINPUT[89]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [90], ABINPUT[90]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [91], ABINPUT[91]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [92], ABINPUT[92]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [93], ABINPUT[93]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [94], ABINPUT[94]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [95], ABINPUT[95]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [96], ABINPUT[96]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [97], ABINPUT[97]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [98], ABINPUT[98]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [99], ABINPUT[99]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [100], ABINPUT[100]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [101], ABINPUT[101]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [102], ABINPUT[102]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [103], ABINPUT[103]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [104], ABINPUT[104]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [105], ABINPUT[105]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [106], ABINPUT[106]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [107], ABINPUT[107]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [108], ABINPUT[108]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [109], ABINPUT[109]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [110], ABINPUT[110]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [111], ABINPUT[111]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [112], ABINPUT[112]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [113], ABINPUT[113]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [114], ABINPUT[114]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [115], ABINPUT[115]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [116], ABINPUT[116]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [117], ABINPUT[117]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [118], ABINPUT[118]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [119], ABINPUT[119]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [120], ABINPUT[120]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [121], ABINPUT[121]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [122], ABINPUT[122]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [123], ABINPUT[123]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [124], ABINPUT[124]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [125], ABINPUT[125]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [126], ABINPUT[126]);
  buf(\oc8051_xiommu_impl_1.ABINPUT [127], ABINPUT[127]);
  buf(\oc8051_xiommu_impl_1.clk , clk);
  buf(\oc8051_xiommu_impl_1.rst , rst);
  buf(\oc8051_xiommu_impl_1.proc_wr , proc_wr);
  buf(\oc8051_xiommu_impl_1.proc_stb , proc_stb);
  buf(\oc8051_xiommu_impl_1.proc_data_in [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.proc_data_in [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.proc_data_in [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.proc_data_in [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.proc_data_in [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.proc_data_in [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.proc_data_in [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.proc_data_in [7], proc_data_in[7]);
  buf(\oc8051_xiommu_impl_1.proc_addr [0], proc_addr[0]);
  buf(\oc8051_xiommu_impl_1.proc_addr [1], proc_addr[1]);
  buf(\oc8051_xiommu_impl_1.proc_addr [2], proc_addr[2]);
  buf(\oc8051_xiommu_impl_1.proc_addr [3], proc_addr[3]);
  buf(\oc8051_xiommu_impl_1.proc_addr [4], proc_addr[4]);
  buf(\oc8051_xiommu_impl_1.proc_addr [5], proc_addr[5]);
  buf(\oc8051_xiommu_impl_1.proc_addr [6], proc_addr[6]);
  buf(\oc8051_xiommu_impl_1.proc_addr [7], proc_addr[7]);
  buf(\oc8051_xiommu_impl_1.proc_addr [8], proc_addr[8]);
  buf(\oc8051_xiommu_impl_1.proc_addr [9], proc_addr[9]);
  buf(\oc8051_xiommu_impl_1.proc_addr [10], proc_addr[10]);
  buf(\oc8051_xiommu_impl_1.proc_addr [11], proc_addr[11]);
  buf(\oc8051_xiommu_impl_1.proc_addr [12], proc_addr[12]);
  buf(\oc8051_xiommu_impl_1.proc_addr [13], proc_addr[13]);
  buf(\oc8051_xiommu_impl_1.proc_addr [14], proc_addr[14]);
  buf(\oc8051_xiommu_impl_1.proc_addr [15], proc_addr[15]);
  buf(\oc8051_xiommu_impl_1.aes_state [0], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [0]);
  buf(\oc8051_xiommu_impl_1.aes_state [1], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [1]);
  buf(\oc8051_xiommu_impl_1.sha_state [0], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0]);
  buf(\oc8051_xiommu_impl_1.sha_state [1], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [1]);
  buf(\oc8051_xiommu_impl_1.aes_len [0], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [0]);
  buf(\oc8051_xiommu_impl_1.aes_len [1], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [1]);
  buf(\oc8051_xiommu_impl_1.aes_len [2], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [2]);
  buf(\oc8051_xiommu_impl_1.aes_len [3], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [3]);
  buf(\oc8051_xiommu_impl_1.aes_len [4], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [4]);
  buf(\oc8051_xiommu_impl_1.aes_len [5], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [5]);
  buf(\oc8051_xiommu_impl_1.aes_len [6], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [6]);
  buf(\oc8051_xiommu_impl_1.aes_len [7], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [7]);
  buf(\oc8051_xiommu_impl_1.aes_len [8], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [8]);
  buf(\oc8051_xiommu_impl_1.aes_len [9], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [9]);
  buf(\oc8051_xiommu_impl_1.aes_len [10], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [10]);
  buf(\oc8051_xiommu_impl_1.aes_len [11], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [11]);
  buf(\oc8051_xiommu_impl_1.aes_len [12], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [12]);
  buf(\oc8051_xiommu_impl_1.aes_len [13], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [13]);
  buf(\oc8051_xiommu_impl_1.aes_len [14], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [14]);
  buf(\oc8051_xiommu_impl_1.aes_len [15], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [15]);
  buf(\oc8051_xiommu_impl_1.sha_len [0], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [0]);
  buf(\oc8051_xiommu_impl_1.sha_len [1], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [1]);
  buf(\oc8051_xiommu_impl_1.sha_len [2], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [2]);
  buf(\oc8051_xiommu_impl_1.sha_len [3], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [3]);
  buf(\oc8051_xiommu_impl_1.sha_len [4], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [4]);
  buf(\oc8051_xiommu_impl_1.sha_len [5], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [5]);
  buf(\oc8051_xiommu_impl_1.sha_len [6], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [6]);
  buf(\oc8051_xiommu_impl_1.sha_len [7], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [7]);
  buf(\oc8051_xiommu_impl_1.sha_len [8], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [8]);
  buf(\oc8051_xiommu_impl_1.sha_len [9], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [9]);
  buf(\oc8051_xiommu_impl_1.sha_len [10], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [10]);
  buf(\oc8051_xiommu_impl_1.sha_len [11], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [11]);
  buf(\oc8051_xiommu_impl_1.sha_len [12], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [12]);
  buf(\oc8051_xiommu_impl_1.sha_len [13], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [13]);
  buf(\oc8051_xiommu_impl_1.sha_len [14], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [14]);
  buf(\oc8051_xiommu_impl_1.sha_len [15], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [15]);
  buf(\xm8051_golden_model_1.n0889 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0889 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0889 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0889 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0889 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0889 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0889 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0889 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0889 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0889 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0889 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0889 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0889 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0889 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0889 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0889 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0889 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0889 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0889 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0889 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0889 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0889 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0889 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0889 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0889 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0889 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0889 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0889 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0889 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0889 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0889 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0889 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0889 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0889 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0889 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0889 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0889 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0889 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0889 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0889 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0889 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0889 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0889 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0889 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0889 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0889 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0889 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0889 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0889 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0889 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0889 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0889 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0889 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0889 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0889 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0889 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0889 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0889 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0889 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0889 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0889 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0889 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0889 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0889 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0889 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0889 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0889 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0889 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0889 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0889 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0889 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0889 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0889 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0889 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0889 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0889 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0889 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0889 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0889 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0889 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0889 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0889 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0889 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0889 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0889 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0889 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0889 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0889 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0889 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0889 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0889 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0889 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0889 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0889 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0889 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0889 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0889 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0889 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0889 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0889 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0889 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0889 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0889 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0889 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0889 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0889 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0889 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0889 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0889 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0889 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0889 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0889 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0889 [112], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0889 [113], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0889 [114], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0889 [115], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0889 [116], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0889 [117], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0889 [118], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0889 [119], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0463 [0], \xm8051_golden_model_1.sha_bytes_processed [0]);
  buf(\xm8051_golden_model_1.n0463 [1], \xm8051_golden_model_1.n0483 [1]);
  buf(\xm8051_golden_model_1.n0888 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0888 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0888 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0888 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0888 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0888 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0888 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0888 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0888 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0888 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0888 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0888 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0888 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0888 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0888 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0888 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0888 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0888 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0888 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0888 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0888 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0888 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0888 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0888 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0888 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0888 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0888 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0888 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0888 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0888 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0888 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0888 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0888 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0888 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0888 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0888 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0888 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0888 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0888 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0888 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0888 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0888 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0888 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0888 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0888 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0888 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0888 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0888 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0888 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0888 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0888 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0888 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0888 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0888 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0888 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0888 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0888 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0888 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0888 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0888 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0888 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0888 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0888 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0888 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0888 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0888 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0888 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0888 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0888 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0888 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0888 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0888 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0888 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0888 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0888 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0888 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0888 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0888 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0888 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0888 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0888 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0888 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0888 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0888 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0888 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0888 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0888 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0888 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0888 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0888 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0888 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0888 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0888 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0888 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0888 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0888 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0888 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0888 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0888 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0888 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0888 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0888 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0888 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0888 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0888 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0888 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0888 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0888 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0888 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0888 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0888 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0888 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0887 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0887 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0887 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0887 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0887 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0887 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0887 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0887 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0887 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0887 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0887 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0887 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0887 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0887 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0887 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0887 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0887 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0887 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0887 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0887 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0887 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0887 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0887 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0887 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0887 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0887 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0887 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0887 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0887 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0887 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0887 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0887 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0887 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0887 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0887 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0887 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0887 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0887 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0887 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0887 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0887 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0887 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0887 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0887 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0887 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0887 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0887 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0887 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0887 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0887 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0887 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0887 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0887 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0887 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0887 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0887 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0887 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0887 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0887 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0887 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0887 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0887 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0887 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0887 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0887 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0887 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0887 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0887 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0887 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0887 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0887 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0887 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0887 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0887 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0887 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0887 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0887 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0887 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0887 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0887 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0887 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0887 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0887 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0887 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0887 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0887 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0887 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0887 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0887 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0887 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0887 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0887 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0887 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0887 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0887 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0887 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0887 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0887 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0887 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0887 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0887 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0887 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0887 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0887 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\xm8051_golden_model_1.n0887 [104], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0887 [105], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0887 [106], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0887 [107], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0887 [108], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0887 [109], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0887 [110], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0887 [111], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0887 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0887 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0887 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0887 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0887 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0887 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0887 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0887 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0887 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0887 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0887 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0887 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0887 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0887 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0887 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0887 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0886 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0886 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0886 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0886 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0886 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0886 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0886 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0886 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0886 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0886 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0886 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0886 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0886 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0886 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0886 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0886 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0886 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0886 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0886 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0886 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0886 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0886 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0886 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0886 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0886 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0886 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0886 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0886 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0886 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0886 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0886 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0886 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0886 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0886 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0886 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0886 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0886 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0886 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0886 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0886 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0886 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0886 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0886 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0886 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0886 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0886 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0886 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0886 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0886 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0886 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0886 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0886 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0886 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0886 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0886 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0886 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0886 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0886 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0886 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0886 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0886 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0886 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0886 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0886 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0886 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0886 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0886 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0886 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0886 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0886 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0886 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0886 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0886 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0886 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0886 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0886 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0886 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0886 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0886 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0886 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0886 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0886 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0886 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0886 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0886 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0886 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0886 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0886 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0886 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0886 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0886 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0886 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0886 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0886 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0886 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0886 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0886 [96], \xm8051_golden_model_1.n0893 [96]);
  buf(\xm8051_golden_model_1.n0886 [97], \xm8051_golden_model_1.n0893 [97]);
  buf(\xm8051_golden_model_1.n0886 [98], \xm8051_golden_model_1.n0893 [98]);
  buf(\xm8051_golden_model_1.n0886 [99], \xm8051_golden_model_1.n0893 [99]);
  buf(\xm8051_golden_model_1.n0886 [100], \xm8051_golden_model_1.n0893 [100]);
  buf(\xm8051_golden_model_1.n0886 [101], \xm8051_golden_model_1.n0893 [101]);
  buf(\xm8051_golden_model_1.n0886 [102], \xm8051_golden_model_1.n0893 [102]);
  buf(\xm8051_golden_model_1.n0886 [103], \xm8051_golden_model_1.n0893 [103]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [0], ABINPUT000[0]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [1], ABINPUT000[1]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [2], ABINPUT000[2]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [3], ABINPUT000[3]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [4], ABINPUT000[4]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [5], ABINPUT000[5]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [6], ABINPUT000[6]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [7], ABINPUT000[7]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [8], ABINPUT000[8]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [9], ABINPUT000[9]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [10], ABINPUT000[10]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [11], ABINPUT000[11]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [12], ABINPUT000[12]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [13], ABINPUT000[13]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [14], ABINPUT000[14]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [15], ABINPUT000[15]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [16], ABINPUT000[16]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [17], ABINPUT000[17]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [18], ABINPUT000[18]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [19], ABINPUT000[19]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [20], ABINPUT000[20]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [21], ABINPUT000[21]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [22], ABINPUT000[22]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [23], ABINPUT000[23]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [24], ABINPUT000[24]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [25], ABINPUT000[25]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [26], ABINPUT000[26]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [27], ABINPUT000[27]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [28], ABINPUT000[28]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [29], ABINPUT000[29]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [30], ABINPUT000[30]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [31], ABINPUT000[31]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [32], ABINPUT000[32]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [33], ABINPUT000[33]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [34], ABINPUT000[34]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [35], ABINPUT000[35]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [36], ABINPUT000[36]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [37], ABINPUT000[37]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [38], ABINPUT000[38]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [39], ABINPUT000[39]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [40], ABINPUT000[40]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [41], ABINPUT000[41]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [42], ABINPUT000[42]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [43], ABINPUT000[43]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [44], ABINPUT000[44]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [45], ABINPUT000[45]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [46], ABINPUT000[46]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [47], ABINPUT000[47]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [48], ABINPUT000[48]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [49], ABINPUT000[49]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [50], ABINPUT000[50]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [51], ABINPUT000[51]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [52], ABINPUT000[52]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [53], ABINPUT000[53]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [54], ABINPUT000[54]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [55], ABINPUT000[55]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [56], ABINPUT000[56]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [57], ABINPUT000[57]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [58], ABINPUT000[58]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [59], ABINPUT000[59]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [60], ABINPUT000[60]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [61], ABINPUT000[61]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [62], ABINPUT000[62]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [63], ABINPUT000[63]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [64], ABINPUT000[64]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [65], ABINPUT000[65]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [66], ABINPUT000[66]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [67], ABINPUT000[67]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [68], ABINPUT000[68]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [69], ABINPUT000[69]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [70], ABINPUT000[70]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [71], ABINPUT000[71]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [72], ABINPUT000[72]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [73], ABINPUT000[73]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [74], ABINPUT000[74]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [75], ABINPUT000[75]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [76], ABINPUT000[76]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [77], ABINPUT000[77]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [78], ABINPUT000[78]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [79], ABINPUT000[79]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [80], ABINPUT000[80]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [81], ABINPUT000[81]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [82], ABINPUT000[82]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [83], ABINPUT000[83]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [84], ABINPUT000[84]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [85], ABINPUT000[85]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [86], ABINPUT000[86]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [87], ABINPUT000[87]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [88], ABINPUT000[88]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [89], ABINPUT000[89]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [90], ABINPUT000[90]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [91], ABINPUT000[91]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [92], ABINPUT000[92]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [93], ABINPUT000[93]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [94], ABINPUT000[94]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [95], ABINPUT000[95]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [96], ABINPUT000[96]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [97], ABINPUT000[97]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [98], ABINPUT000[98]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [99], ABINPUT000[99]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [100], ABINPUT000[100]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [101], ABINPUT000[101]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [102], ABINPUT000[102]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [103], ABINPUT000[103]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [104], ABINPUT000[104]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [105], ABINPUT000[105]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [106], ABINPUT000[106]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [107], ABINPUT000[107]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [108], ABINPUT000[108]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [109], ABINPUT000[109]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [110], ABINPUT000[110]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [111], ABINPUT000[111]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [112], ABINPUT000[112]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [113], ABINPUT000[113]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [114], ABINPUT000[114]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [115], ABINPUT000[115]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [116], ABINPUT000[116]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [117], ABINPUT000[117]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [118], ABINPUT000[118]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [119], ABINPUT000[119]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [120], ABINPUT000[120]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [121], ABINPUT000[121]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [122], ABINPUT000[122]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [123], ABINPUT000[123]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [124], ABINPUT000[124]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [125], ABINPUT000[125]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [126], ABINPUT000[126]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [127], ABINPUT000[127]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [128], ABINPUT000[128]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [129], ABINPUT000[129]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [130], ABINPUT000[130]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [131], ABINPUT000[131]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [132], ABINPUT000[132]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [133], ABINPUT000[133]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [134], ABINPUT000[134]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [135], ABINPUT000[135]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [136], ABINPUT000[136]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [137], ABINPUT000[137]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [138], ABINPUT000[138]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [139], ABINPUT000[139]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [140], ABINPUT000[140]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [141], ABINPUT000[141]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [142], ABINPUT000[142]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [143], ABINPUT000[143]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [144], ABINPUT000[144]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [145], ABINPUT000[145]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [146], ABINPUT000[146]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [147], ABINPUT000[147]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [148], ABINPUT000[148]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [149], ABINPUT000[149]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [150], ABINPUT000[150]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [151], ABINPUT000[151]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [152], ABINPUT000[152]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [153], ABINPUT000[153]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [154], ABINPUT000[154]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [155], ABINPUT000[155]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [156], ABINPUT000[156]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [157], ABINPUT000[157]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [158], ABINPUT000[158]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [159], ABINPUT000[159]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [160], ABINPUT000[160]);
  buf(\oc8051_xiommu_impl_1.ABINPUT000 [161], ABINPUT000[161]);
  buf(sha_state_gm[0], \xm8051_golden_model_1.sha_state [0]);
  buf(sha_state_gm[1], \xm8051_golden_model_1.sha_state [1]);
  buf(sha_state_gm[2], \xm8051_golden_model_1.sha_state [2]);
  buf(sha_state_gm[3], \xm8051_golden_model_1.sha_state [3]);
  buf(sha_state_gm[4], \xm8051_golden_model_1.sha_state [4]);
  buf(sha_state_gm[5], \xm8051_golden_model_1.sha_state [5]);
  buf(sha_state_gm[6], \xm8051_golden_model_1.sha_state [6]);
  buf(sha_state_gm[7], \xm8051_golden_model_1.sha_state [7]);
  buf(aes_state_gm[0], \xm8051_golden_model_1.aes_state [0]);
  buf(aes_state_gm[1], \xm8051_golden_model_1.aes_state [1]);
  buf(aes_state_gm[2], \xm8051_golden_model_1.aes_state [2]);
  buf(aes_state_gm[3], \xm8051_golden_model_1.aes_state [3]);
  buf(aes_state_gm[4], \xm8051_golden_model_1.aes_state [4]);
  buf(aes_state_gm[5], \xm8051_golden_model_1.aes_state [5]);
  buf(aes_state_gm[6], \xm8051_golden_model_1.aes_state [6]);
  buf(aes_state_gm[7], \xm8051_golden_model_1.aes_state [7]);
  buf(sha_len_gm[0], \xm8051_golden_model_1.sha_len [0]);
  buf(sha_len_gm[1], \xm8051_golden_model_1.sha_len [1]);
  buf(sha_len_gm[2], \xm8051_golden_model_1.sha_len [2]);
  buf(sha_len_gm[3], \xm8051_golden_model_1.sha_len [3]);
  buf(sha_len_gm[4], \xm8051_golden_model_1.sha_len [4]);
  buf(sha_len_gm[5], \xm8051_golden_model_1.sha_len [5]);
  buf(sha_len_gm[6], \xm8051_golden_model_1.sha_len [6]);
  buf(sha_len_gm[7], \xm8051_golden_model_1.sha_len [7]);
  buf(sha_len_gm[8], \xm8051_golden_model_1.sha_len [8]);
  buf(sha_len_gm[9], \xm8051_golden_model_1.sha_len [9]);
  buf(sha_len_gm[10], \xm8051_golden_model_1.sha_len [10]);
  buf(sha_len_gm[11], \xm8051_golden_model_1.sha_len [11]);
  buf(sha_len_gm[12], \xm8051_golden_model_1.sha_len [12]);
  buf(sha_len_gm[13], \xm8051_golden_model_1.sha_len [13]);
  buf(sha_len_gm[14], \xm8051_golden_model_1.sha_len [14]);
  buf(sha_len_gm[15], \xm8051_golden_model_1.sha_len [15]);
  buf(aes_len_gm[0], \xm8051_golden_model_1.aes_len [0]);
  buf(aes_len_gm[1], \xm8051_golden_model_1.aes_len [1]);
  buf(aes_len_gm[2], \xm8051_golden_model_1.aes_len [2]);
  buf(aes_len_gm[3], \xm8051_golden_model_1.aes_len [3]);
  buf(aes_len_gm[4], \xm8051_golden_model_1.aes_len [4]);
  buf(aes_len_gm[5], \xm8051_golden_model_1.aes_len [5]);
  buf(aes_len_gm[6], \xm8051_golden_model_1.aes_len [6]);
  buf(aes_len_gm[7], \xm8051_golden_model_1.aes_len [7]);
  buf(aes_len_gm[8], \xm8051_golden_model_1.aes_len [8]);
  buf(aes_len_gm[9], \xm8051_golden_model_1.aes_len [9]);
  buf(aes_len_gm[10], \xm8051_golden_model_1.aes_len [10]);
  buf(aes_len_gm[11], \xm8051_golden_model_1.aes_len [11]);
  buf(aes_len_gm[12], \xm8051_golden_model_1.aes_len [12]);
  buf(aes_len_gm[13], \xm8051_golden_model_1.aes_len [13]);
  buf(aes_len_gm[14], \xm8051_golden_model_1.aes_len [14]);
  buf(aes_len_gm[15], \xm8051_golden_model_1.aes_len [15]);
  buf(sha_len_impl[0], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [0]);
  buf(sha_len_impl[1], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [1]);
  buf(sha_len_impl[2], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [2]);
  buf(sha_len_impl[3], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [3]);
  buf(sha_len_impl[4], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [4]);
  buf(sha_len_impl[5], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [5]);
  buf(sha_len_impl[6], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [6]);
  buf(sha_len_impl[7], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [7]);
  buf(sha_len_impl[8], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [8]);
  buf(sha_len_impl[9], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [9]);
  buf(sha_len_impl[10], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [10]);
  buf(sha_len_impl[11], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [11]);
  buf(sha_len_impl[12], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [12]);
  buf(sha_len_impl[13], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [13]);
  buf(sha_len_impl[14], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [14]);
  buf(sha_len_impl[15], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_len_i.reg_out [15]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.data_in [0], proc_data_in[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.data_in [1], proc_data_in[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.data_in [2], proc_data_in[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.data_in [3], proc_data_in[3]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.data_in [4], proc_data_in[4]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.data_in [5], proc_data_in[5]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.data_in [6], proc_data_in[6]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.data_in [7], proc_data_in[7]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.addr [0], proc_addr[0]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.addr [1], proc_addr[1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.addr [2], proc_addr[2]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.addr [3], proc_addr[3]);
  buf(aes_len_impl[0], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [0]);
  buf(aes_len_impl[1], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [1]);
  buf(aes_len_impl[2], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [2]);
  buf(aes_len_impl[3], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [3]);
  buf(aes_len_impl[4], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [4]);
  buf(aes_len_impl[5], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [5]);
  buf(aes_len_impl[6], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [6]);
  buf(aes_len_impl[7], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [7]);
  buf(aes_len_impl[8], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [8]);
  buf(aes_len_impl[9], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [9]);
  buf(aes_len_impl[10], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [10]);
  buf(aes_len_impl[11], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [11]);
  buf(aes_len_impl[12], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [12]);
  buf(aes_len_impl[13], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [13]);
  buf(aes_len_impl[14], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [14]);
  buf(aes_len_impl[15], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_oplen_i.reg_out [15]);
  buf(\xm8051_golden_model_1.n0885 [0], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0885 [1], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0885 [2], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0885 [3], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0885 [4], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0885 [5], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0885 [6], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0885 [7], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0885 [8], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0885 [9], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0885 [10], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0885 [11], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0885 [12], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0885 [13], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0885 [14], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0885 [15], \xm8051_golden_model_1.n0889 [127]);
  buf(\xm8051_golden_model_1.n0884 [0], \xm8051_golden_model_1.n0905 [0]);
  buf(\xm8051_golden_model_1.n0884 [1], \xm8051_golden_model_1.n0905 [1]);
  buf(\xm8051_golden_model_1.n0884 [2], \xm8051_golden_model_1.n0905 [2]);
  buf(\xm8051_golden_model_1.n0884 [3], \xm8051_golden_model_1.n0905 [3]);
  buf(\xm8051_golden_model_1.n0884 [4], \xm8051_golden_model_1.n0905 [4]);
  buf(\xm8051_golden_model_1.n0884 [5], \xm8051_golden_model_1.n0905 [5]);
  buf(\xm8051_golden_model_1.n0884 [6], \xm8051_golden_model_1.n0905 [6]);
  buf(\xm8051_golden_model_1.n0884 [7], \xm8051_golden_model_1.n0905 [7]);
  buf(\xm8051_golden_model_1.n0884 [8], \xm8051_golden_model_1.n0904 [8]);
  buf(\xm8051_golden_model_1.n0884 [9], \xm8051_golden_model_1.n0904 [9]);
  buf(\xm8051_golden_model_1.n0884 [10], \xm8051_golden_model_1.n0904 [10]);
  buf(\xm8051_golden_model_1.n0884 [11], \xm8051_golden_model_1.n0904 [11]);
  buf(\xm8051_golden_model_1.n0884 [12], \xm8051_golden_model_1.n0904 [12]);
  buf(\xm8051_golden_model_1.n0884 [13], \xm8051_golden_model_1.n0904 [13]);
  buf(\xm8051_golden_model_1.n0884 [14], \xm8051_golden_model_1.n0904 [14]);
  buf(\xm8051_golden_model_1.n0884 [15], \xm8051_golden_model_1.n0904 [15]);
  buf(\xm8051_golden_model_1.n0884 [16], \xm8051_golden_model_1.n0903 [16]);
  buf(\xm8051_golden_model_1.n0884 [17], \xm8051_golden_model_1.n0903 [17]);
  buf(\xm8051_golden_model_1.n0884 [18], \xm8051_golden_model_1.n0903 [18]);
  buf(\xm8051_golden_model_1.n0884 [19], \xm8051_golden_model_1.n0903 [19]);
  buf(\xm8051_golden_model_1.n0884 [20], \xm8051_golden_model_1.n0903 [20]);
  buf(\xm8051_golden_model_1.n0884 [21], \xm8051_golden_model_1.n0903 [21]);
  buf(\xm8051_golden_model_1.n0884 [22], \xm8051_golden_model_1.n0903 [22]);
  buf(\xm8051_golden_model_1.n0884 [23], \xm8051_golden_model_1.n0903 [23]);
  buf(\xm8051_golden_model_1.n0884 [24], \xm8051_golden_model_1.n0902 [24]);
  buf(\xm8051_golden_model_1.n0884 [25], \xm8051_golden_model_1.n0902 [25]);
  buf(\xm8051_golden_model_1.n0884 [26], \xm8051_golden_model_1.n0902 [26]);
  buf(\xm8051_golden_model_1.n0884 [27], \xm8051_golden_model_1.n0902 [27]);
  buf(\xm8051_golden_model_1.n0884 [28], \xm8051_golden_model_1.n0902 [28]);
  buf(\xm8051_golden_model_1.n0884 [29], \xm8051_golden_model_1.n0902 [29]);
  buf(\xm8051_golden_model_1.n0884 [30], \xm8051_golden_model_1.n0902 [30]);
  buf(\xm8051_golden_model_1.n0884 [31], \xm8051_golden_model_1.n0902 [31]);
  buf(\xm8051_golden_model_1.n0884 [32], \xm8051_golden_model_1.n0901 [32]);
  buf(\xm8051_golden_model_1.n0884 [33], \xm8051_golden_model_1.n0901 [33]);
  buf(\xm8051_golden_model_1.n0884 [34], \xm8051_golden_model_1.n0901 [34]);
  buf(\xm8051_golden_model_1.n0884 [35], \xm8051_golden_model_1.n0901 [35]);
  buf(\xm8051_golden_model_1.n0884 [36], \xm8051_golden_model_1.n0901 [36]);
  buf(\xm8051_golden_model_1.n0884 [37], \xm8051_golden_model_1.n0901 [37]);
  buf(\xm8051_golden_model_1.n0884 [38], \xm8051_golden_model_1.n0901 [38]);
  buf(\xm8051_golden_model_1.n0884 [39], \xm8051_golden_model_1.n0901 [39]);
  buf(\xm8051_golden_model_1.n0884 [40], \xm8051_golden_model_1.n0900 [40]);
  buf(\xm8051_golden_model_1.n0884 [41], \xm8051_golden_model_1.n0900 [41]);
  buf(\xm8051_golden_model_1.n0884 [42], \xm8051_golden_model_1.n0900 [42]);
  buf(\xm8051_golden_model_1.n0884 [43], \xm8051_golden_model_1.n0900 [43]);
  buf(\xm8051_golden_model_1.n0884 [44], \xm8051_golden_model_1.n0900 [44]);
  buf(\xm8051_golden_model_1.n0884 [45], \xm8051_golden_model_1.n0900 [45]);
  buf(\xm8051_golden_model_1.n0884 [46], \xm8051_golden_model_1.n0900 [46]);
  buf(\xm8051_golden_model_1.n0884 [47], \xm8051_golden_model_1.n0900 [47]);
  buf(\xm8051_golden_model_1.n0884 [48], \xm8051_golden_model_1.n0899 [48]);
  buf(\xm8051_golden_model_1.n0884 [49], \xm8051_golden_model_1.n0899 [49]);
  buf(\xm8051_golden_model_1.n0884 [50], \xm8051_golden_model_1.n0899 [50]);
  buf(\xm8051_golden_model_1.n0884 [51], \xm8051_golden_model_1.n0899 [51]);
  buf(\xm8051_golden_model_1.n0884 [52], \xm8051_golden_model_1.n0899 [52]);
  buf(\xm8051_golden_model_1.n0884 [53], \xm8051_golden_model_1.n0899 [53]);
  buf(\xm8051_golden_model_1.n0884 [54], \xm8051_golden_model_1.n0899 [54]);
  buf(\xm8051_golden_model_1.n0884 [55], \xm8051_golden_model_1.n0899 [55]);
  buf(\xm8051_golden_model_1.n0884 [56], \xm8051_golden_model_1.n0898 [56]);
  buf(\xm8051_golden_model_1.n0884 [57], \xm8051_golden_model_1.n0898 [57]);
  buf(\xm8051_golden_model_1.n0884 [58], \xm8051_golden_model_1.n0898 [58]);
  buf(\xm8051_golden_model_1.n0884 [59], \xm8051_golden_model_1.n0898 [59]);
  buf(\xm8051_golden_model_1.n0884 [60], \xm8051_golden_model_1.n0898 [60]);
  buf(\xm8051_golden_model_1.n0884 [61], \xm8051_golden_model_1.n0898 [61]);
  buf(\xm8051_golden_model_1.n0884 [62], \xm8051_golden_model_1.n0898 [62]);
  buf(\xm8051_golden_model_1.n0884 [63], \xm8051_golden_model_1.n0898 [63]);
  buf(\xm8051_golden_model_1.n0884 [64], \xm8051_golden_model_1.n0897 [64]);
  buf(\xm8051_golden_model_1.n0884 [65], \xm8051_golden_model_1.n0897 [65]);
  buf(\xm8051_golden_model_1.n0884 [66], \xm8051_golden_model_1.n0897 [66]);
  buf(\xm8051_golden_model_1.n0884 [67], \xm8051_golden_model_1.n0897 [67]);
  buf(\xm8051_golden_model_1.n0884 [68], \xm8051_golden_model_1.n0897 [68]);
  buf(\xm8051_golden_model_1.n0884 [69], \xm8051_golden_model_1.n0897 [69]);
  buf(\xm8051_golden_model_1.n0884 [70], \xm8051_golden_model_1.n0897 [70]);
  buf(\xm8051_golden_model_1.n0884 [71], \xm8051_golden_model_1.n0897 [71]);
  buf(\xm8051_golden_model_1.n0884 [72], \xm8051_golden_model_1.n0896 [72]);
  buf(\xm8051_golden_model_1.n0884 [73], \xm8051_golden_model_1.n0896 [73]);
  buf(\xm8051_golden_model_1.n0884 [74], \xm8051_golden_model_1.n0896 [74]);
  buf(\xm8051_golden_model_1.n0884 [75], \xm8051_golden_model_1.n0896 [75]);
  buf(\xm8051_golden_model_1.n0884 [76], \xm8051_golden_model_1.n0896 [76]);
  buf(\xm8051_golden_model_1.n0884 [77], \xm8051_golden_model_1.n0896 [77]);
  buf(\xm8051_golden_model_1.n0884 [78], \xm8051_golden_model_1.n0896 [78]);
  buf(\xm8051_golden_model_1.n0884 [79], \xm8051_golden_model_1.n0896 [79]);
  buf(\xm8051_golden_model_1.n0884 [80], \xm8051_golden_model_1.n0895 [80]);
  buf(\xm8051_golden_model_1.n0884 [81], \xm8051_golden_model_1.n0895 [81]);
  buf(\xm8051_golden_model_1.n0884 [82], \xm8051_golden_model_1.n0895 [82]);
  buf(\xm8051_golden_model_1.n0884 [83], \xm8051_golden_model_1.n0895 [83]);
  buf(\xm8051_golden_model_1.n0884 [84], \xm8051_golden_model_1.n0895 [84]);
  buf(\xm8051_golden_model_1.n0884 [85], \xm8051_golden_model_1.n0895 [85]);
  buf(\xm8051_golden_model_1.n0884 [86], \xm8051_golden_model_1.n0895 [86]);
  buf(\xm8051_golden_model_1.n0884 [87], \xm8051_golden_model_1.n0895 [87]);
  buf(\xm8051_golden_model_1.n0884 [88], \xm8051_golden_model_1.n0894 [88]);
  buf(\xm8051_golden_model_1.n0884 [89], \xm8051_golden_model_1.n0894 [89]);
  buf(\xm8051_golden_model_1.n0884 [90], \xm8051_golden_model_1.n0894 [90]);
  buf(\xm8051_golden_model_1.n0884 [91], \xm8051_golden_model_1.n0894 [91]);
  buf(\xm8051_golden_model_1.n0884 [92], \xm8051_golden_model_1.n0894 [92]);
  buf(\xm8051_golden_model_1.n0884 [93], \xm8051_golden_model_1.n0894 [93]);
  buf(\xm8051_golden_model_1.n0884 [94], \xm8051_golden_model_1.n0894 [94]);
  buf(\xm8051_golden_model_1.n0884 [95], \xm8051_golden_model_1.n0894 [95]);
  buf(\xm8051_golden_model_1.n0884 [96], proc_data_in[0]);
  buf(\xm8051_golden_model_1.n0884 [97], proc_data_in[1]);
  buf(\xm8051_golden_model_1.n0884 [98], proc_data_in[2]);
  buf(\xm8051_golden_model_1.n0884 [99], proc_data_in[3]);
  buf(\xm8051_golden_model_1.n0884 [100], proc_data_in[4]);
  buf(\xm8051_golden_model_1.n0884 [101], proc_data_in[5]);
  buf(\xm8051_golden_model_1.n0884 [102], proc_data_in[6]);
  buf(\xm8051_golden_model_1.n0884 [103], proc_data_in[7]);
  buf(\xm8051_golden_model_1.n0884 [104], \xm8051_golden_model_1.n0892 [104]);
  buf(\xm8051_golden_model_1.n0884 [105], \xm8051_golden_model_1.n0892 [105]);
  buf(\xm8051_golden_model_1.n0884 [106], \xm8051_golden_model_1.n0892 [106]);
  buf(\xm8051_golden_model_1.n0884 [107], \xm8051_golden_model_1.n0892 [107]);
  buf(\xm8051_golden_model_1.n0884 [108], \xm8051_golden_model_1.n0892 [108]);
  buf(\xm8051_golden_model_1.n0884 [109], \xm8051_golden_model_1.n0892 [109]);
  buf(\xm8051_golden_model_1.n0884 [110], \xm8051_golden_model_1.n0892 [110]);
  buf(\xm8051_golden_model_1.n0884 [111], \xm8051_golden_model_1.n0892 [111]);
  buf(\xm8051_golden_model_1.n0884 [112], \xm8051_golden_model_1.n0891 [112]);
  buf(\xm8051_golden_model_1.n0884 [113], \xm8051_golden_model_1.n0891 [113]);
  buf(\xm8051_golden_model_1.n0884 [114], \xm8051_golden_model_1.n0891 [114]);
  buf(\xm8051_golden_model_1.n0884 [115], \xm8051_golden_model_1.n0891 [115]);
  buf(\xm8051_golden_model_1.n0884 [116], \xm8051_golden_model_1.n0891 [116]);
  buf(\xm8051_golden_model_1.n0884 [117], \xm8051_golden_model_1.n0891 [117]);
  buf(\xm8051_golden_model_1.n0884 [118], \xm8051_golden_model_1.n0891 [118]);
  buf(\xm8051_golden_model_1.n0884 [119], \xm8051_golden_model_1.n0891 [119]);
  buf(\xm8051_golden_model_1.n0884 [120], \xm8051_golden_model_1.n0889 [120]);
  buf(\xm8051_golden_model_1.n0884 [121], \xm8051_golden_model_1.n0889 [121]);
  buf(\xm8051_golden_model_1.n0884 [122], \xm8051_golden_model_1.n0889 [122]);
  buf(\xm8051_golden_model_1.n0884 [123], \xm8051_golden_model_1.n0889 [123]);
  buf(\xm8051_golden_model_1.n0884 [124], \xm8051_golden_model_1.n0889 [124]);
  buf(\xm8051_golden_model_1.n0884 [125], \xm8051_golden_model_1.n0889 [125]);
  buf(\xm8051_golden_model_1.n0884 [126], \xm8051_golden_model_1.n0889 [126]);
  buf(\xm8051_golden_model_1.n0884 [127], \xm8051_golden_model_1.n0889 [127]);
  buf(sha_state_impl[0], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [0]);
  buf(sha_state_impl[1], \oc8051_xiommu_impl_1.sha_top_i.sha_reg_state [1]);
  buf(aes_state_impl[0], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [0]);
  buf(aes_state_impl[1], \oc8051_xiommu_impl_1.aes_top_i.aes_reg_state [1]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.rst , rst);
  buf(datain[0], proc_data_in[0]);
  buf(datain[1], proc_data_in[1]);
  buf(datain[2], proc_data_in[2]);
  buf(datain[3], proc_data_in[3]);
  buf(datain[4], proc_data_in[4]);
  buf(datain[5], proc_data_in[5]);
  buf(datain[6], proc_data_in[6]);
  buf(datain[7], proc_data_in[7]);
  buf(addrin[0], proc_addr[0]);
  buf(addrin[1], proc_addr[1]);
  buf(addrin[2], proc_addr[2]);
  buf(addrin[3], proc_addr[3]);
  buf(addrin[4], proc_addr[4]);
  buf(addrin[5], proc_addr[5]);
  buf(addrin[6], proc_addr[6]);
  buf(addrin[7], proc_addr[7]);
  buf(addrin[8], proc_addr[8]);
  buf(addrin[9], proc_addr[9]);
  buf(addrin[10], proc_addr[10]);
  buf(addrin[11], proc_addr[11]);
  buf(addrin[12], proc_addr[12]);
  buf(addrin[13], proc_addr[13]);
  buf(addrin[14], proc_addr[14]);
  buf(addrin[15], proc_addr[15]);
  buf(\oc8051_xiommu_impl_1.aes_top_i.aes_reg_key1_i.clk , clk);
endmodule
